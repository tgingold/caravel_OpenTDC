magic
tech sky130A
magscale 1 2
timestamp 1607276039
<< viali >>
rect 7389 20349 7423 20383
rect 7573 20213 7607 20247
rect 7941 20213 7975 20247
rect 4353 18581 4387 18615
rect 8401 18173 8435 18207
rect 8953 18173 8987 18207
rect 4169 18105 4203 18139
rect 5457 18037 5491 18071
rect 8585 18037 8619 18071
rect 2789 15045 2823 15079
rect 2605 14909 2639 14943
rect 3249 14773 3283 14807
rect 6837 14569 6871 14603
rect 1409 14433 1443 14467
rect 1593 14229 1627 14263
rect 1593 14025 1627 14059
rect 8125 14025 8159 14059
rect 6837 13821 6871 13855
rect 6837 12733 6871 12767
rect 8401 12733 8435 12767
rect 8953 12733 8987 12767
rect 7021 12597 7055 12631
rect 7389 12597 7423 12631
rect 8585 12597 8619 12631
rect 4997 11849 5031 11883
rect 4813 11713 4847 11747
rect 6929 11169 6963 11203
rect 7113 11033 7147 11067
rect 8585 10761 8619 10795
rect 7481 10557 7515 10591
rect 7757 10557 7791 10591
rect 8401 10557 8435 10591
rect 8953 10557 8987 10591
rect 7113 10421 7147 10455
rect 5733 9061 5767 9095
rect 7021 8789 7055 8823
rect 5825 8585 5859 8619
rect 2421 8041 2455 8075
rect 5733 7973 5767 8007
rect 2237 7905 2271 7939
rect 7021 7701 7055 7735
rect 5825 7497 5859 7531
rect 2329 7157 2363 7191
rect 7021 6409 7055 6443
rect 6837 6205 6871 6239
rect 7481 6069 7515 6103
rect 8585 5865 8619 5899
rect 8401 5729 8435 5763
rect 4445 5321 4479 5355
rect 4905 5321 4939 5355
rect 4261 5117 4295 5151
rect 8401 4981 8435 5015
rect 2789 4165 2823 4199
rect 1409 4029 1443 4063
rect 2053 4029 2087 4063
rect 2605 4029 2639 4063
rect 3249 4029 3283 4063
rect 8309 4029 8343 4063
rect 8861 4029 8895 4063
rect 1593 3893 1627 3927
rect 8493 3893 8527 3927
<< metal1 >>
rect 1104 22330 9752 22352
rect 1104 22278 3872 22330
rect 3924 22278 3936 22330
rect 3988 22278 4000 22330
rect 4052 22278 4064 22330
rect 4116 22278 6763 22330
rect 6815 22278 6827 22330
rect 6879 22278 6891 22330
rect 6943 22278 6955 22330
rect 7007 22278 9752 22330
rect 1104 22256 9752 22278
rect 1104 21786 9752 21808
rect 1104 21734 2427 21786
rect 2479 21734 2491 21786
rect 2543 21734 2555 21786
rect 2607 21734 2619 21786
rect 2671 21734 5318 21786
rect 5370 21734 5382 21786
rect 5434 21734 5446 21786
rect 5498 21734 5510 21786
rect 5562 21734 8208 21786
rect 8260 21734 8272 21786
rect 8324 21734 8336 21786
rect 8388 21734 8400 21786
rect 8452 21734 9752 21786
rect 1104 21712 9752 21734
rect 1104 21242 9752 21264
rect 1104 21190 3872 21242
rect 3924 21190 3936 21242
rect 3988 21190 4000 21242
rect 4052 21190 4064 21242
rect 4116 21190 6763 21242
rect 6815 21190 6827 21242
rect 6879 21190 6891 21242
rect 6943 21190 6955 21242
rect 7007 21190 9752 21242
rect 1104 21168 9752 21190
rect 1104 20698 9752 20720
rect 1104 20646 2427 20698
rect 2479 20646 2491 20698
rect 2543 20646 2555 20698
rect 2607 20646 2619 20698
rect 2671 20646 5318 20698
rect 5370 20646 5382 20698
rect 5434 20646 5446 20698
rect 5498 20646 5510 20698
rect 5562 20646 8208 20698
rect 8260 20646 8272 20698
rect 8324 20646 8336 20698
rect 8388 20646 8400 20698
rect 8452 20646 9752 20698
rect 1104 20624 9752 20646
rect 7377 20383 7435 20389
rect 7377 20349 7389 20383
rect 7423 20380 7435 20383
rect 7423 20352 7972 20380
rect 7423 20349 7435 20352
rect 7377 20343 7435 20349
rect 7944 20256 7972 20352
rect 5166 20204 5172 20256
rect 5224 20244 5230 20256
rect 7561 20247 7619 20253
rect 7561 20244 7573 20247
rect 5224 20216 7573 20244
rect 5224 20204 5230 20216
rect 7561 20213 7573 20216
rect 7607 20213 7619 20247
rect 7926 20244 7932 20256
rect 7887 20216 7932 20244
rect 7561 20207 7619 20213
rect 7926 20204 7932 20216
rect 7984 20204 7990 20256
rect 1104 20154 9752 20176
rect 1104 20102 3872 20154
rect 3924 20102 3936 20154
rect 3988 20102 4000 20154
rect 4052 20102 4064 20154
rect 4116 20102 6763 20154
rect 6815 20102 6827 20154
rect 6879 20102 6891 20154
rect 6943 20102 6955 20154
rect 7007 20102 9752 20154
rect 1104 20080 9752 20102
rect 2314 20000 2320 20052
rect 2372 20040 2378 20052
rect 6270 20040 6276 20052
rect 2372 20012 6276 20040
rect 2372 20000 2378 20012
rect 6270 20000 6276 20012
rect 6328 20000 6334 20052
rect 1104 19610 9752 19632
rect 1104 19558 2427 19610
rect 2479 19558 2491 19610
rect 2543 19558 2555 19610
rect 2607 19558 2619 19610
rect 2671 19558 5318 19610
rect 5370 19558 5382 19610
rect 5434 19558 5446 19610
rect 5498 19558 5510 19610
rect 5562 19558 8208 19610
rect 8260 19558 8272 19610
rect 8324 19558 8336 19610
rect 8388 19558 8400 19610
rect 8452 19558 9752 19610
rect 1104 19536 9752 19558
rect 4430 19320 4436 19372
rect 4488 19360 4494 19372
rect 5626 19360 5632 19372
rect 4488 19332 5632 19360
rect 4488 19320 4494 19332
rect 5626 19320 5632 19332
rect 5684 19320 5690 19372
rect 1104 19066 9752 19088
rect 1104 19014 3872 19066
rect 3924 19014 3936 19066
rect 3988 19014 4000 19066
rect 4052 19014 4064 19066
rect 4116 19014 6763 19066
rect 6815 19014 6827 19066
rect 6879 19014 6891 19066
rect 6943 19014 6955 19066
rect 7007 19014 9752 19066
rect 1104 18992 9752 19014
rect 4338 18612 4344 18624
rect 4299 18584 4344 18612
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 1104 18522 9752 18544
rect 1104 18470 2427 18522
rect 2479 18470 2491 18522
rect 2543 18470 2555 18522
rect 2607 18470 2619 18522
rect 2671 18470 5318 18522
rect 5370 18470 5382 18522
rect 5434 18470 5446 18522
rect 5498 18470 5510 18522
rect 5562 18470 8208 18522
rect 8260 18470 8272 18522
rect 8324 18470 8336 18522
rect 8388 18470 8400 18522
rect 8452 18470 9752 18522
rect 1104 18448 9752 18470
rect 7374 18164 7380 18216
rect 7432 18204 7438 18216
rect 7926 18204 7932 18216
rect 7432 18176 7932 18204
rect 7432 18164 7438 18176
rect 7926 18164 7932 18176
rect 7984 18204 7990 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 7984 18176 8401 18204
rect 7984 18164 7990 18176
rect 8389 18173 8401 18176
rect 8435 18204 8447 18207
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8435 18176 8953 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 4157 18139 4215 18145
rect 4157 18105 4169 18139
rect 4203 18136 4215 18139
rect 4338 18136 4344 18148
rect 4203 18108 4344 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4338 18096 4344 18108
rect 4396 18136 4402 18148
rect 6546 18136 6552 18148
rect 4396 18108 6552 18136
rect 4396 18096 4402 18108
rect 6546 18096 6552 18108
rect 6604 18096 6610 18148
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 5445 18071 5503 18077
rect 5445 18068 5457 18071
rect 5132 18040 5457 18068
rect 5132 18028 5138 18040
rect 5445 18037 5457 18040
rect 5491 18037 5503 18071
rect 5445 18031 5503 18037
rect 8202 18028 8208 18080
rect 8260 18068 8266 18080
rect 8573 18071 8631 18077
rect 8573 18068 8585 18071
rect 8260 18040 8585 18068
rect 8260 18028 8266 18040
rect 8573 18037 8585 18040
rect 8619 18037 8631 18071
rect 8573 18031 8631 18037
rect 1104 17978 9752 18000
rect 1104 17926 3872 17978
rect 3924 17926 3936 17978
rect 3988 17926 4000 17978
rect 4052 17926 4064 17978
rect 4116 17926 6763 17978
rect 6815 17926 6827 17978
rect 6879 17926 6891 17978
rect 6943 17926 6955 17978
rect 7007 17926 9752 17978
rect 1104 17904 9752 17926
rect 1104 17434 9752 17456
rect 1104 17382 2427 17434
rect 2479 17382 2491 17434
rect 2543 17382 2555 17434
rect 2607 17382 2619 17434
rect 2671 17382 5318 17434
rect 5370 17382 5382 17434
rect 5434 17382 5446 17434
rect 5498 17382 5510 17434
rect 5562 17382 8208 17434
rect 8260 17382 8272 17434
rect 8324 17382 8336 17434
rect 8388 17382 8400 17434
rect 8452 17382 9752 17434
rect 1104 17360 9752 17382
rect 1104 16890 9752 16912
rect 1104 16838 3872 16890
rect 3924 16838 3936 16890
rect 3988 16838 4000 16890
rect 4052 16838 4064 16890
rect 4116 16838 6763 16890
rect 6815 16838 6827 16890
rect 6879 16838 6891 16890
rect 6943 16838 6955 16890
rect 7007 16838 9752 16890
rect 1104 16816 9752 16838
rect 1104 16346 9752 16368
rect 1104 16294 2427 16346
rect 2479 16294 2491 16346
rect 2543 16294 2555 16346
rect 2607 16294 2619 16346
rect 2671 16294 5318 16346
rect 5370 16294 5382 16346
rect 5434 16294 5446 16346
rect 5498 16294 5510 16346
rect 5562 16294 8208 16346
rect 8260 16294 8272 16346
rect 8324 16294 8336 16346
rect 8388 16294 8400 16346
rect 8452 16294 9752 16346
rect 1104 16272 9752 16294
rect 1104 15802 9752 15824
rect 1104 15750 3872 15802
rect 3924 15750 3936 15802
rect 3988 15750 4000 15802
rect 4052 15750 4064 15802
rect 4116 15750 6763 15802
rect 6815 15750 6827 15802
rect 6879 15750 6891 15802
rect 6943 15750 6955 15802
rect 7007 15750 9752 15802
rect 1104 15728 9752 15750
rect 1104 15258 9752 15280
rect 1104 15206 2427 15258
rect 2479 15206 2491 15258
rect 2543 15206 2555 15258
rect 2607 15206 2619 15258
rect 2671 15206 5318 15258
rect 5370 15206 5382 15258
rect 5434 15206 5446 15258
rect 5498 15206 5510 15258
rect 5562 15206 8208 15258
rect 8260 15206 8272 15258
rect 8324 15206 8336 15258
rect 8388 15206 8400 15258
rect 8452 15206 9752 15258
rect 1104 15184 9752 15206
rect 2777 15079 2835 15085
rect 2777 15045 2789 15079
rect 2823 15076 2835 15079
rect 6178 15076 6184 15088
rect 2823 15048 6184 15076
rect 2823 15045 2835 15048
rect 2777 15039 2835 15045
rect 6178 15036 6184 15048
rect 6236 15036 6242 15088
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 2593 14943 2651 14949
rect 2593 14940 2605 14943
rect 1452 14912 2605 14940
rect 1452 14900 1458 14912
rect 2593 14909 2605 14912
rect 2639 14940 2651 14943
rect 2639 14912 3280 14940
rect 2639 14909 2651 14912
rect 2593 14903 2651 14909
rect 3252 14813 3280 14912
rect 3237 14807 3295 14813
rect 3237 14773 3249 14807
rect 3283 14804 3295 14807
rect 7374 14804 7380 14816
rect 3283 14776 7380 14804
rect 3283 14773 3295 14776
rect 3237 14767 3295 14773
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 1104 14714 9752 14736
rect 1104 14662 3872 14714
rect 3924 14662 3936 14714
rect 3988 14662 4000 14714
rect 4052 14662 4064 14714
rect 4116 14662 6763 14714
rect 6815 14662 6827 14714
rect 6879 14662 6891 14714
rect 6943 14662 6955 14714
rect 7007 14662 9752 14714
rect 1104 14640 9752 14662
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6604 14572 6837 14600
rect 6604 14560 6610 14572
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 5626 14260 5632 14272
rect 1627 14232 5632 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 1104 14170 9752 14192
rect 1104 14118 2427 14170
rect 2479 14118 2491 14170
rect 2543 14118 2555 14170
rect 2607 14118 2619 14170
rect 2671 14118 5318 14170
rect 5370 14118 5382 14170
rect 5434 14118 5446 14170
rect 5498 14118 5510 14170
rect 5562 14118 8208 14170
rect 8260 14118 8272 14170
rect 8324 14118 8336 14170
rect 8388 14118 8400 14170
rect 8452 14118 9752 14170
rect 1104 14096 9752 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1452 14028 1593 14056
rect 1452 14016 1458 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 6328 14028 8125 14056
rect 6328 14016 6334 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 8113 14019 8171 14025
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6546 13852 6552 13864
rect 6420 13824 6552 13852
rect 6420 13812 6426 13824
rect 6546 13812 6552 13824
rect 6604 13852 6610 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6604 13824 6837 13852
rect 6604 13812 6610 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 1104 13626 9752 13648
rect 1104 13574 3872 13626
rect 3924 13574 3936 13626
rect 3988 13574 4000 13626
rect 4052 13574 4064 13626
rect 4116 13574 6763 13626
rect 6815 13574 6827 13626
rect 6879 13574 6891 13626
rect 6943 13574 6955 13626
rect 7007 13574 9752 13626
rect 1104 13552 9752 13574
rect 1104 13082 9752 13104
rect 1104 13030 2427 13082
rect 2479 13030 2491 13082
rect 2543 13030 2555 13082
rect 2607 13030 2619 13082
rect 2671 13030 5318 13082
rect 5370 13030 5382 13082
rect 5434 13030 5446 13082
rect 5498 13030 5510 13082
rect 5562 13030 8208 13082
rect 8260 13030 8272 13082
rect 8324 13030 8336 13082
rect 8388 13030 8400 13082
rect 8452 13030 9752 13082
rect 1104 13008 9752 13030
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 6871 12736 8401 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7392 12640 7420 12736
rect 8389 12733 8401 12736
rect 8435 12764 8447 12767
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8435 12736 8953 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 6604 12600 7021 12628
rect 6604 12588 6610 12600
rect 7009 12597 7021 12600
rect 7055 12597 7067 12631
rect 7374 12628 7380 12640
rect 7335 12600 7380 12628
rect 7009 12591 7067 12597
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 8570 12628 8576 12640
rect 8531 12600 8576 12628
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 1104 12538 9752 12560
rect 1104 12486 3872 12538
rect 3924 12486 3936 12538
rect 3988 12486 4000 12538
rect 4052 12486 4064 12538
rect 4116 12486 6763 12538
rect 6815 12486 6827 12538
rect 6879 12486 6891 12538
rect 6943 12486 6955 12538
rect 7007 12486 9752 12538
rect 1104 12464 9752 12486
rect 1104 11994 9752 12016
rect 1104 11942 2427 11994
rect 2479 11942 2491 11994
rect 2543 11942 2555 11994
rect 2607 11942 2619 11994
rect 2671 11942 5318 11994
rect 5370 11942 5382 11994
rect 5434 11942 5446 11994
rect 5498 11942 5510 11994
rect 5562 11942 8208 11994
rect 8260 11942 8272 11994
rect 8324 11942 8336 11994
rect 8388 11942 8400 11994
rect 8452 11942 9752 11994
rect 1104 11920 9752 11942
rect 4985 11883 5043 11889
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 7374 11880 7380 11892
rect 5031 11852 7380 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 3476 11716 4813 11744
rect 3476 11704 3482 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 1104 11450 9752 11472
rect 1104 11398 3872 11450
rect 3924 11398 3936 11450
rect 3988 11398 4000 11450
rect 4052 11398 4064 11450
rect 4116 11398 6763 11450
rect 6815 11398 6827 11450
rect 6879 11398 6891 11450
rect 6943 11398 6955 11450
rect 7007 11398 9752 11450
rect 1104 11376 9752 11398
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7374 11200 7380 11212
rect 6963 11172 7380 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 5626 11064 5632 11076
rect 2832 11036 5632 11064
rect 2832 11024 2838 11036
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 6696 11036 7113 11064
rect 6696 11024 6702 11036
rect 7101 11033 7113 11036
rect 7147 11033 7159 11067
rect 7101 11027 7159 11033
rect 1104 10906 9752 10928
rect 1104 10854 2427 10906
rect 2479 10854 2491 10906
rect 2543 10854 2555 10906
rect 2607 10854 2619 10906
rect 2671 10854 5318 10906
rect 5370 10854 5382 10906
rect 5434 10854 5446 10906
rect 5498 10854 5510 10906
rect 5562 10854 8208 10906
rect 8260 10854 8272 10906
rect 8324 10854 8336 10906
rect 8388 10854 8400 10906
rect 8452 10854 9752 10906
rect 1104 10832 9752 10854
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 6788 10764 8585 10792
rect 6788 10752 6794 10764
rect 8573 10761 8585 10764
rect 8619 10761 8631 10795
rect 8573 10755 8631 10761
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 6420 10560 7481 10588
rect 6420 10548 6426 10560
rect 7469 10557 7481 10560
rect 7515 10588 7527 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7515 10560 7757 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8435 10560 8953 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 8404 10520 8432 10551
rect 7392 10492 8432 10520
rect 7392 10464 7420 10492
rect 7101 10455 7159 10461
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 7374 10452 7380 10464
rect 7147 10424 7380 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 1104 10362 9752 10384
rect 1104 10310 3872 10362
rect 3924 10310 3936 10362
rect 3988 10310 4000 10362
rect 4052 10310 4064 10362
rect 4116 10310 6763 10362
rect 6815 10310 6827 10362
rect 6879 10310 6891 10362
rect 6943 10310 6955 10362
rect 7007 10310 9752 10362
rect 1104 10288 9752 10310
rect 1104 9818 9752 9840
rect 1104 9766 2427 9818
rect 2479 9766 2491 9818
rect 2543 9766 2555 9818
rect 2607 9766 2619 9818
rect 2671 9766 5318 9818
rect 5370 9766 5382 9818
rect 5434 9766 5446 9818
rect 5498 9766 5510 9818
rect 5562 9766 8208 9818
rect 8260 9766 8272 9818
rect 8324 9766 8336 9818
rect 8388 9766 8400 9818
rect 8452 9766 9752 9818
rect 1104 9744 9752 9766
rect 1104 9274 9752 9296
rect 1104 9222 3872 9274
rect 3924 9222 3936 9274
rect 3988 9222 4000 9274
rect 4052 9222 4064 9274
rect 4116 9222 6763 9274
rect 6815 9222 6827 9274
rect 6879 9222 6891 9274
rect 6943 9222 6955 9274
rect 7007 9222 9752 9274
rect 1104 9200 9752 9222
rect 5721 9095 5779 9101
rect 5721 9061 5733 9095
rect 5767 9092 5779 9095
rect 5810 9092 5816 9104
rect 5767 9064 5816 9092
rect 5767 9061 5779 9064
rect 5721 9055 5779 9061
rect 5810 9052 5816 9064
rect 5868 9092 5874 9104
rect 6362 9092 6368 9104
rect 5868 9064 6368 9092
rect 5868 9052 5874 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 3384 8792 7021 8820
rect 3384 8780 3390 8792
rect 7009 8789 7021 8792
rect 7055 8789 7067 8823
rect 7009 8783 7067 8789
rect 1104 8730 9752 8752
rect 1104 8678 2427 8730
rect 2479 8678 2491 8730
rect 2543 8678 2555 8730
rect 2607 8678 2619 8730
rect 2671 8678 5318 8730
rect 5370 8678 5382 8730
rect 5434 8678 5446 8730
rect 5498 8678 5510 8730
rect 5562 8678 8208 8730
rect 8260 8678 8272 8730
rect 8324 8678 8336 8730
rect 8388 8678 8400 8730
rect 8452 8678 9752 8730
rect 1104 8656 9752 8678
rect 5810 8616 5816 8628
rect 5771 8588 5816 8616
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 1104 8186 9752 8208
rect 1104 8134 3872 8186
rect 3924 8134 3936 8186
rect 3988 8134 4000 8186
rect 4052 8134 4064 8186
rect 4116 8134 6763 8186
rect 6815 8134 6827 8186
rect 6879 8134 6891 8186
rect 6943 8134 6955 8186
rect 7007 8134 9752 8186
rect 1104 8112 9752 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2774 8072 2780 8084
rect 2455 8044 2780 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 8004 5779 8007
rect 5810 8004 5816 8016
rect 5767 7976 5816 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 5810 7964 5816 7976
rect 5868 7964 5874 8016
rect 2222 7936 2228 7948
rect 2183 7908 2228 7936
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 5776 7704 7021 7732
rect 5776 7692 5782 7704
rect 7009 7701 7021 7704
rect 7055 7701 7067 7735
rect 7009 7695 7067 7701
rect 1104 7642 9752 7664
rect 1104 7590 2427 7642
rect 2479 7590 2491 7642
rect 2543 7590 2555 7642
rect 2607 7590 2619 7642
rect 2671 7590 5318 7642
rect 5370 7590 5382 7642
rect 5434 7590 5446 7642
rect 5498 7590 5510 7642
rect 5562 7590 8208 7642
rect 8260 7590 8272 7642
rect 8324 7590 8336 7642
rect 8388 7590 8400 7642
rect 8452 7590 9752 7642
rect 1104 7568 9752 7590
rect 5810 7528 5816 7540
rect 5771 7500 5816 7528
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2317 7191 2375 7197
rect 2317 7188 2329 7191
rect 2280 7160 2329 7188
rect 2280 7148 2286 7160
rect 2317 7157 2329 7160
rect 2363 7188 2375 7191
rect 4890 7188 4896 7200
rect 2363 7160 4896 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 1104 7098 9752 7120
rect 1104 7046 3872 7098
rect 3924 7046 3936 7098
rect 3988 7046 4000 7098
rect 4052 7046 4064 7098
rect 4116 7046 6763 7098
rect 6815 7046 6827 7098
rect 6879 7046 6891 7098
rect 6943 7046 6955 7098
rect 7007 7046 9752 7098
rect 1104 7024 9752 7046
rect 1104 6554 9752 6576
rect 1104 6502 2427 6554
rect 2479 6502 2491 6554
rect 2543 6502 2555 6554
rect 2607 6502 2619 6554
rect 2671 6502 5318 6554
rect 5370 6502 5382 6554
rect 5434 6502 5446 6554
rect 5498 6502 5510 6554
rect 5562 6502 8208 6554
rect 8260 6502 8272 6554
rect 8324 6502 8336 6554
rect 8388 6502 8400 6554
rect 8452 6502 9752 6554
rect 1104 6480 9752 6502
rect 7009 6443 7067 6449
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 7098 6440 7104 6452
rect 7055 6412 7104 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 4948 6208 6837 6236
rect 4948 6196 4954 6208
rect 6825 6205 6837 6208
rect 6871 6236 6883 6239
rect 7374 6236 7380 6248
rect 6871 6208 7380 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7374 6196 7380 6208
rect 7432 6236 7438 6248
rect 7432 6208 7512 6236
rect 7432 6196 7438 6208
rect 7484 6109 7512 6208
rect 7469 6103 7527 6109
rect 7469 6069 7481 6103
rect 7515 6100 7527 6103
rect 7926 6100 7932 6112
rect 7515 6072 7932 6100
rect 7515 6069 7527 6072
rect 7469 6063 7527 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 1104 6010 9752 6032
rect 1104 5958 3872 6010
rect 3924 5958 3936 6010
rect 3988 5958 4000 6010
rect 4052 5958 4064 6010
rect 4116 5958 6763 6010
rect 6815 5958 6827 6010
rect 6879 5958 6891 6010
rect 6943 5958 6955 6010
rect 7007 5958 9752 6010
rect 1104 5936 9752 5958
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 6512 5868 8585 5896
rect 6512 5856 6518 5868
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 8573 5859 8631 5865
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 7984 5732 8401 5760
rect 7984 5720 7990 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 8389 5723 8447 5729
rect 1104 5466 9752 5488
rect 1104 5414 2427 5466
rect 2479 5414 2491 5466
rect 2543 5414 2555 5466
rect 2607 5414 2619 5466
rect 2671 5414 5318 5466
rect 5370 5414 5382 5466
rect 5434 5414 5446 5466
rect 5498 5414 5510 5466
rect 5562 5414 8208 5466
rect 8260 5414 8272 5466
rect 8324 5414 8336 5466
rect 8388 5414 8400 5466
rect 8452 5414 9752 5466
rect 1104 5392 9752 5414
rect 4430 5352 4436 5364
rect 4391 5324 4436 5352
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 4890 5352 4896 5364
rect 4851 5324 4896 5352
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 4246 5148 4252 5160
rect 4159 5120 4252 5148
rect 4246 5108 4252 5120
rect 4304 5148 4310 5160
rect 4890 5148 4896 5160
rect 4304 5120 4896 5148
rect 4304 5108 4310 5120
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 7984 4984 8401 5012
rect 7984 4972 7990 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8389 4975 8447 4981
rect 1104 4922 9752 4944
rect 1104 4870 3872 4922
rect 3924 4870 3936 4922
rect 3988 4870 4000 4922
rect 4052 4870 4064 4922
rect 4116 4870 6763 4922
rect 6815 4870 6827 4922
rect 6879 4870 6891 4922
rect 6943 4870 6955 4922
rect 7007 4870 9752 4922
rect 1104 4848 9752 4870
rect 1104 4378 9752 4400
rect 1104 4326 2427 4378
rect 2479 4326 2491 4378
rect 2543 4326 2555 4378
rect 2607 4326 2619 4378
rect 2671 4326 5318 4378
rect 5370 4326 5382 4378
rect 5434 4326 5446 4378
rect 5498 4326 5510 4378
rect 5562 4326 8208 4378
rect 8260 4326 8272 4378
rect 8324 4326 8336 4378
rect 8388 4326 8400 4378
rect 8452 4326 9752 4378
rect 1104 4304 9752 4326
rect 2777 4199 2835 4205
rect 2777 4165 2789 4199
rect 2823 4165 2835 4199
rect 5626 4196 5632 4208
rect 2777 4159 2835 4165
rect 4816 4168 5632 4196
rect 2792 4128 2820 4159
rect 4816 4128 4844 4168
rect 5626 4156 5632 4168
rect 5684 4156 5690 4208
rect 2792 4100 4844 4128
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 8938 4128 8944 4140
rect 5868 4100 8944 4128
rect 5868 4088 5874 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1443 4032 2053 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2041 4029 2053 4032
rect 2087 4060 2099 4063
rect 2593 4063 2651 4069
rect 2593 4060 2605 4063
rect 2087 4032 2605 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 2593 4029 2605 4032
rect 2639 4060 2651 4063
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 2639 4032 3249 4060
rect 2639 4029 2651 4032
rect 2593 4023 2651 4029
rect 3237 4029 3249 4032
rect 3283 4060 3295 4063
rect 4246 4060 4252 4072
rect 3283 4032 4252 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 4246 4020 4252 4032
rect 4304 4020 4310 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 7984 4032 8309 4060
rect 7984 4020 7990 4032
rect 8297 4029 8309 4032
rect 8343 4060 8355 4063
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8343 4032 8861 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 2866 3992 2872 4004
rect 1596 3964 2872 3992
rect 1596 3933 1624 3964
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8481 3927 8539 3933
rect 8481 3924 8493 3927
rect 8076 3896 8493 3924
rect 8076 3884 8082 3896
rect 8481 3893 8493 3896
rect 8527 3893 8539 3927
rect 8481 3887 8539 3893
rect 1104 3834 9752 3856
rect 1104 3782 3872 3834
rect 3924 3782 3936 3834
rect 3988 3782 4000 3834
rect 4052 3782 4064 3834
rect 4116 3782 6763 3834
rect 6815 3782 6827 3834
rect 6879 3782 6891 3834
rect 6943 3782 6955 3834
rect 7007 3782 9752 3834
rect 1104 3760 9752 3782
rect 1104 3290 9752 3312
rect 1104 3238 2427 3290
rect 2479 3238 2491 3290
rect 2543 3238 2555 3290
rect 2607 3238 2619 3290
rect 2671 3238 5318 3290
rect 5370 3238 5382 3290
rect 5434 3238 5446 3290
rect 5498 3238 5510 3290
rect 5562 3238 8208 3290
rect 8260 3238 8272 3290
rect 8324 3238 8336 3290
rect 8388 3238 8400 3290
rect 8452 3238 9752 3290
rect 1104 3216 9752 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 5718 3176 5724 3188
rect 1820 3148 5724 3176
rect 1820 3136 1826 3148
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 1104 2746 9752 2768
rect 1104 2694 3872 2746
rect 3924 2694 3936 2746
rect 3988 2694 4000 2746
rect 4052 2694 4064 2746
rect 4116 2694 6763 2746
rect 6815 2694 6827 2746
rect 6879 2694 6891 2746
rect 6943 2694 6955 2746
rect 7007 2694 9752 2746
rect 1104 2672 9752 2694
rect 1104 2202 9752 2224
rect 1104 2150 2427 2202
rect 2479 2150 2491 2202
rect 2543 2150 2555 2202
rect 2607 2150 2619 2202
rect 2671 2150 5318 2202
rect 5370 2150 5382 2202
rect 5434 2150 5446 2202
rect 5498 2150 5510 2202
rect 5562 2150 8208 2202
rect 8260 2150 8272 2202
rect 8324 2150 8336 2202
rect 8388 2150 8400 2202
rect 8452 2150 9752 2202
rect 1104 2128 9752 2150
<< via1 >>
rect 3872 22278 3924 22330
rect 3936 22278 3988 22330
rect 4000 22278 4052 22330
rect 4064 22278 4116 22330
rect 6763 22278 6815 22330
rect 6827 22278 6879 22330
rect 6891 22278 6943 22330
rect 6955 22278 7007 22330
rect 2427 21734 2479 21786
rect 2491 21734 2543 21786
rect 2555 21734 2607 21786
rect 2619 21734 2671 21786
rect 5318 21734 5370 21786
rect 5382 21734 5434 21786
rect 5446 21734 5498 21786
rect 5510 21734 5562 21786
rect 8208 21734 8260 21786
rect 8272 21734 8324 21786
rect 8336 21734 8388 21786
rect 8400 21734 8452 21786
rect 3872 21190 3924 21242
rect 3936 21190 3988 21242
rect 4000 21190 4052 21242
rect 4064 21190 4116 21242
rect 6763 21190 6815 21242
rect 6827 21190 6879 21242
rect 6891 21190 6943 21242
rect 6955 21190 7007 21242
rect 2427 20646 2479 20698
rect 2491 20646 2543 20698
rect 2555 20646 2607 20698
rect 2619 20646 2671 20698
rect 5318 20646 5370 20698
rect 5382 20646 5434 20698
rect 5446 20646 5498 20698
rect 5510 20646 5562 20698
rect 8208 20646 8260 20698
rect 8272 20646 8324 20698
rect 8336 20646 8388 20698
rect 8400 20646 8452 20698
rect 5172 20204 5224 20256
rect 7932 20247 7984 20256
rect 7932 20213 7941 20247
rect 7941 20213 7975 20247
rect 7975 20213 7984 20247
rect 7932 20204 7984 20213
rect 3872 20102 3924 20154
rect 3936 20102 3988 20154
rect 4000 20102 4052 20154
rect 4064 20102 4116 20154
rect 6763 20102 6815 20154
rect 6827 20102 6879 20154
rect 6891 20102 6943 20154
rect 6955 20102 7007 20154
rect 2320 20000 2372 20052
rect 6276 20000 6328 20052
rect 2427 19558 2479 19610
rect 2491 19558 2543 19610
rect 2555 19558 2607 19610
rect 2619 19558 2671 19610
rect 5318 19558 5370 19610
rect 5382 19558 5434 19610
rect 5446 19558 5498 19610
rect 5510 19558 5562 19610
rect 8208 19558 8260 19610
rect 8272 19558 8324 19610
rect 8336 19558 8388 19610
rect 8400 19558 8452 19610
rect 4436 19320 4488 19372
rect 5632 19320 5684 19372
rect 3872 19014 3924 19066
rect 3936 19014 3988 19066
rect 4000 19014 4052 19066
rect 4064 19014 4116 19066
rect 6763 19014 6815 19066
rect 6827 19014 6879 19066
rect 6891 19014 6943 19066
rect 6955 19014 7007 19066
rect 4344 18615 4396 18624
rect 4344 18581 4353 18615
rect 4353 18581 4387 18615
rect 4387 18581 4396 18615
rect 4344 18572 4396 18581
rect 2427 18470 2479 18522
rect 2491 18470 2543 18522
rect 2555 18470 2607 18522
rect 2619 18470 2671 18522
rect 5318 18470 5370 18522
rect 5382 18470 5434 18522
rect 5446 18470 5498 18522
rect 5510 18470 5562 18522
rect 8208 18470 8260 18522
rect 8272 18470 8324 18522
rect 8336 18470 8388 18522
rect 8400 18470 8452 18522
rect 7380 18164 7432 18216
rect 7932 18164 7984 18216
rect 4344 18096 4396 18148
rect 6552 18096 6604 18148
rect 5080 18028 5132 18080
rect 8208 18028 8260 18080
rect 3872 17926 3924 17978
rect 3936 17926 3988 17978
rect 4000 17926 4052 17978
rect 4064 17926 4116 17978
rect 6763 17926 6815 17978
rect 6827 17926 6879 17978
rect 6891 17926 6943 17978
rect 6955 17926 7007 17978
rect 2427 17382 2479 17434
rect 2491 17382 2543 17434
rect 2555 17382 2607 17434
rect 2619 17382 2671 17434
rect 5318 17382 5370 17434
rect 5382 17382 5434 17434
rect 5446 17382 5498 17434
rect 5510 17382 5562 17434
rect 8208 17382 8260 17434
rect 8272 17382 8324 17434
rect 8336 17382 8388 17434
rect 8400 17382 8452 17434
rect 3872 16838 3924 16890
rect 3936 16838 3988 16890
rect 4000 16838 4052 16890
rect 4064 16838 4116 16890
rect 6763 16838 6815 16890
rect 6827 16838 6879 16890
rect 6891 16838 6943 16890
rect 6955 16838 7007 16890
rect 2427 16294 2479 16346
rect 2491 16294 2543 16346
rect 2555 16294 2607 16346
rect 2619 16294 2671 16346
rect 5318 16294 5370 16346
rect 5382 16294 5434 16346
rect 5446 16294 5498 16346
rect 5510 16294 5562 16346
rect 8208 16294 8260 16346
rect 8272 16294 8324 16346
rect 8336 16294 8388 16346
rect 8400 16294 8452 16346
rect 3872 15750 3924 15802
rect 3936 15750 3988 15802
rect 4000 15750 4052 15802
rect 4064 15750 4116 15802
rect 6763 15750 6815 15802
rect 6827 15750 6879 15802
rect 6891 15750 6943 15802
rect 6955 15750 7007 15802
rect 2427 15206 2479 15258
rect 2491 15206 2543 15258
rect 2555 15206 2607 15258
rect 2619 15206 2671 15258
rect 5318 15206 5370 15258
rect 5382 15206 5434 15258
rect 5446 15206 5498 15258
rect 5510 15206 5562 15258
rect 8208 15206 8260 15258
rect 8272 15206 8324 15258
rect 8336 15206 8388 15258
rect 8400 15206 8452 15258
rect 6184 15036 6236 15088
rect 1400 14900 1452 14952
rect 7380 14764 7432 14816
rect 3872 14662 3924 14714
rect 3936 14662 3988 14714
rect 4000 14662 4052 14714
rect 4064 14662 4116 14714
rect 6763 14662 6815 14714
rect 6827 14662 6879 14714
rect 6891 14662 6943 14714
rect 6955 14662 7007 14714
rect 6552 14560 6604 14612
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 5632 14220 5684 14272
rect 2427 14118 2479 14170
rect 2491 14118 2543 14170
rect 2555 14118 2607 14170
rect 2619 14118 2671 14170
rect 5318 14118 5370 14170
rect 5382 14118 5434 14170
rect 5446 14118 5498 14170
rect 5510 14118 5562 14170
rect 8208 14118 8260 14170
rect 8272 14118 8324 14170
rect 8336 14118 8388 14170
rect 8400 14118 8452 14170
rect 1400 14016 1452 14068
rect 6276 14016 6328 14068
rect 6368 13812 6420 13864
rect 6552 13812 6604 13864
rect 3872 13574 3924 13626
rect 3936 13574 3988 13626
rect 4000 13574 4052 13626
rect 4064 13574 4116 13626
rect 6763 13574 6815 13626
rect 6827 13574 6879 13626
rect 6891 13574 6943 13626
rect 6955 13574 7007 13626
rect 2427 13030 2479 13082
rect 2491 13030 2543 13082
rect 2555 13030 2607 13082
rect 2619 13030 2671 13082
rect 5318 13030 5370 13082
rect 5382 13030 5434 13082
rect 5446 13030 5498 13082
rect 5510 13030 5562 13082
rect 8208 13030 8260 13082
rect 8272 13030 8324 13082
rect 8336 13030 8388 13082
rect 8400 13030 8452 13082
rect 6552 12588 6604 12640
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 3872 12486 3924 12538
rect 3936 12486 3988 12538
rect 4000 12486 4052 12538
rect 4064 12486 4116 12538
rect 6763 12486 6815 12538
rect 6827 12486 6879 12538
rect 6891 12486 6943 12538
rect 6955 12486 7007 12538
rect 2427 11942 2479 11994
rect 2491 11942 2543 11994
rect 2555 11942 2607 11994
rect 2619 11942 2671 11994
rect 5318 11942 5370 11994
rect 5382 11942 5434 11994
rect 5446 11942 5498 11994
rect 5510 11942 5562 11994
rect 8208 11942 8260 11994
rect 8272 11942 8324 11994
rect 8336 11942 8388 11994
rect 8400 11942 8452 11994
rect 7380 11840 7432 11892
rect 3424 11704 3476 11756
rect 3872 11398 3924 11450
rect 3936 11398 3988 11450
rect 4000 11398 4052 11450
rect 4064 11398 4116 11450
rect 6763 11398 6815 11450
rect 6827 11398 6879 11450
rect 6891 11398 6943 11450
rect 6955 11398 7007 11450
rect 7380 11160 7432 11212
rect 2780 11024 2832 11076
rect 5632 11024 5684 11076
rect 6644 11024 6696 11076
rect 2427 10854 2479 10906
rect 2491 10854 2543 10906
rect 2555 10854 2607 10906
rect 2619 10854 2671 10906
rect 5318 10854 5370 10906
rect 5382 10854 5434 10906
rect 5446 10854 5498 10906
rect 5510 10854 5562 10906
rect 8208 10854 8260 10906
rect 8272 10854 8324 10906
rect 8336 10854 8388 10906
rect 8400 10854 8452 10906
rect 6736 10752 6788 10804
rect 6368 10548 6420 10600
rect 7380 10412 7432 10464
rect 3872 10310 3924 10362
rect 3936 10310 3988 10362
rect 4000 10310 4052 10362
rect 4064 10310 4116 10362
rect 6763 10310 6815 10362
rect 6827 10310 6879 10362
rect 6891 10310 6943 10362
rect 6955 10310 7007 10362
rect 2427 9766 2479 9818
rect 2491 9766 2543 9818
rect 2555 9766 2607 9818
rect 2619 9766 2671 9818
rect 5318 9766 5370 9818
rect 5382 9766 5434 9818
rect 5446 9766 5498 9818
rect 5510 9766 5562 9818
rect 8208 9766 8260 9818
rect 8272 9766 8324 9818
rect 8336 9766 8388 9818
rect 8400 9766 8452 9818
rect 3872 9222 3924 9274
rect 3936 9222 3988 9274
rect 4000 9222 4052 9274
rect 4064 9222 4116 9274
rect 6763 9222 6815 9274
rect 6827 9222 6879 9274
rect 6891 9222 6943 9274
rect 6955 9222 7007 9274
rect 5816 9052 5868 9104
rect 6368 9052 6420 9104
rect 3332 8780 3384 8832
rect 2427 8678 2479 8730
rect 2491 8678 2543 8730
rect 2555 8678 2607 8730
rect 2619 8678 2671 8730
rect 5318 8678 5370 8730
rect 5382 8678 5434 8730
rect 5446 8678 5498 8730
rect 5510 8678 5562 8730
rect 8208 8678 8260 8730
rect 8272 8678 8324 8730
rect 8336 8678 8388 8730
rect 8400 8678 8452 8730
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 3872 8134 3924 8186
rect 3936 8134 3988 8186
rect 4000 8134 4052 8186
rect 4064 8134 4116 8186
rect 6763 8134 6815 8186
rect 6827 8134 6879 8186
rect 6891 8134 6943 8186
rect 6955 8134 7007 8186
rect 2780 8032 2832 8084
rect 5816 7964 5868 8016
rect 2228 7939 2280 7948
rect 2228 7905 2237 7939
rect 2237 7905 2271 7939
rect 2271 7905 2280 7939
rect 2228 7896 2280 7905
rect 5724 7692 5776 7744
rect 2427 7590 2479 7642
rect 2491 7590 2543 7642
rect 2555 7590 2607 7642
rect 2619 7590 2671 7642
rect 5318 7590 5370 7642
rect 5382 7590 5434 7642
rect 5446 7590 5498 7642
rect 5510 7590 5562 7642
rect 8208 7590 8260 7642
rect 8272 7590 8324 7642
rect 8336 7590 8388 7642
rect 8400 7590 8452 7642
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 2228 7148 2280 7200
rect 4896 7148 4948 7200
rect 3872 7046 3924 7098
rect 3936 7046 3988 7098
rect 4000 7046 4052 7098
rect 4064 7046 4116 7098
rect 6763 7046 6815 7098
rect 6827 7046 6879 7098
rect 6891 7046 6943 7098
rect 6955 7046 7007 7098
rect 2427 6502 2479 6554
rect 2491 6502 2543 6554
rect 2555 6502 2607 6554
rect 2619 6502 2671 6554
rect 5318 6502 5370 6554
rect 5382 6502 5434 6554
rect 5446 6502 5498 6554
rect 5510 6502 5562 6554
rect 8208 6502 8260 6554
rect 8272 6502 8324 6554
rect 8336 6502 8388 6554
rect 8400 6502 8452 6554
rect 7104 6400 7156 6452
rect 4896 6196 4948 6248
rect 7380 6196 7432 6248
rect 7932 6060 7984 6112
rect 3872 5958 3924 6010
rect 3936 5958 3988 6010
rect 4000 5958 4052 6010
rect 4064 5958 4116 6010
rect 6763 5958 6815 6010
rect 6827 5958 6879 6010
rect 6891 5958 6943 6010
rect 6955 5958 7007 6010
rect 6460 5856 6512 5908
rect 7932 5720 7984 5772
rect 2427 5414 2479 5466
rect 2491 5414 2543 5466
rect 2555 5414 2607 5466
rect 2619 5414 2671 5466
rect 5318 5414 5370 5466
rect 5382 5414 5434 5466
rect 5446 5414 5498 5466
rect 5510 5414 5562 5466
rect 8208 5414 8260 5466
rect 8272 5414 8324 5466
rect 8336 5414 8388 5466
rect 8400 5414 8452 5466
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 4896 5108 4948 5160
rect 7932 4972 7984 5024
rect 3872 4870 3924 4922
rect 3936 4870 3988 4922
rect 4000 4870 4052 4922
rect 4064 4870 4116 4922
rect 6763 4870 6815 4922
rect 6827 4870 6879 4922
rect 6891 4870 6943 4922
rect 6955 4870 7007 4922
rect 2427 4326 2479 4378
rect 2491 4326 2543 4378
rect 2555 4326 2607 4378
rect 2619 4326 2671 4378
rect 5318 4326 5370 4378
rect 5382 4326 5434 4378
rect 5446 4326 5498 4378
rect 5510 4326 5562 4378
rect 8208 4326 8260 4378
rect 8272 4326 8324 4378
rect 8336 4326 8388 4378
rect 8400 4326 8452 4378
rect 5632 4156 5684 4208
rect 5816 4088 5868 4140
rect 8944 4088 8996 4140
rect 4252 4020 4304 4072
rect 7932 4020 7984 4072
rect 2872 3952 2924 4004
rect 8024 3884 8076 3936
rect 3872 3782 3924 3834
rect 3936 3782 3988 3834
rect 4000 3782 4052 3834
rect 4064 3782 4116 3834
rect 6763 3782 6815 3834
rect 6827 3782 6879 3834
rect 6891 3782 6943 3834
rect 6955 3782 7007 3834
rect 2427 3238 2479 3290
rect 2491 3238 2543 3290
rect 2555 3238 2607 3290
rect 2619 3238 2671 3290
rect 5318 3238 5370 3290
rect 5382 3238 5434 3290
rect 5446 3238 5498 3290
rect 5510 3238 5562 3290
rect 8208 3238 8260 3290
rect 8272 3238 8324 3290
rect 8336 3238 8388 3290
rect 8400 3238 8452 3290
rect 1768 3136 1820 3188
rect 5724 3136 5776 3188
rect 3872 2694 3924 2746
rect 3936 2694 3988 2746
rect 4000 2694 4052 2746
rect 4064 2694 4116 2746
rect 6763 2694 6815 2746
rect 6827 2694 6879 2746
rect 6891 2694 6943 2746
rect 6955 2694 7007 2746
rect 2427 2150 2479 2202
rect 2491 2150 2543 2202
rect 2555 2150 2607 2202
rect 2619 2150 2671 2202
rect 5318 2150 5370 2202
rect 5382 2150 5434 2202
rect 5446 2150 5498 2202
rect 5510 2150 5562 2202
rect 8208 2150 8260 2202
rect 8272 2150 8324 2202
rect 8336 2150 8388 2202
rect 8400 2150 8452 2202
<< metal2 >>
rect 2686 23680 2742 24480
rect 8114 23680 8170 24480
rect 2700 21978 2728 23680
rect 6642 23488 6698 23497
rect 6642 23423 6698 23432
rect 3846 22332 4142 22352
rect 3902 22330 3926 22332
rect 3982 22330 4006 22332
rect 4062 22330 4086 22332
rect 3924 22278 3926 22330
rect 3988 22278 4000 22330
rect 4062 22278 4064 22330
rect 3902 22276 3926 22278
rect 3982 22276 4006 22278
rect 4062 22276 4086 22278
rect 3846 22256 4142 22276
rect 2332 21950 2728 21978
rect 2332 20058 2360 21950
rect 2401 21788 2697 21808
rect 2457 21786 2481 21788
rect 2537 21786 2561 21788
rect 2617 21786 2641 21788
rect 2479 21734 2481 21786
rect 2543 21734 2555 21786
rect 2617 21734 2619 21786
rect 2457 21732 2481 21734
rect 2537 21732 2561 21734
rect 2617 21732 2641 21734
rect 2401 21712 2697 21732
rect 5292 21788 5588 21808
rect 5348 21786 5372 21788
rect 5428 21786 5452 21788
rect 5508 21786 5532 21788
rect 5370 21734 5372 21786
rect 5434 21734 5446 21786
rect 5508 21734 5510 21786
rect 5348 21732 5372 21734
rect 5428 21732 5452 21734
rect 5508 21732 5532 21734
rect 5292 21712 5588 21732
rect 3846 21244 4142 21264
rect 3902 21242 3926 21244
rect 3982 21242 4006 21244
rect 4062 21242 4086 21244
rect 3924 21190 3926 21242
rect 3988 21190 4000 21242
rect 4062 21190 4064 21242
rect 3902 21188 3926 21190
rect 3982 21188 4006 21190
rect 4062 21188 4086 21190
rect 3846 21168 4142 21188
rect 2401 20700 2697 20720
rect 2457 20698 2481 20700
rect 2537 20698 2561 20700
rect 2617 20698 2641 20700
rect 2479 20646 2481 20698
rect 2543 20646 2555 20698
rect 2617 20646 2619 20698
rect 2457 20644 2481 20646
rect 2537 20644 2561 20646
rect 2617 20644 2641 20646
rect 2401 20624 2697 20644
rect 5292 20700 5588 20720
rect 5348 20698 5372 20700
rect 5428 20698 5452 20700
rect 5508 20698 5532 20700
rect 5370 20646 5372 20698
rect 5434 20646 5446 20698
rect 5508 20646 5510 20698
rect 5348 20644 5372 20646
rect 5428 20644 5452 20646
rect 5508 20644 5532 20646
rect 5292 20624 5588 20644
rect 3422 20496 3478 20505
rect 3422 20431 3478 20440
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2401 19612 2697 19632
rect 2457 19610 2481 19612
rect 2537 19610 2561 19612
rect 2617 19610 2641 19612
rect 2479 19558 2481 19610
rect 2543 19558 2555 19610
rect 2617 19558 2619 19610
rect 2457 19556 2481 19558
rect 2537 19556 2561 19558
rect 2617 19556 2641 19558
rect 2401 19536 2697 19556
rect 2401 18524 2697 18544
rect 2457 18522 2481 18524
rect 2537 18522 2561 18524
rect 2617 18522 2641 18524
rect 2479 18470 2481 18522
rect 2543 18470 2555 18522
rect 2617 18470 2619 18522
rect 2457 18468 2481 18470
rect 2537 18468 2561 18470
rect 2617 18468 2641 18470
rect 2401 18448 2697 18468
rect 2401 17436 2697 17456
rect 2457 17434 2481 17436
rect 2537 17434 2561 17436
rect 2617 17434 2641 17436
rect 2479 17382 2481 17434
rect 2543 17382 2555 17434
rect 2617 17382 2619 17434
rect 2457 17380 2481 17382
rect 2537 17380 2561 17382
rect 2617 17380 2641 17382
rect 2401 17360 2697 17380
rect 2401 16348 2697 16368
rect 2457 16346 2481 16348
rect 2537 16346 2561 16348
rect 2617 16346 2641 16348
rect 2479 16294 2481 16346
rect 2543 16294 2555 16346
rect 2617 16294 2619 16346
rect 2457 16292 2481 16294
rect 2537 16292 2561 16294
rect 2617 16292 2641 16294
rect 2401 16272 2697 16292
rect 2401 15260 2697 15280
rect 2457 15258 2481 15260
rect 2537 15258 2561 15260
rect 2617 15258 2641 15260
rect 2479 15206 2481 15258
rect 2543 15206 2555 15258
rect 2617 15206 2619 15258
rect 2457 15204 2481 15206
rect 2537 15204 2561 15206
rect 2617 15204 2641 15206
rect 2401 15184 2697 15204
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14482 1440 14894
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 14074 1440 14418
rect 2401 14172 2697 14192
rect 2457 14170 2481 14172
rect 2537 14170 2561 14172
rect 2617 14170 2641 14172
rect 2479 14118 2481 14170
rect 2543 14118 2555 14170
rect 2617 14118 2619 14170
rect 2457 14116 2481 14118
rect 2537 14116 2561 14118
rect 2617 14116 2641 14118
rect 2401 14096 2697 14116
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 2401 13084 2697 13104
rect 2457 13082 2481 13084
rect 2537 13082 2561 13084
rect 2617 13082 2641 13084
rect 2479 13030 2481 13082
rect 2543 13030 2555 13082
rect 2617 13030 2619 13082
rect 2457 13028 2481 13030
rect 2537 13028 2561 13030
rect 2617 13028 2641 13030
rect 2401 13008 2697 13028
rect 2870 12336 2926 12345
rect 2870 12271 2926 12280
rect 2401 11996 2697 12016
rect 2457 11994 2481 11996
rect 2537 11994 2561 11996
rect 2617 11994 2641 11996
rect 2479 11942 2481 11994
rect 2543 11942 2555 11994
rect 2617 11942 2619 11994
rect 2457 11940 2481 11942
rect 2537 11940 2561 11942
rect 2617 11940 2641 11942
rect 2401 11920 2697 11940
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2401 10908 2697 10928
rect 2457 10906 2481 10908
rect 2537 10906 2561 10908
rect 2617 10906 2641 10908
rect 2479 10854 2481 10906
rect 2543 10854 2555 10906
rect 2617 10854 2619 10906
rect 2457 10852 2481 10854
rect 2537 10852 2561 10854
rect 2617 10852 2641 10854
rect 2401 10832 2697 10852
rect 2401 9820 2697 9840
rect 2457 9818 2481 9820
rect 2537 9818 2561 9820
rect 2617 9818 2641 9820
rect 2479 9766 2481 9818
rect 2543 9766 2555 9818
rect 2617 9766 2619 9818
rect 2457 9764 2481 9766
rect 2537 9764 2561 9766
rect 2617 9764 2641 9766
rect 2401 9744 2697 9764
rect 2401 8732 2697 8752
rect 2457 8730 2481 8732
rect 2537 8730 2561 8732
rect 2617 8730 2641 8732
rect 2479 8678 2481 8730
rect 2543 8678 2555 8730
rect 2617 8678 2619 8730
rect 2457 8676 2481 8678
rect 2537 8676 2561 8678
rect 2617 8676 2641 8678
rect 2401 8656 2697 8676
rect 2792 8090 2820 11018
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7206 2268 7890
rect 2401 7644 2697 7664
rect 2457 7642 2481 7644
rect 2537 7642 2561 7644
rect 2617 7642 2641 7644
rect 2479 7590 2481 7642
rect 2543 7590 2555 7642
rect 2617 7590 2619 7642
rect 2457 7588 2481 7590
rect 2537 7588 2561 7590
rect 2617 7588 2641 7590
rect 2401 7568 2697 7588
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2401 6556 2697 6576
rect 2457 6554 2481 6556
rect 2537 6554 2561 6556
rect 2617 6554 2641 6556
rect 2479 6502 2481 6554
rect 2543 6502 2555 6554
rect 2617 6502 2619 6554
rect 2457 6500 2481 6502
rect 2537 6500 2561 6502
rect 2617 6500 2641 6502
rect 2401 6480 2697 6500
rect 2401 5468 2697 5488
rect 2457 5466 2481 5468
rect 2537 5466 2561 5468
rect 2617 5466 2641 5468
rect 2479 5414 2481 5466
rect 2543 5414 2555 5466
rect 2617 5414 2619 5466
rect 2457 5412 2481 5414
rect 2537 5412 2561 5414
rect 2617 5412 2641 5414
rect 2401 5392 2697 5412
rect 2401 4380 2697 4400
rect 2457 4378 2481 4380
rect 2537 4378 2561 4380
rect 2617 4378 2641 4380
rect 2479 4326 2481 4378
rect 2543 4326 2555 4378
rect 2617 4326 2619 4378
rect 2457 4324 2481 4326
rect 2537 4324 2561 4326
rect 2617 4324 2641 4326
rect 2401 4304 2697 4324
rect 2884 4010 2912 12271
rect 3436 11762 3464 20431
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 3846 20156 4142 20176
rect 3902 20154 3926 20156
rect 3982 20154 4006 20156
rect 4062 20154 4086 20156
rect 3924 20102 3926 20154
rect 3988 20102 4000 20154
rect 4062 20102 4064 20154
rect 3902 20100 3926 20102
rect 3982 20100 4006 20102
rect 4062 20100 4086 20102
rect 3846 20080 4142 20100
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 3846 19068 4142 19088
rect 3902 19066 3926 19068
rect 3982 19066 4006 19068
rect 4062 19066 4086 19068
rect 3924 19014 3926 19066
rect 3988 19014 4000 19066
rect 4062 19014 4064 19066
rect 3902 19012 3926 19014
rect 3982 19012 4006 19014
rect 4062 19012 4086 19014
rect 3846 18992 4142 19012
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18154 4384 18566
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 3846 17980 4142 18000
rect 3902 17978 3926 17980
rect 3982 17978 4006 17980
rect 4062 17978 4086 17980
rect 3924 17926 3926 17978
rect 3988 17926 4000 17978
rect 4062 17926 4064 17978
rect 3902 17924 3926 17926
rect 3982 17924 4006 17926
rect 4062 17924 4086 17926
rect 3846 17904 4142 17924
rect 3846 16892 4142 16912
rect 3902 16890 3926 16892
rect 3982 16890 4006 16892
rect 4062 16890 4086 16892
rect 3924 16838 3926 16890
rect 3988 16838 4000 16890
rect 4062 16838 4064 16890
rect 3902 16836 3926 16838
rect 3982 16836 4006 16838
rect 4062 16836 4086 16838
rect 3846 16816 4142 16836
rect 3846 15804 4142 15824
rect 3902 15802 3926 15804
rect 3982 15802 4006 15804
rect 4062 15802 4086 15804
rect 3924 15750 3926 15802
rect 3988 15750 4000 15802
rect 4062 15750 4064 15802
rect 3902 15748 3926 15750
rect 3982 15748 4006 15750
rect 4062 15748 4086 15750
rect 3846 15728 4142 15748
rect 3846 14716 4142 14736
rect 3902 14714 3926 14716
rect 3982 14714 4006 14716
rect 4062 14714 4086 14716
rect 3924 14662 3926 14714
rect 3988 14662 4000 14714
rect 4062 14662 4064 14714
rect 3902 14660 3926 14662
rect 3982 14660 4006 14662
rect 4062 14660 4086 14662
rect 3846 14640 4142 14660
rect 3846 13628 4142 13648
rect 3902 13626 3926 13628
rect 3982 13626 4006 13628
rect 4062 13626 4086 13628
rect 3924 13574 3926 13626
rect 3988 13574 4000 13626
rect 4062 13574 4064 13626
rect 3902 13572 3926 13574
rect 3982 13572 4006 13574
rect 4062 13572 4086 13574
rect 3846 13552 4142 13572
rect 3846 12540 4142 12560
rect 3902 12538 3926 12540
rect 3982 12538 4006 12540
rect 4062 12538 4086 12540
rect 3924 12486 3926 12538
rect 3988 12486 4000 12538
rect 4062 12486 4064 12538
rect 3902 12484 3926 12486
rect 3982 12484 4006 12486
rect 4062 12484 4086 12486
rect 3846 12464 4142 12484
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3846 11452 4142 11472
rect 3902 11450 3926 11452
rect 3982 11450 4006 11452
rect 4062 11450 4086 11452
rect 3924 11398 3926 11450
rect 3988 11398 4000 11450
rect 4062 11398 4064 11450
rect 3902 11396 3926 11398
rect 3982 11396 4006 11398
rect 4062 11396 4086 11398
rect 3846 11376 4142 11396
rect 3846 10364 4142 10384
rect 3902 10362 3926 10364
rect 3982 10362 4006 10364
rect 4062 10362 4086 10364
rect 3924 10310 3926 10362
rect 3988 10310 4000 10362
rect 4062 10310 4064 10362
rect 3902 10308 3926 10310
rect 3982 10308 4006 10310
rect 4062 10308 4086 10310
rect 3846 10288 4142 10308
rect 3846 9276 4142 9296
rect 3902 9274 3926 9276
rect 3982 9274 4006 9276
rect 4062 9274 4086 9276
rect 3924 9222 3926 9274
rect 3988 9222 4000 9274
rect 4062 9222 4064 9274
rect 3902 9220 3926 9222
rect 3982 9220 4006 9222
rect 4062 9220 4086 9222
rect 3846 9200 4142 9220
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 4185 3372 8774
rect 3846 8188 4142 8208
rect 3902 8186 3926 8188
rect 3982 8186 4006 8188
rect 4062 8186 4086 8188
rect 3924 8134 3926 8186
rect 3988 8134 4000 8186
rect 4062 8134 4064 8186
rect 3902 8132 3926 8134
rect 3982 8132 4006 8134
rect 4062 8132 4086 8134
rect 3846 8112 4142 8132
rect 3846 7100 4142 7120
rect 3902 7098 3926 7100
rect 3982 7098 4006 7100
rect 4062 7098 4086 7100
rect 3924 7046 3926 7098
rect 3988 7046 4000 7098
rect 4062 7046 4064 7098
rect 3902 7044 3926 7046
rect 3982 7044 4006 7046
rect 4062 7044 4086 7046
rect 3846 7024 4142 7044
rect 3846 6012 4142 6032
rect 3902 6010 3926 6012
rect 3982 6010 4006 6012
rect 4062 6010 4086 6012
rect 3924 5958 3926 6010
rect 3988 5958 4000 6010
rect 4062 5958 4064 6010
rect 3902 5956 3926 5958
rect 3982 5956 4006 5958
rect 4062 5956 4086 5958
rect 3846 5936 4142 5956
rect 4448 5370 4476 19314
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6254 4936 7142
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4908 5370 4936 6190
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 5166 4936 5306
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 3846 4924 4142 4944
rect 3902 4922 3926 4924
rect 3982 4922 4006 4924
rect 4062 4922 4086 4924
rect 3924 4870 3926 4922
rect 3988 4870 4000 4922
rect 4062 4870 4064 4922
rect 3902 4868 3926 4870
rect 3982 4868 4006 4870
rect 4062 4868 4086 4870
rect 3846 4848 4142 4868
rect 3330 4176 3386 4185
rect 3330 4111 3386 4120
rect 4264 4078 4292 5102
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 3846 3836 4142 3856
rect 3902 3834 3926 3836
rect 3982 3834 4006 3836
rect 4062 3834 4086 3836
rect 3924 3782 3926 3834
rect 3988 3782 4000 3834
rect 4062 3782 4064 3834
rect 3902 3780 3926 3782
rect 3982 3780 4006 3782
rect 4062 3780 4086 3782
rect 3846 3760 4142 3780
rect 2401 3292 2697 3312
rect 2457 3290 2481 3292
rect 2537 3290 2561 3292
rect 2617 3290 2641 3292
rect 2479 3238 2481 3290
rect 2543 3238 2555 3290
rect 2617 3238 2619 3290
rect 2457 3236 2481 3238
rect 2537 3236 2561 3238
rect 2617 3236 2641 3238
rect 2401 3216 2697 3236
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1780 800 1808 3130
rect 3846 2748 4142 2768
rect 3902 2746 3926 2748
rect 3982 2746 4006 2748
rect 4062 2746 4086 2748
rect 3924 2694 3926 2746
rect 3988 2694 4000 2746
rect 4062 2694 4064 2746
rect 3902 2692 3926 2694
rect 3982 2692 4006 2694
rect 4062 2692 4086 2694
rect 3846 2672 4142 2692
rect 2401 2204 2697 2224
rect 2457 2202 2481 2204
rect 2537 2202 2561 2204
rect 2617 2202 2641 2204
rect 2479 2150 2481 2202
rect 2543 2150 2555 2202
rect 2617 2150 2619 2202
rect 2457 2148 2481 2150
rect 2537 2148 2561 2150
rect 2617 2148 2641 2150
rect 2401 2128 2697 2148
rect 5092 921 5120 18022
rect 5184 1986 5212 20198
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 5630 19816 5686 19825
rect 5630 19751 5686 19760
rect 5292 19612 5588 19632
rect 5348 19610 5372 19612
rect 5428 19610 5452 19612
rect 5508 19610 5532 19612
rect 5370 19558 5372 19610
rect 5434 19558 5446 19610
rect 5508 19558 5510 19610
rect 5348 19556 5372 19558
rect 5428 19556 5452 19558
rect 5508 19556 5532 19558
rect 5292 19536 5588 19556
rect 5644 19378 5672 19751
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5292 18524 5588 18544
rect 5348 18522 5372 18524
rect 5428 18522 5452 18524
rect 5508 18522 5532 18524
rect 5370 18470 5372 18522
rect 5434 18470 5446 18522
rect 5508 18470 5510 18522
rect 5348 18468 5372 18470
rect 5428 18468 5452 18470
rect 5508 18468 5532 18470
rect 5292 18448 5588 18468
rect 5292 17436 5588 17456
rect 5348 17434 5372 17436
rect 5428 17434 5452 17436
rect 5508 17434 5532 17436
rect 5370 17382 5372 17434
rect 5434 17382 5446 17434
rect 5508 17382 5510 17434
rect 5348 17380 5372 17382
rect 5428 17380 5452 17382
rect 5508 17380 5532 17382
rect 5292 17360 5588 17380
rect 5292 16348 5588 16368
rect 5348 16346 5372 16348
rect 5428 16346 5452 16348
rect 5508 16346 5532 16348
rect 5370 16294 5372 16346
rect 5434 16294 5446 16346
rect 5508 16294 5510 16346
rect 5348 16292 5372 16294
rect 5428 16292 5452 16294
rect 5508 16292 5532 16294
rect 5292 16272 5588 16292
rect 5292 15260 5588 15280
rect 5348 15258 5372 15260
rect 5428 15258 5452 15260
rect 5508 15258 5532 15260
rect 5370 15206 5372 15258
rect 5434 15206 5446 15258
rect 5508 15206 5510 15258
rect 5348 15204 5372 15206
rect 5428 15204 5452 15206
rect 5508 15204 5532 15206
rect 5292 15184 5588 15204
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5292 14172 5588 14192
rect 5348 14170 5372 14172
rect 5428 14170 5452 14172
rect 5508 14170 5532 14172
rect 5370 14118 5372 14170
rect 5434 14118 5446 14170
rect 5508 14118 5510 14170
rect 5348 14116 5372 14118
rect 5428 14116 5452 14118
rect 5508 14116 5532 14118
rect 5292 14096 5588 14116
rect 5644 13977 5672 14214
rect 5630 13968 5686 13977
rect 5630 13903 5686 13912
rect 5292 13084 5588 13104
rect 5348 13082 5372 13084
rect 5428 13082 5452 13084
rect 5508 13082 5532 13084
rect 5370 13030 5372 13082
rect 5434 13030 5446 13082
rect 5508 13030 5510 13082
rect 5348 13028 5372 13030
rect 5428 13028 5452 13030
rect 5508 13028 5532 13030
rect 5292 13008 5588 13028
rect 5630 12200 5686 12209
rect 5630 12135 5686 12144
rect 5292 11996 5588 12016
rect 5348 11994 5372 11996
rect 5428 11994 5452 11996
rect 5508 11994 5532 11996
rect 5370 11942 5372 11994
rect 5434 11942 5446 11994
rect 5508 11942 5510 11994
rect 5348 11940 5372 11942
rect 5428 11940 5452 11942
rect 5508 11940 5532 11942
rect 5292 11920 5588 11940
rect 5644 11082 5672 12135
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5292 10908 5588 10928
rect 5348 10906 5372 10908
rect 5428 10906 5452 10908
rect 5508 10906 5532 10908
rect 5370 10854 5372 10906
rect 5434 10854 5446 10906
rect 5508 10854 5510 10906
rect 5348 10852 5372 10854
rect 5428 10852 5452 10854
rect 5508 10852 5532 10854
rect 5292 10832 5588 10852
rect 5292 9820 5588 9840
rect 5348 9818 5372 9820
rect 5428 9818 5452 9820
rect 5508 9818 5532 9820
rect 5370 9766 5372 9818
rect 5434 9766 5446 9818
rect 5508 9766 5510 9818
rect 5348 9764 5372 9766
rect 5428 9764 5452 9766
rect 5508 9764 5532 9766
rect 5292 9744 5588 9764
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5292 8732 5588 8752
rect 5348 8730 5372 8732
rect 5428 8730 5452 8732
rect 5508 8730 5532 8732
rect 5370 8678 5372 8730
rect 5434 8678 5446 8730
rect 5508 8678 5510 8730
rect 5348 8676 5372 8678
rect 5428 8676 5452 8678
rect 5508 8676 5532 8678
rect 5292 8656 5588 8676
rect 5828 8634 5856 9046
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5828 8022 5856 8570
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5292 7644 5588 7664
rect 5348 7642 5372 7644
rect 5428 7642 5452 7644
rect 5508 7642 5532 7644
rect 5370 7590 5372 7642
rect 5434 7590 5446 7642
rect 5508 7590 5510 7642
rect 5348 7588 5372 7590
rect 5428 7588 5452 7590
rect 5508 7588 5532 7590
rect 5292 7568 5588 7588
rect 5292 6556 5588 6576
rect 5348 6554 5372 6556
rect 5428 6554 5452 6556
rect 5508 6554 5532 6556
rect 5370 6502 5372 6554
rect 5434 6502 5446 6554
rect 5508 6502 5510 6554
rect 5348 6500 5372 6502
rect 5428 6500 5452 6502
rect 5508 6500 5532 6502
rect 5292 6480 5588 6500
rect 5292 5468 5588 5488
rect 5348 5466 5372 5468
rect 5428 5466 5452 5468
rect 5508 5466 5532 5468
rect 5370 5414 5372 5466
rect 5434 5414 5446 5466
rect 5508 5414 5510 5466
rect 5348 5412 5372 5414
rect 5428 5412 5452 5414
rect 5508 5412 5532 5414
rect 5292 5392 5588 5412
rect 5630 4584 5686 4593
rect 5630 4519 5686 4528
rect 5292 4380 5588 4400
rect 5348 4378 5372 4380
rect 5428 4378 5452 4380
rect 5508 4378 5532 4380
rect 5370 4326 5372 4378
rect 5434 4326 5446 4378
rect 5508 4326 5510 4378
rect 5348 4324 5372 4326
rect 5428 4324 5452 4326
rect 5508 4324 5532 4326
rect 5292 4304 5588 4324
rect 5644 4214 5672 4519
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5292 3292 5588 3312
rect 5348 3290 5372 3292
rect 5428 3290 5452 3292
rect 5508 3290 5532 3292
rect 5370 3238 5372 3290
rect 5434 3238 5446 3290
rect 5508 3238 5510 3290
rect 5348 3236 5372 3238
rect 5428 3236 5452 3238
rect 5508 3236 5532 3238
rect 5292 3216 5588 3236
rect 5736 3194 5764 7686
rect 5828 7546 5856 7958
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5828 4146 5856 7482
rect 6196 6769 6224 15030
rect 6288 14074 6316 19994
rect 6552 18148 6604 18154
rect 6552 18090 6604 18096
rect 6458 15600 6514 15609
rect 6458 15535 6514 15544
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6380 10606 6408 13806
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 9110 6408 10542
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6182 6760 6238 6769
rect 6182 6695 6238 6704
rect 6472 5914 6500 15535
rect 6564 14618 6592 18090
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6564 13870 6592 14554
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 10577 6592 12582
rect 6656 11234 6684 23423
rect 6737 22332 7033 22352
rect 6793 22330 6817 22332
rect 6873 22330 6897 22332
rect 6953 22330 6977 22332
rect 6815 22278 6817 22330
rect 6879 22278 6891 22330
rect 6953 22278 6955 22330
rect 6793 22276 6817 22278
rect 6873 22276 6897 22278
rect 6953 22276 6977 22278
rect 6737 22256 7033 22276
rect 8128 21978 8156 23680
rect 8036 21950 8156 21978
rect 7102 21584 7158 21593
rect 7102 21519 7158 21528
rect 6737 21244 7033 21264
rect 6793 21242 6817 21244
rect 6873 21242 6897 21244
rect 6953 21242 6977 21244
rect 6815 21190 6817 21242
rect 6879 21190 6891 21242
rect 6953 21190 6955 21242
rect 6793 21188 6817 21190
rect 6873 21188 6897 21190
rect 6953 21188 6977 21190
rect 6737 21168 7033 21188
rect 6737 20156 7033 20176
rect 6793 20154 6817 20156
rect 6873 20154 6897 20156
rect 6953 20154 6977 20156
rect 6815 20102 6817 20154
rect 6879 20102 6891 20154
rect 6953 20102 6955 20154
rect 6793 20100 6817 20102
rect 6873 20100 6897 20102
rect 6953 20100 6977 20102
rect 6737 20080 7033 20100
rect 6737 19068 7033 19088
rect 6793 19066 6817 19068
rect 6873 19066 6897 19068
rect 6953 19066 6977 19068
rect 6815 19014 6817 19066
rect 6879 19014 6891 19066
rect 6953 19014 6955 19066
rect 6793 19012 6817 19014
rect 6873 19012 6897 19014
rect 6953 19012 6977 19014
rect 6737 18992 7033 19012
rect 6737 17980 7033 18000
rect 6793 17978 6817 17980
rect 6873 17978 6897 17980
rect 6953 17978 6977 17980
rect 6815 17926 6817 17978
rect 6879 17926 6891 17978
rect 6953 17926 6955 17978
rect 6793 17924 6817 17926
rect 6873 17924 6897 17926
rect 6953 17924 6977 17926
rect 6737 17904 7033 17924
rect 6737 16892 7033 16912
rect 6793 16890 6817 16892
rect 6873 16890 6897 16892
rect 6953 16890 6977 16892
rect 6815 16838 6817 16890
rect 6879 16838 6891 16890
rect 6953 16838 6955 16890
rect 6793 16836 6817 16838
rect 6873 16836 6897 16838
rect 6953 16836 6977 16838
rect 6737 16816 7033 16836
rect 6737 15804 7033 15824
rect 6793 15802 6817 15804
rect 6873 15802 6897 15804
rect 6953 15802 6977 15804
rect 6815 15750 6817 15802
rect 6879 15750 6891 15802
rect 6953 15750 6955 15802
rect 6793 15748 6817 15750
rect 6873 15748 6897 15750
rect 6953 15748 6977 15750
rect 6737 15728 7033 15748
rect 6737 14716 7033 14736
rect 6793 14714 6817 14716
rect 6873 14714 6897 14716
rect 6953 14714 6977 14716
rect 6815 14662 6817 14714
rect 6879 14662 6891 14714
rect 6953 14662 6955 14714
rect 6793 14660 6817 14662
rect 6873 14660 6897 14662
rect 6953 14660 6977 14662
rect 6737 14640 7033 14660
rect 6737 13628 7033 13648
rect 6793 13626 6817 13628
rect 6873 13626 6897 13628
rect 6953 13626 6977 13628
rect 6815 13574 6817 13626
rect 6879 13574 6891 13626
rect 6953 13574 6955 13626
rect 6793 13572 6817 13574
rect 6873 13572 6897 13574
rect 6953 13572 6977 13574
rect 6737 13552 7033 13572
rect 6737 12540 7033 12560
rect 6793 12538 6817 12540
rect 6873 12538 6897 12540
rect 6953 12538 6977 12540
rect 6815 12486 6817 12538
rect 6879 12486 6891 12538
rect 6953 12486 6955 12538
rect 6793 12484 6817 12486
rect 6873 12484 6897 12486
rect 6953 12484 6977 12486
rect 6737 12464 7033 12484
rect 6737 11452 7033 11472
rect 6793 11450 6817 11452
rect 6873 11450 6897 11452
rect 6953 11450 6977 11452
rect 6815 11398 6817 11450
rect 6879 11398 6891 11450
rect 6953 11398 6955 11450
rect 6793 11396 6817 11398
rect 6873 11396 6897 11398
rect 6953 11396 6977 11398
rect 6737 11376 7033 11396
rect 6656 11206 6776 11234
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6550 10568 6606 10577
rect 6550 10503 6606 10512
rect 6656 8401 6684 11018
rect 6748 10810 6776 11206
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6737 10364 7033 10384
rect 6793 10362 6817 10364
rect 6873 10362 6897 10364
rect 6953 10362 6977 10364
rect 6815 10310 6817 10362
rect 6879 10310 6891 10362
rect 6953 10310 6955 10362
rect 6793 10308 6817 10310
rect 6873 10308 6897 10310
rect 6953 10308 6977 10310
rect 6737 10288 7033 10308
rect 6737 9276 7033 9296
rect 6793 9274 6817 9276
rect 6873 9274 6897 9276
rect 6953 9274 6977 9276
rect 6815 9222 6817 9274
rect 6879 9222 6891 9274
rect 6953 9222 6955 9274
rect 6793 9220 6817 9222
rect 6873 9220 6897 9222
rect 6953 9220 6977 9222
rect 6737 9200 7033 9220
rect 6642 8392 6698 8401
rect 6642 8327 6698 8336
rect 6737 8188 7033 8208
rect 6793 8186 6817 8188
rect 6873 8186 6897 8188
rect 6953 8186 6977 8188
rect 6815 8134 6817 8186
rect 6879 8134 6891 8186
rect 6953 8134 6955 8186
rect 6793 8132 6817 8134
rect 6873 8132 6897 8134
rect 6953 8132 6977 8134
rect 6737 8112 7033 8132
rect 6737 7100 7033 7120
rect 6793 7098 6817 7100
rect 6873 7098 6897 7100
rect 6953 7098 6977 7100
rect 6815 7046 6817 7098
rect 6879 7046 6891 7098
rect 6953 7046 6955 7098
rect 6793 7044 6817 7046
rect 6873 7044 6897 7046
rect 6953 7044 6977 7046
rect 6737 7024 7033 7044
rect 7116 6458 7144 21519
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 18222 7972 20198
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7392 14822 7420 18158
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 12646 7420 14758
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 11898 7420 12582
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7392 11218 7420 11834
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7392 10470 7420 11154
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7392 6254 7420 10406
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 6737 6012 7033 6032
rect 6793 6010 6817 6012
rect 6873 6010 6897 6012
rect 6953 6010 6977 6012
rect 6815 5958 6817 6010
rect 6879 5958 6891 6010
rect 6953 5958 6955 6010
rect 6793 5956 6817 5958
rect 6873 5956 6897 5958
rect 6953 5956 6977 5958
rect 6737 5936 7033 5956
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 7944 5778 7972 6054
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7944 5030 7972 5714
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 6737 4924 7033 4944
rect 6793 4922 6817 4924
rect 6873 4922 6897 4924
rect 6953 4922 6977 4924
rect 6815 4870 6817 4922
rect 6879 4870 6891 4922
rect 6953 4870 6955 4922
rect 6793 4868 6817 4870
rect 6873 4868 6897 4870
rect 6953 4868 6977 4870
rect 6737 4848 7033 4868
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 7944 4078 7972 4966
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8036 3942 8064 21950
rect 8182 21788 8478 21808
rect 8238 21786 8262 21788
rect 8318 21786 8342 21788
rect 8398 21786 8422 21788
rect 8260 21734 8262 21786
rect 8324 21734 8336 21786
rect 8398 21734 8400 21786
rect 8238 21732 8262 21734
rect 8318 21732 8342 21734
rect 8398 21732 8422 21734
rect 8182 21712 8478 21732
rect 8182 20700 8478 20720
rect 8238 20698 8262 20700
rect 8318 20698 8342 20700
rect 8398 20698 8422 20700
rect 8260 20646 8262 20698
rect 8324 20646 8336 20698
rect 8398 20646 8400 20698
rect 8238 20644 8262 20646
rect 8318 20644 8342 20646
rect 8398 20644 8422 20646
rect 8182 20624 8478 20644
rect 8182 19612 8478 19632
rect 8238 19610 8262 19612
rect 8318 19610 8342 19612
rect 8398 19610 8422 19612
rect 8260 19558 8262 19610
rect 8324 19558 8336 19610
rect 8398 19558 8400 19610
rect 8238 19556 8262 19558
rect 8318 19556 8342 19558
rect 8398 19556 8422 19558
rect 8182 19536 8478 19556
rect 8182 18524 8478 18544
rect 8238 18522 8262 18524
rect 8318 18522 8342 18524
rect 8398 18522 8422 18524
rect 8260 18470 8262 18522
rect 8324 18470 8336 18522
rect 8398 18470 8400 18522
rect 8238 18468 8262 18470
rect 8318 18468 8342 18470
rect 8398 18468 8422 18470
rect 8182 18448 8478 18468
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17785 8248 18022
rect 8206 17776 8262 17785
rect 8206 17711 8262 17720
rect 8182 17436 8478 17456
rect 8238 17434 8262 17436
rect 8318 17434 8342 17436
rect 8398 17434 8422 17436
rect 8260 17382 8262 17434
rect 8324 17382 8336 17434
rect 8398 17382 8400 17434
rect 8238 17380 8262 17382
rect 8318 17380 8342 17382
rect 8398 17380 8422 17382
rect 8182 17360 8478 17380
rect 8182 16348 8478 16368
rect 8238 16346 8262 16348
rect 8318 16346 8342 16348
rect 8398 16346 8422 16348
rect 8260 16294 8262 16346
rect 8324 16294 8336 16346
rect 8398 16294 8400 16346
rect 8238 16292 8262 16294
rect 8318 16292 8342 16294
rect 8398 16292 8422 16294
rect 8182 16272 8478 16292
rect 8182 15260 8478 15280
rect 8238 15258 8262 15260
rect 8318 15258 8342 15260
rect 8398 15258 8422 15260
rect 8260 15206 8262 15258
rect 8324 15206 8336 15258
rect 8398 15206 8400 15258
rect 8238 15204 8262 15206
rect 8318 15204 8342 15206
rect 8398 15204 8422 15206
rect 8182 15184 8478 15204
rect 8182 14172 8478 14192
rect 8238 14170 8262 14172
rect 8318 14170 8342 14172
rect 8398 14170 8422 14172
rect 8260 14118 8262 14170
rect 8324 14118 8336 14170
rect 8398 14118 8400 14170
rect 8238 14116 8262 14118
rect 8318 14116 8342 14118
rect 8398 14116 8422 14118
rect 8182 14096 8478 14116
rect 8182 13084 8478 13104
rect 8238 13082 8262 13084
rect 8318 13082 8342 13084
rect 8398 13082 8422 13084
rect 8260 13030 8262 13082
rect 8324 13030 8336 13082
rect 8398 13030 8400 13082
rect 8238 13028 8262 13030
rect 8318 13028 8342 13030
rect 8398 13028 8422 13030
rect 8182 13008 8478 13028
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8182 11996 8478 12016
rect 8238 11994 8262 11996
rect 8318 11994 8342 11996
rect 8398 11994 8422 11996
rect 8260 11942 8262 11994
rect 8324 11942 8336 11994
rect 8398 11942 8400 11994
rect 8238 11940 8262 11942
rect 8318 11940 8342 11942
rect 8398 11940 8422 11942
rect 8182 11920 8478 11940
rect 8182 10908 8478 10928
rect 8238 10906 8262 10908
rect 8318 10906 8342 10908
rect 8398 10906 8422 10908
rect 8260 10854 8262 10906
rect 8324 10854 8336 10906
rect 8398 10854 8400 10906
rect 8238 10852 8262 10854
rect 8318 10852 8342 10854
rect 8398 10852 8422 10854
rect 8182 10832 8478 10852
rect 8182 9820 8478 9840
rect 8238 9818 8262 9820
rect 8318 9818 8342 9820
rect 8398 9818 8422 9820
rect 8260 9766 8262 9818
rect 8324 9766 8336 9818
rect 8398 9766 8400 9818
rect 8238 9764 8262 9766
rect 8318 9764 8342 9766
rect 8398 9764 8422 9766
rect 8182 9744 8478 9764
rect 8182 8732 8478 8752
rect 8238 8730 8262 8732
rect 8318 8730 8342 8732
rect 8398 8730 8422 8732
rect 8260 8678 8262 8730
rect 8324 8678 8336 8730
rect 8398 8678 8400 8730
rect 8238 8676 8262 8678
rect 8318 8676 8342 8678
rect 8398 8676 8422 8678
rect 8182 8656 8478 8676
rect 8182 7644 8478 7664
rect 8238 7642 8262 7644
rect 8318 7642 8342 7644
rect 8398 7642 8422 7644
rect 8260 7590 8262 7642
rect 8324 7590 8336 7642
rect 8398 7590 8400 7642
rect 8238 7588 8262 7590
rect 8318 7588 8342 7590
rect 8398 7588 8422 7590
rect 8182 7568 8478 7588
rect 8182 6556 8478 6576
rect 8238 6554 8262 6556
rect 8318 6554 8342 6556
rect 8398 6554 8422 6556
rect 8260 6502 8262 6554
rect 8324 6502 8336 6554
rect 8398 6502 8400 6554
rect 8238 6500 8262 6502
rect 8318 6500 8342 6502
rect 8398 6500 8422 6502
rect 8182 6480 8478 6500
rect 8182 5468 8478 5488
rect 8238 5466 8262 5468
rect 8318 5466 8342 5468
rect 8398 5466 8422 5468
rect 8260 5414 8262 5466
rect 8324 5414 8336 5466
rect 8398 5414 8400 5466
rect 8238 5412 8262 5414
rect 8318 5412 8342 5414
rect 8398 5412 8422 5414
rect 8182 5392 8478 5412
rect 8182 4380 8478 4400
rect 8238 4378 8262 4380
rect 8318 4378 8342 4380
rect 8398 4378 8422 4380
rect 8260 4326 8262 4378
rect 8324 4326 8336 4378
rect 8398 4326 8400 4378
rect 8238 4324 8262 4326
rect 8318 4324 8342 4326
rect 8398 4324 8422 4326
rect 8182 4304 8478 4324
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 6737 3836 7033 3856
rect 6793 3834 6817 3836
rect 6873 3834 6897 3836
rect 6953 3834 6977 3836
rect 6815 3782 6817 3834
rect 6879 3782 6891 3834
rect 6953 3782 6955 3834
rect 6793 3780 6817 3782
rect 6873 3780 6897 3782
rect 6953 3780 6977 3782
rect 6737 3760 7033 3780
rect 8182 3292 8478 3312
rect 8238 3290 8262 3292
rect 8318 3290 8342 3292
rect 8398 3290 8422 3292
rect 8260 3238 8262 3290
rect 8324 3238 8336 3290
rect 8398 3238 8400 3290
rect 8238 3236 8262 3238
rect 8318 3236 8342 3238
rect 8398 3236 8422 3238
rect 8182 3216 8478 3236
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 6737 2748 7033 2768
rect 6793 2746 6817 2748
rect 6873 2746 6897 2748
rect 6953 2746 6977 2748
rect 6815 2694 6817 2746
rect 6879 2694 6891 2746
rect 6953 2694 6955 2746
rect 6793 2692 6817 2694
rect 6873 2692 6897 2694
rect 6953 2692 6977 2694
rect 6737 2672 7033 2692
rect 8588 2689 8616 12582
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8574 2680 8630 2689
rect 8574 2615 8630 2624
rect 5292 2204 5588 2224
rect 5348 2202 5372 2204
rect 5428 2202 5452 2204
rect 5508 2202 5532 2204
rect 5370 2150 5372 2202
rect 5434 2150 5446 2202
rect 5508 2150 5510 2202
rect 5348 2148 5372 2150
rect 5428 2148 5452 2150
rect 5508 2148 5532 2150
rect 5292 2128 5588 2148
rect 8182 2204 8478 2224
rect 8238 2202 8262 2204
rect 8318 2202 8342 2204
rect 8398 2202 8422 2204
rect 8260 2150 8262 2202
rect 8324 2150 8336 2202
rect 8398 2150 8400 2202
rect 8238 2148 8262 2150
rect 8318 2148 8342 2150
rect 8398 2148 8422 2150
rect 8182 2128 8478 2148
rect 5184 1958 5396 1986
rect 5078 912 5134 921
rect 5078 847 5134 856
rect 5368 800 5396 1958
rect 8956 800 8984 4082
rect 1766 0 1822 800
rect 5354 0 5410 800
rect 8942 0 8998 800
<< via2 >>
rect 6642 23432 6698 23488
rect 3846 22330 3902 22332
rect 3926 22330 3982 22332
rect 4006 22330 4062 22332
rect 4086 22330 4142 22332
rect 3846 22278 3872 22330
rect 3872 22278 3902 22330
rect 3926 22278 3936 22330
rect 3936 22278 3982 22330
rect 4006 22278 4052 22330
rect 4052 22278 4062 22330
rect 4086 22278 4116 22330
rect 4116 22278 4142 22330
rect 3846 22276 3902 22278
rect 3926 22276 3982 22278
rect 4006 22276 4062 22278
rect 4086 22276 4142 22278
rect 2401 21786 2457 21788
rect 2481 21786 2537 21788
rect 2561 21786 2617 21788
rect 2641 21786 2697 21788
rect 2401 21734 2427 21786
rect 2427 21734 2457 21786
rect 2481 21734 2491 21786
rect 2491 21734 2537 21786
rect 2561 21734 2607 21786
rect 2607 21734 2617 21786
rect 2641 21734 2671 21786
rect 2671 21734 2697 21786
rect 2401 21732 2457 21734
rect 2481 21732 2537 21734
rect 2561 21732 2617 21734
rect 2641 21732 2697 21734
rect 5292 21786 5348 21788
rect 5372 21786 5428 21788
rect 5452 21786 5508 21788
rect 5532 21786 5588 21788
rect 5292 21734 5318 21786
rect 5318 21734 5348 21786
rect 5372 21734 5382 21786
rect 5382 21734 5428 21786
rect 5452 21734 5498 21786
rect 5498 21734 5508 21786
rect 5532 21734 5562 21786
rect 5562 21734 5588 21786
rect 5292 21732 5348 21734
rect 5372 21732 5428 21734
rect 5452 21732 5508 21734
rect 5532 21732 5588 21734
rect 3846 21242 3902 21244
rect 3926 21242 3982 21244
rect 4006 21242 4062 21244
rect 4086 21242 4142 21244
rect 3846 21190 3872 21242
rect 3872 21190 3902 21242
rect 3926 21190 3936 21242
rect 3936 21190 3982 21242
rect 4006 21190 4052 21242
rect 4052 21190 4062 21242
rect 4086 21190 4116 21242
rect 4116 21190 4142 21242
rect 3846 21188 3902 21190
rect 3926 21188 3982 21190
rect 4006 21188 4062 21190
rect 4086 21188 4142 21190
rect 2401 20698 2457 20700
rect 2481 20698 2537 20700
rect 2561 20698 2617 20700
rect 2641 20698 2697 20700
rect 2401 20646 2427 20698
rect 2427 20646 2457 20698
rect 2481 20646 2491 20698
rect 2491 20646 2537 20698
rect 2561 20646 2607 20698
rect 2607 20646 2617 20698
rect 2641 20646 2671 20698
rect 2671 20646 2697 20698
rect 2401 20644 2457 20646
rect 2481 20644 2537 20646
rect 2561 20644 2617 20646
rect 2641 20644 2697 20646
rect 5292 20698 5348 20700
rect 5372 20698 5428 20700
rect 5452 20698 5508 20700
rect 5532 20698 5588 20700
rect 5292 20646 5318 20698
rect 5318 20646 5348 20698
rect 5372 20646 5382 20698
rect 5382 20646 5428 20698
rect 5452 20646 5498 20698
rect 5498 20646 5508 20698
rect 5532 20646 5562 20698
rect 5562 20646 5588 20698
rect 5292 20644 5348 20646
rect 5372 20644 5428 20646
rect 5452 20644 5508 20646
rect 5532 20644 5588 20646
rect 3422 20440 3478 20496
rect 2401 19610 2457 19612
rect 2481 19610 2537 19612
rect 2561 19610 2617 19612
rect 2641 19610 2697 19612
rect 2401 19558 2427 19610
rect 2427 19558 2457 19610
rect 2481 19558 2491 19610
rect 2491 19558 2537 19610
rect 2561 19558 2607 19610
rect 2607 19558 2617 19610
rect 2641 19558 2671 19610
rect 2671 19558 2697 19610
rect 2401 19556 2457 19558
rect 2481 19556 2537 19558
rect 2561 19556 2617 19558
rect 2641 19556 2697 19558
rect 2401 18522 2457 18524
rect 2481 18522 2537 18524
rect 2561 18522 2617 18524
rect 2641 18522 2697 18524
rect 2401 18470 2427 18522
rect 2427 18470 2457 18522
rect 2481 18470 2491 18522
rect 2491 18470 2537 18522
rect 2561 18470 2607 18522
rect 2607 18470 2617 18522
rect 2641 18470 2671 18522
rect 2671 18470 2697 18522
rect 2401 18468 2457 18470
rect 2481 18468 2537 18470
rect 2561 18468 2617 18470
rect 2641 18468 2697 18470
rect 2401 17434 2457 17436
rect 2481 17434 2537 17436
rect 2561 17434 2617 17436
rect 2641 17434 2697 17436
rect 2401 17382 2427 17434
rect 2427 17382 2457 17434
rect 2481 17382 2491 17434
rect 2491 17382 2537 17434
rect 2561 17382 2607 17434
rect 2607 17382 2617 17434
rect 2641 17382 2671 17434
rect 2671 17382 2697 17434
rect 2401 17380 2457 17382
rect 2481 17380 2537 17382
rect 2561 17380 2617 17382
rect 2641 17380 2697 17382
rect 2401 16346 2457 16348
rect 2481 16346 2537 16348
rect 2561 16346 2617 16348
rect 2641 16346 2697 16348
rect 2401 16294 2427 16346
rect 2427 16294 2457 16346
rect 2481 16294 2491 16346
rect 2491 16294 2537 16346
rect 2561 16294 2607 16346
rect 2607 16294 2617 16346
rect 2641 16294 2671 16346
rect 2671 16294 2697 16346
rect 2401 16292 2457 16294
rect 2481 16292 2537 16294
rect 2561 16292 2617 16294
rect 2641 16292 2697 16294
rect 2401 15258 2457 15260
rect 2481 15258 2537 15260
rect 2561 15258 2617 15260
rect 2641 15258 2697 15260
rect 2401 15206 2427 15258
rect 2427 15206 2457 15258
rect 2481 15206 2491 15258
rect 2491 15206 2537 15258
rect 2561 15206 2607 15258
rect 2607 15206 2617 15258
rect 2641 15206 2671 15258
rect 2671 15206 2697 15258
rect 2401 15204 2457 15206
rect 2481 15204 2537 15206
rect 2561 15204 2617 15206
rect 2641 15204 2697 15206
rect 2401 14170 2457 14172
rect 2481 14170 2537 14172
rect 2561 14170 2617 14172
rect 2641 14170 2697 14172
rect 2401 14118 2427 14170
rect 2427 14118 2457 14170
rect 2481 14118 2491 14170
rect 2491 14118 2537 14170
rect 2561 14118 2607 14170
rect 2607 14118 2617 14170
rect 2641 14118 2671 14170
rect 2671 14118 2697 14170
rect 2401 14116 2457 14118
rect 2481 14116 2537 14118
rect 2561 14116 2617 14118
rect 2641 14116 2697 14118
rect 2401 13082 2457 13084
rect 2481 13082 2537 13084
rect 2561 13082 2617 13084
rect 2641 13082 2697 13084
rect 2401 13030 2427 13082
rect 2427 13030 2457 13082
rect 2481 13030 2491 13082
rect 2491 13030 2537 13082
rect 2561 13030 2607 13082
rect 2607 13030 2617 13082
rect 2641 13030 2671 13082
rect 2671 13030 2697 13082
rect 2401 13028 2457 13030
rect 2481 13028 2537 13030
rect 2561 13028 2617 13030
rect 2641 13028 2697 13030
rect 2870 12280 2926 12336
rect 2401 11994 2457 11996
rect 2481 11994 2537 11996
rect 2561 11994 2617 11996
rect 2641 11994 2697 11996
rect 2401 11942 2427 11994
rect 2427 11942 2457 11994
rect 2481 11942 2491 11994
rect 2491 11942 2537 11994
rect 2561 11942 2607 11994
rect 2607 11942 2617 11994
rect 2641 11942 2671 11994
rect 2671 11942 2697 11994
rect 2401 11940 2457 11942
rect 2481 11940 2537 11942
rect 2561 11940 2617 11942
rect 2641 11940 2697 11942
rect 2401 10906 2457 10908
rect 2481 10906 2537 10908
rect 2561 10906 2617 10908
rect 2641 10906 2697 10908
rect 2401 10854 2427 10906
rect 2427 10854 2457 10906
rect 2481 10854 2491 10906
rect 2491 10854 2537 10906
rect 2561 10854 2607 10906
rect 2607 10854 2617 10906
rect 2641 10854 2671 10906
rect 2671 10854 2697 10906
rect 2401 10852 2457 10854
rect 2481 10852 2537 10854
rect 2561 10852 2617 10854
rect 2641 10852 2697 10854
rect 2401 9818 2457 9820
rect 2481 9818 2537 9820
rect 2561 9818 2617 9820
rect 2641 9818 2697 9820
rect 2401 9766 2427 9818
rect 2427 9766 2457 9818
rect 2481 9766 2491 9818
rect 2491 9766 2537 9818
rect 2561 9766 2607 9818
rect 2607 9766 2617 9818
rect 2641 9766 2671 9818
rect 2671 9766 2697 9818
rect 2401 9764 2457 9766
rect 2481 9764 2537 9766
rect 2561 9764 2617 9766
rect 2641 9764 2697 9766
rect 2401 8730 2457 8732
rect 2481 8730 2537 8732
rect 2561 8730 2617 8732
rect 2641 8730 2697 8732
rect 2401 8678 2427 8730
rect 2427 8678 2457 8730
rect 2481 8678 2491 8730
rect 2491 8678 2537 8730
rect 2561 8678 2607 8730
rect 2607 8678 2617 8730
rect 2641 8678 2671 8730
rect 2671 8678 2697 8730
rect 2401 8676 2457 8678
rect 2481 8676 2537 8678
rect 2561 8676 2617 8678
rect 2641 8676 2697 8678
rect 2401 7642 2457 7644
rect 2481 7642 2537 7644
rect 2561 7642 2617 7644
rect 2641 7642 2697 7644
rect 2401 7590 2427 7642
rect 2427 7590 2457 7642
rect 2481 7590 2491 7642
rect 2491 7590 2537 7642
rect 2561 7590 2607 7642
rect 2607 7590 2617 7642
rect 2641 7590 2671 7642
rect 2671 7590 2697 7642
rect 2401 7588 2457 7590
rect 2481 7588 2537 7590
rect 2561 7588 2617 7590
rect 2641 7588 2697 7590
rect 2401 6554 2457 6556
rect 2481 6554 2537 6556
rect 2561 6554 2617 6556
rect 2641 6554 2697 6556
rect 2401 6502 2427 6554
rect 2427 6502 2457 6554
rect 2481 6502 2491 6554
rect 2491 6502 2537 6554
rect 2561 6502 2607 6554
rect 2607 6502 2617 6554
rect 2641 6502 2671 6554
rect 2671 6502 2697 6554
rect 2401 6500 2457 6502
rect 2481 6500 2537 6502
rect 2561 6500 2617 6502
rect 2641 6500 2697 6502
rect 2401 5466 2457 5468
rect 2481 5466 2537 5468
rect 2561 5466 2617 5468
rect 2641 5466 2697 5468
rect 2401 5414 2427 5466
rect 2427 5414 2457 5466
rect 2481 5414 2491 5466
rect 2491 5414 2537 5466
rect 2561 5414 2607 5466
rect 2607 5414 2617 5466
rect 2641 5414 2671 5466
rect 2671 5414 2697 5466
rect 2401 5412 2457 5414
rect 2481 5412 2537 5414
rect 2561 5412 2617 5414
rect 2641 5412 2697 5414
rect 2401 4378 2457 4380
rect 2481 4378 2537 4380
rect 2561 4378 2617 4380
rect 2641 4378 2697 4380
rect 2401 4326 2427 4378
rect 2427 4326 2457 4378
rect 2481 4326 2491 4378
rect 2491 4326 2537 4378
rect 2561 4326 2607 4378
rect 2607 4326 2617 4378
rect 2641 4326 2671 4378
rect 2671 4326 2697 4378
rect 2401 4324 2457 4326
rect 2481 4324 2537 4326
rect 2561 4324 2617 4326
rect 2641 4324 2697 4326
rect 3846 20154 3902 20156
rect 3926 20154 3982 20156
rect 4006 20154 4062 20156
rect 4086 20154 4142 20156
rect 3846 20102 3872 20154
rect 3872 20102 3902 20154
rect 3926 20102 3936 20154
rect 3936 20102 3982 20154
rect 4006 20102 4052 20154
rect 4052 20102 4062 20154
rect 4086 20102 4116 20154
rect 4116 20102 4142 20154
rect 3846 20100 3902 20102
rect 3926 20100 3982 20102
rect 4006 20100 4062 20102
rect 4086 20100 4142 20102
rect 3846 19066 3902 19068
rect 3926 19066 3982 19068
rect 4006 19066 4062 19068
rect 4086 19066 4142 19068
rect 3846 19014 3872 19066
rect 3872 19014 3902 19066
rect 3926 19014 3936 19066
rect 3936 19014 3982 19066
rect 4006 19014 4052 19066
rect 4052 19014 4062 19066
rect 4086 19014 4116 19066
rect 4116 19014 4142 19066
rect 3846 19012 3902 19014
rect 3926 19012 3982 19014
rect 4006 19012 4062 19014
rect 4086 19012 4142 19014
rect 3846 17978 3902 17980
rect 3926 17978 3982 17980
rect 4006 17978 4062 17980
rect 4086 17978 4142 17980
rect 3846 17926 3872 17978
rect 3872 17926 3902 17978
rect 3926 17926 3936 17978
rect 3936 17926 3982 17978
rect 4006 17926 4052 17978
rect 4052 17926 4062 17978
rect 4086 17926 4116 17978
rect 4116 17926 4142 17978
rect 3846 17924 3902 17926
rect 3926 17924 3982 17926
rect 4006 17924 4062 17926
rect 4086 17924 4142 17926
rect 3846 16890 3902 16892
rect 3926 16890 3982 16892
rect 4006 16890 4062 16892
rect 4086 16890 4142 16892
rect 3846 16838 3872 16890
rect 3872 16838 3902 16890
rect 3926 16838 3936 16890
rect 3936 16838 3982 16890
rect 4006 16838 4052 16890
rect 4052 16838 4062 16890
rect 4086 16838 4116 16890
rect 4116 16838 4142 16890
rect 3846 16836 3902 16838
rect 3926 16836 3982 16838
rect 4006 16836 4062 16838
rect 4086 16836 4142 16838
rect 3846 15802 3902 15804
rect 3926 15802 3982 15804
rect 4006 15802 4062 15804
rect 4086 15802 4142 15804
rect 3846 15750 3872 15802
rect 3872 15750 3902 15802
rect 3926 15750 3936 15802
rect 3936 15750 3982 15802
rect 4006 15750 4052 15802
rect 4052 15750 4062 15802
rect 4086 15750 4116 15802
rect 4116 15750 4142 15802
rect 3846 15748 3902 15750
rect 3926 15748 3982 15750
rect 4006 15748 4062 15750
rect 4086 15748 4142 15750
rect 3846 14714 3902 14716
rect 3926 14714 3982 14716
rect 4006 14714 4062 14716
rect 4086 14714 4142 14716
rect 3846 14662 3872 14714
rect 3872 14662 3902 14714
rect 3926 14662 3936 14714
rect 3936 14662 3982 14714
rect 4006 14662 4052 14714
rect 4052 14662 4062 14714
rect 4086 14662 4116 14714
rect 4116 14662 4142 14714
rect 3846 14660 3902 14662
rect 3926 14660 3982 14662
rect 4006 14660 4062 14662
rect 4086 14660 4142 14662
rect 3846 13626 3902 13628
rect 3926 13626 3982 13628
rect 4006 13626 4062 13628
rect 4086 13626 4142 13628
rect 3846 13574 3872 13626
rect 3872 13574 3902 13626
rect 3926 13574 3936 13626
rect 3936 13574 3982 13626
rect 4006 13574 4052 13626
rect 4052 13574 4062 13626
rect 4086 13574 4116 13626
rect 4116 13574 4142 13626
rect 3846 13572 3902 13574
rect 3926 13572 3982 13574
rect 4006 13572 4062 13574
rect 4086 13572 4142 13574
rect 3846 12538 3902 12540
rect 3926 12538 3982 12540
rect 4006 12538 4062 12540
rect 4086 12538 4142 12540
rect 3846 12486 3872 12538
rect 3872 12486 3902 12538
rect 3926 12486 3936 12538
rect 3936 12486 3982 12538
rect 4006 12486 4052 12538
rect 4052 12486 4062 12538
rect 4086 12486 4116 12538
rect 4116 12486 4142 12538
rect 3846 12484 3902 12486
rect 3926 12484 3982 12486
rect 4006 12484 4062 12486
rect 4086 12484 4142 12486
rect 3846 11450 3902 11452
rect 3926 11450 3982 11452
rect 4006 11450 4062 11452
rect 4086 11450 4142 11452
rect 3846 11398 3872 11450
rect 3872 11398 3902 11450
rect 3926 11398 3936 11450
rect 3936 11398 3982 11450
rect 4006 11398 4052 11450
rect 4052 11398 4062 11450
rect 4086 11398 4116 11450
rect 4116 11398 4142 11450
rect 3846 11396 3902 11398
rect 3926 11396 3982 11398
rect 4006 11396 4062 11398
rect 4086 11396 4142 11398
rect 3846 10362 3902 10364
rect 3926 10362 3982 10364
rect 4006 10362 4062 10364
rect 4086 10362 4142 10364
rect 3846 10310 3872 10362
rect 3872 10310 3902 10362
rect 3926 10310 3936 10362
rect 3936 10310 3982 10362
rect 4006 10310 4052 10362
rect 4052 10310 4062 10362
rect 4086 10310 4116 10362
rect 4116 10310 4142 10362
rect 3846 10308 3902 10310
rect 3926 10308 3982 10310
rect 4006 10308 4062 10310
rect 4086 10308 4142 10310
rect 3846 9274 3902 9276
rect 3926 9274 3982 9276
rect 4006 9274 4062 9276
rect 4086 9274 4142 9276
rect 3846 9222 3872 9274
rect 3872 9222 3902 9274
rect 3926 9222 3936 9274
rect 3936 9222 3982 9274
rect 4006 9222 4052 9274
rect 4052 9222 4062 9274
rect 4086 9222 4116 9274
rect 4116 9222 4142 9274
rect 3846 9220 3902 9222
rect 3926 9220 3982 9222
rect 4006 9220 4062 9222
rect 4086 9220 4142 9222
rect 3846 8186 3902 8188
rect 3926 8186 3982 8188
rect 4006 8186 4062 8188
rect 4086 8186 4142 8188
rect 3846 8134 3872 8186
rect 3872 8134 3902 8186
rect 3926 8134 3936 8186
rect 3936 8134 3982 8186
rect 4006 8134 4052 8186
rect 4052 8134 4062 8186
rect 4086 8134 4116 8186
rect 4116 8134 4142 8186
rect 3846 8132 3902 8134
rect 3926 8132 3982 8134
rect 4006 8132 4062 8134
rect 4086 8132 4142 8134
rect 3846 7098 3902 7100
rect 3926 7098 3982 7100
rect 4006 7098 4062 7100
rect 4086 7098 4142 7100
rect 3846 7046 3872 7098
rect 3872 7046 3902 7098
rect 3926 7046 3936 7098
rect 3936 7046 3982 7098
rect 4006 7046 4052 7098
rect 4052 7046 4062 7098
rect 4086 7046 4116 7098
rect 4116 7046 4142 7098
rect 3846 7044 3902 7046
rect 3926 7044 3982 7046
rect 4006 7044 4062 7046
rect 4086 7044 4142 7046
rect 3846 6010 3902 6012
rect 3926 6010 3982 6012
rect 4006 6010 4062 6012
rect 4086 6010 4142 6012
rect 3846 5958 3872 6010
rect 3872 5958 3902 6010
rect 3926 5958 3936 6010
rect 3936 5958 3982 6010
rect 4006 5958 4052 6010
rect 4052 5958 4062 6010
rect 4086 5958 4116 6010
rect 4116 5958 4142 6010
rect 3846 5956 3902 5958
rect 3926 5956 3982 5958
rect 4006 5956 4062 5958
rect 4086 5956 4142 5958
rect 3846 4922 3902 4924
rect 3926 4922 3982 4924
rect 4006 4922 4062 4924
rect 4086 4922 4142 4924
rect 3846 4870 3872 4922
rect 3872 4870 3902 4922
rect 3926 4870 3936 4922
rect 3936 4870 3982 4922
rect 4006 4870 4052 4922
rect 4052 4870 4062 4922
rect 4086 4870 4116 4922
rect 4116 4870 4142 4922
rect 3846 4868 3902 4870
rect 3926 4868 3982 4870
rect 4006 4868 4062 4870
rect 4086 4868 4142 4870
rect 3330 4120 3386 4176
rect 3846 3834 3902 3836
rect 3926 3834 3982 3836
rect 4006 3834 4062 3836
rect 4086 3834 4142 3836
rect 3846 3782 3872 3834
rect 3872 3782 3902 3834
rect 3926 3782 3936 3834
rect 3936 3782 3982 3834
rect 4006 3782 4052 3834
rect 4052 3782 4062 3834
rect 4086 3782 4116 3834
rect 4116 3782 4142 3834
rect 3846 3780 3902 3782
rect 3926 3780 3982 3782
rect 4006 3780 4062 3782
rect 4086 3780 4142 3782
rect 2401 3290 2457 3292
rect 2481 3290 2537 3292
rect 2561 3290 2617 3292
rect 2641 3290 2697 3292
rect 2401 3238 2427 3290
rect 2427 3238 2457 3290
rect 2481 3238 2491 3290
rect 2491 3238 2537 3290
rect 2561 3238 2607 3290
rect 2607 3238 2617 3290
rect 2641 3238 2671 3290
rect 2671 3238 2697 3290
rect 2401 3236 2457 3238
rect 2481 3236 2537 3238
rect 2561 3236 2617 3238
rect 2641 3236 2697 3238
rect 3846 2746 3902 2748
rect 3926 2746 3982 2748
rect 4006 2746 4062 2748
rect 4086 2746 4142 2748
rect 3846 2694 3872 2746
rect 3872 2694 3902 2746
rect 3926 2694 3936 2746
rect 3936 2694 3982 2746
rect 4006 2694 4052 2746
rect 4052 2694 4062 2746
rect 4086 2694 4116 2746
rect 4116 2694 4142 2746
rect 3846 2692 3902 2694
rect 3926 2692 3982 2694
rect 4006 2692 4062 2694
rect 4086 2692 4142 2694
rect 2401 2202 2457 2204
rect 2481 2202 2537 2204
rect 2561 2202 2617 2204
rect 2641 2202 2697 2204
rect 2401 2150 2427 2202
rect 2427 2150 2457 2202
rect 2481 2150 2491 2202
rect 2491 2150 2537 2202
rect 2561 2150 2607 2202
rect 2607 2150 2617 2202
rect 2641 2150 2671 2202
rect 2671 2150 2697 2202
rect 2401 2148 2457 2150
rect 2481 2148 2537 2150
rect 2561 2148 2617 2150
rect 2641 2148 2697 2150
rect 5630 19760 5686 19816
rect 5292 19610 5348 19612
rect 5372 19610 5428 19612
rect 5452 19610 5508 19612
rect 5532 19610 5588 19612
rect 5292 19558 5318 19610
rect 5318 19558 5348 19610
rect 5372 19558 5382 19610
rect 5382 19558 5428 19610
rect 5452 19558 5498 19610
rect 5498 19558 5508 19610
rect 5532 19558 5562 19610
rect 5562 19558 5588 19610
rect 5292 19556 5348 19558
rect 5372 19556 5428 19558
rect 5452 19556 5508 19558
rect 5532 19556 5588 19558
rect 5292 18522 5348 18524
rect 5372 18522 5428 18524
rect 5452 18522 5508 18524
rect 5532 18522 5588 18524
rect 5292 18470 5318 18522
rect 5318 18470 5348 18522
rect 5372 18470 5382 18522
rect 5382 18470 5428 18522
rect 5452 18470 5498 18522
rect 5498 18470 5508 18522
rect 5532 18470 5562 18522
rect 5562 18470 5588 18522
rect 5292 18468 5348 18470
rect 5372 18468 5428 18470
rect 5452 18468 5508 18470
rect 5532 18468 5588 18470
rect 5292 17434 5348 17436
rect 5372 17434 5428 17436
rect 5452 17434 5508 17436
rect 5532 17434 5588 17436
rect 5292 17382 5318 17434
rect 5318 17382 5348 17434
rect 5372 17382 5382 17434
rect 5382 17382 5428 17434
rect 5452 17382 5498 17434
rect 5498 17382 5508 17434
rect 5532 17382 5562 17434
rect 5562 17382 5588 17434
rect 5292 17380 5348 17382
rect 5372 17380 5428 17382
rect 5452 17380 5508 17382
rect 5532 17380 5588 17382
rect 5292 16346 5348 16348
rect 5372 16346 5428 16348
rect 5452 16346 5508 16348
rect 5532 16346 5588 16348
rect 5292 16294 5318 16346
rect 5318 16294 5348 16346
rect 5372 16294 5382 16346
rect 5382 16294 5428 16346
rect 5452 16294 5498 16346
rect 5498 16294 5508 16346
rect 5532 16294 5562 16346
rect 5562 16294 5588 16346
rect 5292 16292 5348 16294
rect 5372 16292 5428 16294
rect 5452 16292 5508 16294
rect 5532 16292 5588 16294
rect 5292 15258 5348 15260
rect 5372 15258 5428 15260
rect 5452 15258 5508 15260
rect 5532 15258 5588 15260
rect 5292 15206 5318 15258
rect 5318 15206 5348 15258
rect 5372 15206 5382 15258
rect 5382 15206 5428 15258
rect 5452 15206 5498 15258
rect 5498 15206 5508 15258
rect 5532 15206 5562 15258
rect 5562 15206 5588 15258
rect 5292 15204 5348 15206
rect 5372 15204 5428 15206
rect 5452 15204 5508 15206
rect 5532 15204 5588 15206
rect 5292 14170 5348 14172
rect 5372 14170 5428 14172
rect 5452 14170 5508 14172
rect 5532 14170 5588 14172
rect 5292 14118 5318 14170
rect 5318 14118 5348 14170
rect 5372 14118 5382 14170
rect 5382 14118 5428 14170
rect 5452 14118 5498 14170
rect 5498 14118 5508 14170
rect 5532 14118 5562 14170
rect 5562 14118 5588 14170
rect 5292 14116 5348 14118
rect 5372 14116 5428 14118
rect 5452 14116 5508 14118
rect 5532 14116 5588 14118
rect 5630 13912 5686 13968
rect 5292 13082 5348 13084
rect 5372 13082 5428 13084
rect 5452 13082 5508 13084
rect 5532 13082 5588 13084
rect 5292 13030 5318 13082
rect 5318 13030 5348 13082
rect 5372 13030 5382 13082
rect 5382 13030 5428 13082
rect 5452 13030 5498 13082
rect 5498 13030 5508 13082
rect 5532 13030 5562 13082
rect 5562 13030 5588 13082
rect 5292 13028 5348 13030
rect 5372 13028 5428 13030
rect 5452 13028 5508 13030
rect 5532 13028 5588 13030
rect 5630 12144 5686 12200
rect 5292 11994 5348 11996
rect 5372 11994 5428 11996
rect 5452 11994 5508 11996
rect 5532 11994 5588 11996
rect 5292 11942 5318 11994
rect 5318 11942 5348 11994
rect 5372 11942 5382 11994
rect 5382 11942 5428 11994
rect 5452 11942 5498 11994
rect 5498 11942 5508 11994
rect 5532 11942 5562 11994
rect 5562 11942 5588 11994
rect 5292 11940 5348 11942
rect 5372 11940 5428 11942
rect 5452 11940 5508 11942
rect 5532 11940 5588 11942
rect 5292 10906 5348 10908
rect 5372 10906 5428 10908
rect 5452 10906 5508 10908
rect 5532 10906 5588 10908
rect 5292 10854 5318 10906
rect 5318 10854 5348 10906
rect 5372 10854 5382 10906
rect 5382 10854 5428 10906
rect 5452 10854 5498 10906
rect 5498 10854 5508 10906
rect 5532 10854 5562 10906
rect 5562 10854 5588 10906
rect 5292 10852 5348 10854
rect 5372 10852 5428 10854
rect 5452 10852 5508 10854
rect 5532 10852 5588 10854
rect 5292 9818 5348 9820
rect 5372 9818 5428 9820
rect 5452 9818 5508 9820
rect 5532 9818 5588 9820
rect 5292 9766 5318 9818
rect 5318 9766 5348 9818
rect 5372 9766 5382 9818
rect 5382 9766 5428 9818
rect 5452 9766 5498 9818
rect 5498 9766 5508 9818
rect 5532 9766 5562 9818
rect 5562 9766 5588 9818
rect 5292 9764 5348 9766
rect 5372 9764 5428 9766
rect 5452 9764 5508 9766
rect 5532 9764 5588 9766
rect 5292 8730 5348 8732
rect 5372 8730 5428 8732
rect 5452 8730 5508 8732
rect 5532 8730 5588 8732
rect 5292 8678 5318 8730
rect 5318 8678 5348 8730
rect 5372 8678 5382 8730
rect 5382 8678 5428 8730
rect 5452 8678 5498 8730
rect 5498 8678 5508 8730
rect 5532 8678 5562 8730
rect 5562 8678 5588 8730
rect 5292 8676 5348 8678
rect 5372 8676 5428 8678
rect 5452 8676 5508 8678
rect 5532 8676 5588 8678
rect 5292 7642 5348 7644
rect 5372 7642 5428 7644
rect 5452 7642 5508 7644
rect 5532 7642 5588 7644
rect 5292 7590 5318 7642
rect 5318 7590 5348 7642
rect 5372 7590 5382 7642
rect 5382 7590 5428 7642
rect 5452 7590 5498 7642
rect 5498 7590 5508 7642
rect 5532 7590 5562 7642
rect 5562 7590 5588 7642
rect 5292 7588 5348 7590
rect 5372 7588 5428 7590
rect 5452 7588 5508 7590
rect 5532 7588 5588 7590
rect 5292 6554 5348 6556
rect 5372 6554 5428 6556
rect 5452 6554 5508 6556
rect 5532 6554 5588 6556
rect 5292 6502 5318 6554
rect 5318 6502 5348 6554
rect 5372 6502 5382 6554
rect 5382 6502 5428 6554
rect 5452 6502 5498 6554
rect 5498 6502 5508 6554
rect 5532 6502 5562 6554
rect 5562 6502 5588 6554
rect 5292 6500 5348 6502
rect 5372 6500 5428 6502
rect 5452 6500 5508 6502
rect 5532 6500 5588 6502
rect 5292 5466 5348 5468
rect 5372 5466 5428 5468
rect 5452 5466 5508 5468
rect 5532 5466 5588 5468
rect 5292 5414 5318 5466
rect 5318 5414 5348 5466
rect 5372 5414 5382 5466
rect 5382 5414 5428 5466
rect 5452 5414 5498 5466
rect 5498 5414 5508 5466
rect 5532 5414 5562 5466
rect 5562 5414 5588 5466
rect 5292 5412 5348 5414
rect 5372 5412 5428 5414
rect 5452 5412 5508 5414
rect 5532 5412 5588 5414
rect 5630 4528 5686 4584
rect 5292 4378 5348 4380
rect 5372 4378 5428 4380
rect 5452 4378 5508 4380
rect 5532 4378 5588 4380
rect 5292 4326 5318 4378
rect 5318 4326 5348 4378
rect 5372 4326 5382 4378
rect 5382 4326 5428 4378
rect 5452 4326 5498 4378
rect 5498 4326 5508 4378
rect 5532 4326 5562 4378
rect 5562 4326 5588 4378
rect 5292 4324 5348 4326
rect 5372 4324 5428 4326
rect 5452 4324 5508 4326
rect 5532 4324 5588 4326
rect 5292 3290 5348 3292
rect 5372 3290 5428 3292
rect 5452 3290 5508 3292
rect 5532 3290 5588 3292
rect 5292 3238 5318 3290
rect 5318 3238 5348 3290
rect 5372 3238 5382 3290
rect 5382 3238 5428 3290
rect 5452 3238 5498 3290
rect 5498 3238 5508 3290
rect 5532 3238 5562 3290
rect 5562 3238 5588 3290
rect 5292 3236 5348 3238
rect 5372 3236 5428 3238
rect 5452 3236 5508 3238
rect 5532 3236 5588 3238
rect 6458 15544 6514 15600
rect 6182 6704 6238 6760
rect 6737 22330 6793 22332
rect 6817 22330 6873 22332
rect 6897 22330 6953 22332
rect 6977 22330 7033 22332
rect 6737 22278 6763 22330
rect 6763 22278 6793 22330
rect 6817 22278 6827 22330
rect 6827 22278 6873 22330
rect 6897 22278 6943 22330
rect 6943 22278 6953 22330
rect 6977 22278 7007 22330
rect 7007 22278 7033 22330
rect 6737 22276 6793 22278
rect 6817 22276 6873 22278
rect 6897 22276 6953 22278
rect 6977 22276 7033 22278
rect 7102 21528 7158 21584
rect 6737 21242 6793 21244
rect 6817 21242 6873 21244
rect 6897 21242 6953 21244
rect 6977 21242 7033 21244
rect 6737 21190 6763 21242
rect 6763 21190 6793 21242
rect 6817 21190 6827 21242
rect 6827 21190 6873 21242
rect 6897 21190 6943 21242
rect 6943 21190 6953 21242
rect 6977 21190 7007 21242
rect 7007 21190 7033 21242
rect 6737 21188 6793 21190
rect 6817 21188 6873 21190
rect 6897 21188 6953 21190
rect 6977 21188 7033 21190
rect 6737 20154 6793 20156
rect 6817 20154 6873 20156
rect 6897 20154 6953 20156
rect 6977 20154 7033 20156
rect 6737 20102 6763 20154
rect 6763 20102 6793 20154
rect 6817 20102 6827 20154
rect 6827 20102 6873 20154
rect 6897 20102 6943 20154
rect 6943 20102 6953 20154
rect 6977 20102 7007 20154
rect 7007 20102 7033 20154
rect 6737 20100 6793 20102
rect 6817 20100 6873 20102
rect 6897 20100 6953 20102
rect 6977 20100 7033 20102
rect 6737 19066 6793 19068
rect 6817 19066 6873 19068
rect 6897 19066 6953 19068
rect 6977 19066 7033 19068
rect 6737 19014 6763 19066
rect 6763 19014 6793 19066
rect 6817 19014 6827 19066
rect 6827 19014 6873 19066
rect 6897 19014 6943 19066
rect 6943 19014 6953 19066
rect 6977 19014 7007 19066
rect 7007 19014 7033 19066
rect 6737 19012 6793 19014
rect 6817 19012 6873 19014
rect 6897 19012 6953 19014
rect 6977 19012 7033 19014
rect 6737 17978 6793 17980
rect 6817 17978 6873 17980
rect 6897 17978 6953 17980
rect 6977 17978 7033 17980
rect 6737 17926 6763 17978
rect 6763 17926 6793 17978
rect 6817 17926 6827 17978
rect 6827 17926 6873 17978
rect 6897 17926 6943 17978
rect 6943 17926 6953 17978
rect 6977 17926 7007 17978
rect 7007 17926 7033 17978
rect 6737 17924 6793 17926
rect 6817 17924 6873 17926
rect 6897 17924 6953 17926
rect 6977 17924 7033 17926
rect 6737 16890 6793 16892
rect 6817 16890 6873 16892
rect 6897 16890 6953 16892
rect 6977 16890 7033 16892
rect 6737 16838 6763 16890
rect 6763 16838 6793 16890
rect 6817 16838 6827 16890
rect 6827 16838 6873 16890
rect 6897 16838 6943 16890
rect 6943 16838 6953 16890
rect 6977 16838 7007 16890
rect 7007 16838 7033 16890
rect 6737 16836 6793 16838
rect 6817 16836 6873 16838
rect 6897 16836 6953 16838
rect 6977 16836 7033 16838
rect 6737 15802 6793 15804
rect 6817 15802 6873 15804
rect 6897 15802 6953 15804
rect 6977 15802 7033 15804
rect 6737 15750 6763 15802
rect 6763 15750 6793 15802
rect 6817 15750 6827 15802
rect 6827 15750 6873 15802
rect 6897 15750 6943 15802
rect 6943 15750 6953 15802
rect 6977 15750 7007 15802
rect 7007 15750 7033 15802
rect 6737 15748 6793 15750
rect 6817 15748 6873 15750
rect 6897 15748 6953 15750
rect 6977 15748 7033 15750
rect 6737 14714 6793 14716
rect 6817 14714 6873 14716
rect 6897 14714 6953 14716
rect 6977 14714 7033 14716
rect 6737 14662 6763 14714
rect 6763 14662 6793 14714
rect 6817 14662 6827 14714
rect 6827 14662 6873 14714
rect 6897 14662 6943 14714
rect 6943 14662 6953 14714
rect 6977 14662 7007 14714
rect 7007 14662 7033 14714
rect 6737 14660 6793 14662
rect 6817 14660 6873 14662
rect 6897 14660 6953 14662
rect 6977 14660 7033 14662
rect 6737 13626 6793 13628
rect 6817 13626 6873 13628
rect 6897 13626 6953 13628
rect 6977 13626 7033 13628
rect 6737 13574 6763 13626
rect 6763 13574 6793 13626
rect 6817 13574 6827 13626
rect 6827 13574 6873 13626
rect 6897 13574 6943 13626
rect 6943 13574 6953 13626
rect 6977 13574 7007 13626
rect 7007 13574 7033 13626
rect 6737 13572 6793 13574
rect 6817 13572 6873 13574
rect 6897 13572 6953 13574
rect 6977 13572 7033 13574
rect 6737 12538 6793 12540
rect 6817 12538 6873 12540
rect 6897 12538 6953 12540
rect 6977 12538 7033 12540
rect 6737 12486 6763 12538
rect 6763 12486 6793 12538
rect 6817 12486 6827 12538
rect 6827 12486 6873 12538
rect 6897 12486 6943 12538
rect 6943 12486 6953 12538
rect 6977 12486 7007 12538
rect 7007 12486 7033 12538
rect 6737 12484 6793 12486
rect 6817 12484 6873 12486
rect 6897 12484 6953 12486
rect 6977 12484 7033 12486
rect 6737 11450 6793 11452
rect 6817 11450 6873 11452
rect 6897 11450 6953 11452
rect 6977 11450 7033 11452
rect 6737 11398 6763 11450
rect 6763 11398 6793 11450
rect 6817 11398 6827 11450
rect 6827 11398 6873 11450
rect 6897 11398 6943 11450
rect 6943 11398 6953 11450
rect 6977 11398 7007 11450
rect 7007 11398 7033 11450
rect 6737 11396 6793 11398
rect 6817 11396 6873 11398
rect 6897 11396 6953 11398
rect 6977 11396 7033 11398
rect 6550 10512 6606 10568
rect 6737 10362 6793 10364
rect 6817 10362 6873 10364
rect 6897 10362 6953 10364
rect 6977 10362 7033 10364
rect 6737 10310 6763 10362
rect 6763 10310 6793 10362
rect 6817 10310 6827 10362
rect 6827 10310 6873 10362
rect 6897 10310 6943 10362
rect 6943 10310 6953 10362
rect 6977 10310 7007 10362
rect 7007 10310 7033 10362
rect 6737 10308 6793 10310
rect 6817 10308 6873 10310
rect 6897 10308 6953 10310
rect 6977 10308 7033 10310
rect 6737 9274 6793 9276
rect 6817 9274 6873 9276
rect 6897 9274 6953 9276
rect 6977 9274 7033 9276
rect 6737 9222 6763 9274
rect 6763 9222 6793 9274
rect 6817 9222 6827 9274
rect 6827 9222 6873 9274
rect 6897 9222 6943 9274
rect 6943 9222 6953 9274
rect 6977 9222 7007 9274
rect 7007 9222 7033 9274
rect 6737 9220 6793 9222
rect 6817 9220 6873 9222
rect 6897 9220 6953 9222
rect 6977 9220 7033 9222
rect 6642 8336 6698 8392
rect 6737 8186 6793 8188
rect 6817 8186 6873 8188
rect 6897 8186 6953 8188
rect 6977 8186 7033 8188
rect 6737 8134 6763 8186
rect 6763 8134 6793 8186
rect 6817 8134 6827 8186
rect 6827 8134 6873 8186
rect 6897 8134 6943 8186
rect 6943 8134 6953 8186
rect 6977 8134 7007 8186
rect 7007 8134 7033 8186
rect 6737 8132 6793 8134
rect 6817 8132 6873 8134
rect 6897 8132 6953 8134
rect 6977 8132 7033 8134
rect 6737 7098 6793 7100
rect 6817 7098 6873 7100
rect 6897 7098 6953 7100
rect 6977 7098 7033 7100
rect 6737 7046 6763 7098
rect 6763 7046 6793 7098
rect 6817 7046 6827 7098
rect 6827 7046 6873 7098
rect 6897 7046 6943 7098
rect 6943 7046 6953 7098
rect 6977 7046 7007 7098
rect 7007 7046 7033 7098
rect 6737 7044 6793 7046
rect 6817 7044 6873 7046
rect 6897 7044 6953 7046
rect 6977 7044 7033 7046
rect 6737 6010 6793 6012
rect 6817 6010 6873 6012
rect 6897 6010 6953 6012
rect 6977 6010 7033 6012
rect 6737 5958 6763 6010
rect 6763 5958 6793 6010
rect 6817 5958 6827 6010
rect 6827 5958 6873 6010
rect 6897 5958 6943 6010
rect 6943 5958 6953 6010
rect 6977 5958 7007 6010
rect 7007 5958 7033 6010
rect 6737 5956 6793 5958
rect 6817 5956 6873 5958
rect 6897 5956 6953 5958
rect 6977 5956 7033 5958
rect 6737 4922 6793 4924
rect 6817 4922 6873 4924
rect 6897 4922 6953 4924
rect 6977 4922 7033 4924
rect 6737 4870 6763 4922
rect 6763 4870 6793 4922
rect 6817 4870 6827 4922
rect 6827 4870 6873 4922
rect 6897 4870 6943 4922
rect 6943 4870 6953 4922
rect 6977 4870 7007 4922
rect 7007 4870 7033 4922
rect 6737 4868 6793 4870
rect 6817 4868 6873 4870
rect 6897 4868 6953 4870
rect 6977 4868 7033 4870
rect 8182 21786 8238 21788
rect 8262 21786 8318 21788
rect 8342 21786 8398 21788
rect 8422 21786 8478 21788
rect 8182 21734 8208 21786
rect 8208 21734 8238 21786
rect 8262 21734 8272 21786
rect 8272 21734 8318 21786
rect 8342 21734 8388 21786
rect 8388 21734 8398 21786
rect 8422 21734 8452 21786
rect 8452 21734 8478 21786
rect 8182 21732 8238 21734
rect 8262 21732 8318 21734
rect 8342 21732 8398 21734
rect 8422 21732 8478 21734
rect 8182 20698 8238 20700
rect 8262 20698 8318 20700
rect 8342 20698 8398 20700
rect 8422 20698 8478 20700
rect 8182 20646 8208 20698
rect 8208 20646 8238 20698
rect 8262 20646 8272 20698
rect 8272 20646 8318 20698
rect 8342 20646 8388 20698
rect 8388 20646 8398 20698
rect 8422 20646 8452 20698
rect 8452 20646 8478 20698
rect 8182 20644 8238 20646
rect 8262 20644 8318 20646
rect 8342 20644 8398 20646
rect 8422 20644 8478 20646
rect 8182 19610 8238 19612
rect 8262 19610 8318 19612
rect 8342 19610 8398 19612
rect 8422 19610 8478 19612
rect 8182 19558 8208 19610
rect 8208 19558 8238 19610
rect 8262 19558 8272 19610
rect 8272 19558 8318 19610
rect 8342 19558 8388 19610
rect 8388 19558 8398 19610
rect 8422 19558 8452 19610
rect 8452 19558 8478 19610
rect 8182 19556 8238 19558
rect 8262 19556 8318 19558
rect 8342 19556 8398 19558
rect 8422 19556 8478 19558
rect 8182 18522 8238 18524
rect 8262 18522 8318 18524
rect 8342 18522 8398 18524
rect 8422 18522 8478 18524
rect 8182 18470 8208 18522
rect 8208 18470 8238 18522
rect 8262 18470 8272 18522
rect 8272 18470 8318 18522
rect 8342 18470 8388 18522
rect 8388 18470 8398 18522
rect 8422 18470 8452 18522
rect 8452 18470 8478 18522
rect 8182 18468 8238 18470
rect 8262 18468 8318 18470
rect 8342 18468 8398 18470
rect 8422 18468 8478 18470
rect 8206 17720 8262 17776
rect 8182 17434 8238 17436
rect 8262 17434 8318 17436
rect 8342 17434 8398 17436
rect 8422 17434 8478 17436
rect 8182 17382 8208 17434
rect 8208 17382 8238 17434
rect 8262 17382 8272 17434
rect 8272 17382 8318 17434
rect 8342 17382 8388 17434
rect 8388 17382 8398 17434
rect 8422 17382 8452 17434
rect 8452 17382 8478 17434
rect 8182 17380 8238 17382
rect 8262 17380 8318 17382
rect 8342 17380 8398 17382
rect 8422 17380 8478 17382
rect 8182 16346 8238 16348
rect 8262 16346 8318 16348
rect 8342 16346 8398 16348
rect 8422 16346 8478 16348
rect 8182 16294 8208 16346
rect 8208 16294 8238 16346
rect 8262 16294 8272 16346
rect 8272 16294 8318 16346
rect 8342 16294 8388 16346
rect 8388 16294 8398 16346
rect 8422 16294 8452 16346
rect 8452 16294 8478 16346
rect 8182 16292 8238 16294
rect 8262 16292 8318 16294
rect 8342 16292 8398 16294
rect 8422 16292 8478 16294
rect 8182 15258 8238 15260
rect 8262 15258 8318 15260
rect 8342 15258 8398 15260
rect 8422 15258 8478 15260
rect 8182 15206 8208 15258
rect 8208 15206 8238 15258
rect 8262 15206 8272 15258
rect 8272 15206 8318 15258
rect 8342 15206 8388 15258
rect 8388 15206 8398 15258
rect 8422 15206 8452 15258
rect 8452 15206 8478 15258
rect 8182 15204 8238 15206
rect 8262 15204 8318 15206
rect 8342 15204 8398 15206
rect 8422 15204 8478 15206
rect 8182 14170 8238 14172
rect 8262 14170 8318 14172
rect 8342 14170 8398 14172
rect 8422 14170 8478 14172
rect 8182 14118 8208 14170
rect 8208 14118 8238 14170
rect 8262 14118 8272 14170
rect 8272 14118 8318 14170
rect 8342 14118 8388 14170
rect 8388 14118 8398 14170
rect 8422 14118 8452 14170
rect 8452 14118 8478 14170
rect 8182 14116 8238 14118
rect 8262 14116 8318 14118
rect 8342 14116 8398 14118
rect 8422 14116 8478 14118
rect 8182 13082 8238 13084
rect 8262 13082 8318 13084
rect 8342 13082 8398 13084
rect 8422 13082 8478 13084
rect 8182 13030 8208 13082
rect 8208 13030 8238 13082
rect 8262 13030 8272 13082
rect 8272 13030 8318 13082
rect 8342 13030 8388 13082
rect 8388 13030 8398 13082
rect 8422 13030 8452 13082
rect 8452 13030 8478 13082
rect 8182 13028 8238 13030
rect 8262 13028 8318 13030
rect 8342 13028 8398 13030
rect 8422 13028 8478 13030
rect 8182 11994 8238 11996
rect 8262 11994 8318 11996
rect 8342 11994 8398 11996
rect 8422 11994 8478 11996
rect 8182 11942 8208 11994
rect 8208 11942 8238 11994
rect 8262 11942 8272 11994
rect 8272 11942 8318 11994
rect 8342 11942 8388 11994
rect 8388 11942 8398 11994
rect 8422 11942 8452 11994
rect 8452 11942 8478 11994
rect 8182 11940 8238 11942
rect 8262 11940 8318 11942
rect 8342 11940 8398 11942
rect 8422 11940 8478 11942
rect 8182 10906 8238 10908
rect 8262 10906 8318 10908
rect 8342 10906 8398 10908
rect 8422 10906 8478 10908
rect 8182 10854 8208 10906
rect 8208 10854 8238 10906
rect 8262 10854 8272 10906
rect 8272 10854 8318 10906
rect 8342 10854 8388 10906
rect 8388 10854 8398 10906
rect 8422 10854 8452 10906
rect 8452 10854 8478 10906
rect 8182 10852 8238 10854
rect 8262 10852 8318 10854
rect 8342 10852 8398 10854
rect 8422 10852 8478 10854
rect 8182 9818 8238 9820
rect 8262 9818 8318 9820
rect 8342 9818 8398 9820
rect 8422 9818 8478 9820
rect 8182 9766 8208 9818
rect 8208 9766 8238 9818
rect 8262 9766 8272 9818
rect 8272 9766 8318 9818
rect 8342 9766 8388 9818
rect 8388 9766 8398 9818
rect 8422 9766 8452 9818
rect 8452 9766 8478 9818
rect 8182 9764 8238 9766
rect 8262 9764 8318 9766
rect 8342 9764 8398 9766
rect 8422 9764 8478 9766
rect 8182 8730 8238 8732
rect 8262 8730 8318 8732
rect 8342 8730 8398 8732
rect 8422 8730 8478 8732
rect 8182 8678 8208 8730
rect 8208 8678 8238 8730
rect 8262 8678 8272 8730
rect 8272 8678 8318 8730
rect 8342 8678 8388 8730
rect 8388 8678 8398 8730
rect 8422 8678 8452 8730
rect 8452 8678 8478 8730
rect 8182 8676 8238 8678
rect 8262 8676 8318 8678
rect 8342 8676 8398 8678
rect 8422 8676 8478 8678
rect 8182 7642 8238 7644
rect 8262 7642 8318 7644
rect 8342 7642 8398 7644
rect 8422 7642 8478 7644
rect 8182 7590 8208 7642
rect 8208 7590 8238 7642
rect 8262 7590 8272 7642
rect 8272 7590 8318 7642
rect 8342 7590 8388 7642
rect 8388 7590 8398 7642
rect 8422 7590 8452 7642
rect 8452 7590 8478 7642
rect 8182 7588 8238 7590
rect 8262 7588 8318 7590
rect 8342 7588 8398 7590
rect 8422 7588 8478 7590
rect 8182 6554 8238 6556
rect 8262 6554 8318 6556
rect 8342 6554 8398 6556
rect 8422 6554 8478 6556
rect 8182 6502 8208 6554
rect 8208 6502 8238 6554
rect 8262 6502 8272 6554
rect 8272 6502 8318 6554
rect 8342 6502 8388 6554
rect 8388 6502 8398 6554
rect 8422 6502 8452 6554
rect 8452 6502 8478 6554
rect 8182 6500 8238 6502
rect 8262 6500 8318 6502
rect 8342 6500 8398 6502
rect 8422 6500 8478 6502
rect 8182 5466 8238 5468
rect 8262 5466 8318 5468
rect 8342 5466 8398 5468
rect 8422 5466 8478 5468
rect 8182 5414 8208 5466
rect 8208 5414 8238 5466
rect 8262 5414 8272 5466
rect 8272 5414 8318 5466
rect 8342 5414 8388 5466
rect 8388 5414 8398 5466
rect 8422 5414 8452 5466
rect 8452 5414 8478 5466
rect 8182 5412 8238 5414
rect 8262 5412 8318 5414
rect 8342 5412 8398 5414
rect 8422 5412 8478 5414
rect 8182 4378 8238 4380
rect 8262 4378 8318 4380
rect 8342 4378 8398 4380
rect 8422 4378 8478 4380
rect 8182 4326 8208 4378
rect 8208 4326 8238 4378
rect 8262 4326 8272 4378
rect 8272 4326 8318 4378
rect 8342 4326 8388 4378
rect 8388 4326 8398 4378
rect 8422 4326 8452 4378
rect 8452 4326 8478 4378
rect 8182 4324 8238 4326
rect 8262 4324 8318 4326
rect 8342 4324 8398 4326
rect 8422 4324 8478 4326
rect 6737 3834 6793 3836
rect 6817 3834 6873 3836
rect 6897 3834 6953 3836
rect 6977 3834 7033 3836
rect 6737 3782 6763 3834
rect 6763 3782 6793 3834
rect 6817 3782 6827 3834
rect 6827 3782 6873 3834
rect 6897 3782 6943 3834
rect 6943 3782 6953 3834
rect 6977 3782 7007 3834
rect 7007 3782 7033 3834
rect 6737 3780 6793 3782
rect 6817 3780 6873 3782
rect 6897 3780 6953 3782
rect 6977 3780 7033 3782
rect 8182 3290 8238 3292
rect 8262 3290 8318 3292
rect 8342 3290 8398 3292
rect 8422 3290 8478 3292
rect 8182 3238 8208 3290
rect 8208 3238 8238 3290
rect 8262 3238 8272 3290
rect 8272 3238 8318 3290
rect 8342 3238 8388 3290
rect 8388 3238 8398 3290
rect 8422 3238 8452 3290
rect 8452 3238 8478 3290
rect 8182 3236 8238 3238
rect 8262 3236 8318 3238
rect 8342 3236 8398 3238
rect 8422 3236 8478 3238
rect 6737 2746 6793 2748
rect 6817 2746 6873 2748
rect 6897 2746 6953 2748
rect 6977 2746 7033 2748
rect 6737 2694 6763 2746
rect 6763 2694 6793 2746
rect 6817 2694 6827 2746
rect 6827 2694 6873 2746
rect 6897 2694 6943 2746
rect 6943 2694 6953 2746
rect 6977 2694 7007 2746
rect 7007 2694 7033 2746
rect 6737 2692 6793 2694
rect 6817 2692 6873 2694
rect 6897 2692 6953 2694
rect 6977 2692 7033 2694
rect 8574 2624 8630 2680
rect 5292 2202 5348 2204
rect 5372 2202 5428 2204
rect 5452 2202 5508 2204
rect 5532 2202 5588 2204
rect 5292 2150 5318 2202
rect 5318 2150 5348 2202
rect 5372 2150 5382 2202
rect 5382 2150 5428 2202
rect 5452 2150 5498 2202
rect 5498 2150 5508 2202
rect 5532 2150 5562 2202
rect 5562 2150 5588 2202
rect 5292 2148 5348 2150
rect 5372 2148 5428 2150
rect 5452 2148 5508 2150
rect 5532 2148 5588 2150
rect 8182 2202 8238 2204
rect 8262 2202 8318 2204
rect 8342 2202 8398 2204
rect 8422 2202 8478 2204
rect 8182 2150 8208 2202
rect 8208 2150 8238 2202
rect 8262 2150 8272 2202
rect 8272 2150 8318 2202
rect 8342 2150 8388 2202
rect 8388 2150 8398 2202
rect 8422 2150 8452 2202
rect 8452 2150 8478 2202
rect 8182 2148 8238 2150
rect 8262 2148 8318 2150
rect 8342 2148 8398 2150
rect 8422 2148 8478 2150
rect 5078 856 5134 912
<< metal3 >>
rect 6637 23490 6703 23493
rect 10080 23490 10880 23520
rect 6637 23488 10880 23490
rect 6637 23432 6642 23488
rect 6698 23432 10880 23488
rect 6637 23430 10880 23432
rect 6637 23427 6703 23430
rect 10080 23400 10880 23430
rect 3834 22336 4154 22337
rect 3834 22272 3842 22336
rect 3906 22272 3922 22336
rect 3986 22272 4002 22336
rect 4066 22272 4082 22336
rect 4146 22272 4154 22336
rect 3834 22271 4154 22272
rect 6725 22336 7045 22337
rect 6725 22272 6733 22336
rect 6797 22272 6813 22336
rect 6877 22272 6893 22336
rect 6957 22272 6973 22336
rect 7037 22272 7045 22336
rect 6725 22271 7045 22272
rect 2389 21792 2709 21793
rect 2389 21728 2397 21792
rect 2461 21728 2477 21792
rect 2541 21728 2557 21792
rect 2621 21728 2637 21792
rect 2701 21728 2709 21792
rect 2389 21727 2709 21728
rect 5280 21792 5600 21793
rect 5280 21728 5288 21792
rect 5352 21728 5368 21792
rect 5432 21728 5448 21792
rect 5512 21728 5528 21792
rect 5592 21728 5600 21792
rect 5280 21727 5600 21728
rect 8170 21792 8490 21793
rect 8170 21728 8178 21792
rect 8242 21728 8258 21792
rect 8322 21728 8338 21792
rect 8402 21728 8418 21792
rect 8482 21728 8490 21792
rect 8170 21727 8490 21728
rect 7097 21586 7163 21589
rect 10080 21586 10880 21616
rect 7097 21584 10880 21586
rect 7097 21528 7102 21584
rect 7158 21528 10880 21584
rect 7097 21526 10880 21528
rect 7097 21523 7163 21526
rect 10080 21496 10880 21526
rect 3834 21248 4154 21249
rect 3834 21184 3842 21248
rect 3906 21184 3922 21248
rect 3986 21184 4002 21248
rect 4066 21184 4082 21248
rect 4146 21184 4154 21248
rect 3834 21183 4154 21184
rect 6725 21248 7045 21249
rect 6725 21184 6733 21248
rect 6797 21184 6813 21248
rect 6877 21184 6893 21248
rect 6957 21184 6973 21248
rect 7037 21184 7045 21248
rect 6725 21183 7045 21184
rect 2389 20704 2709 20705
rect 2389 20640 2397 20704
rect 2461 20640 2477 20704
rect 2541 20640 2557 20704
rect 2621 20640 2637 20704
rect 2701 20640 2709 20704
rect 2389 20639 2709 20640
rect 5280 20704 5600 20705
rect 5280 20640 5288 20704
rect 5352 20640 5368 20704
rect 5432 20640 5448 20704
rect 5512 20640 5528 20704
rect 5592 20640 5600 20704
rect 5280 20639 5600 20640
rect 8170 20704 8490 20705
rect 8170 20640 8178 20704
rect 8242 20640 8258 20704
rect 8322 20640 8338 20704
rect 8402 20640 8418 20704
rect 8482 20640 8490 20704
rect 8170 20639 8490 20640
rect 0 20498 800 20528
rect 3417 20498 3483 20501
rect 0 20496 3483 20498
rect 0 20440 3422 20496
rect 3478 20440 3483 20496
rect 0 20438 3483 20440
rect 0 20408 800 20438
rect 3417 20435 3483 20438
rect 3834 20160 4154 20161
rect 3834 20096 3842 20160
rect 3906 20096 3922 20160
rect 3986 20096 4002 20160
rect 4066 20096 4082 20160
rect 4146 20096 4154 20160
rect 3834 20095 4154 20096
rect 6725 20160 7045 20161
rect 6725 20096 6733 20160
rect 6797 20096 6813 20160
rect 6877 20096 6893 20160
rect 6957 20096 6973 20160
rect 7037 20096 7045 20160
rect 6725 20095 7045 20096
rect 5625 19818 5691 19821
rect 5625 19816 8770 19818
rect 5625 19760 5630 19816
rect 5686 19760 8770 19816
rect 5625 19758 8770 19760
rect 5625 19755 5691 19758
rect 8710 19682 8770 19758
rect 10080 19682 10880 19712
rect 8710 19622 10880 19682
rect 2389 19616 2709 19617
rect 2389 19552 2397 19616
rect 2461 19552 2477 19616
rect 2541 19552 2557 19616
rect 2621 19552 2637 19616
rect 2701 19552 2709 19616
rect 2389 19551 2709 19552
rect 5280 19616 5600 19617
rect 5280 19552 5288 19616
rect 5352 19552 5368 19616
rect 5432 19552 5448 19616
rect 5512 19552 5528 19616
rect 5592 19552 5600 19616
rect 5280 19551 5600 19552
rect 8170 19616 8490 19617
rect 8170 19552 8178 19616
rect 8242 19552 8258 19616
rect 8322 19552 8338 19616
rect 8402 19552 8418 19616
rect 8482 19552 8490 19616
rect 10080 19592 10880 19622
rect 8170 19551 8490 19552
rect 3834 19072 4154 19073
rect 3834 19008 3842 19072
rect 3906 19008 3922 19072
rect 3986 19008 4002 19072
rect 4066 19008 4082 19072
rect 4146 19008 4154 19072
rect 3834 19007 4154 19008
rect 6725 19072 7045 19073
rect 6725 19008 6733 19072
rect 6797 19008 6813 19072
rect 6877 19008 6893 19072
rect 6957 19008 6973 19072
rect 7037 19008 7045 19072
rect 6725 19007 7045 19008
rect 2389 18528 2709 18529
rect 2389 18464 2397 18528
rect 2461 18464 2477 18528
rect 2541 18464 2557 18528
rect 2621 18464 2637 18528
rect 2701 18464 2709 18528
rect 2389 18463 2709 18464
rect 5280 18528 5600 18529
rect 5280 18464 5288 18528
rect 5352 18464 5368 18528
rect 5432 18464 5448 18528
rect 5512 18464 5528 18528
rect 5592 18464 5600 18528
rect 5280 18463 5600 18464
rect 8170 18528 8490 18529
rect 8170 18464 8178 18528
rect 8242 18464 8258 18528
rect 8322 18464 8338 18528
rect 8402 18464 8418 18528
rect 8482 18464 8490 18528
rect 8170 18463 8490 18464
rect 3834 17984 4154 17985
rect 3834 17920 3842 17984
rect 3906 17920 3922 17984
rect 3986 17920 4002 17984
rect 4066 17920 4082 17984
rect 4146 17920 4154 17984
rect 3834 17919 4154 17920
rect 6725 17984 7045 17985
rect 6725 17920 6733 17984
rect 6797 17920 6813 17984
rect 6877 17920 6893 17984
rect 6957 17920 6973 17984
rect 7037 17920 7045 17984
rect 6725 17919 7045 17920
rect 8201 17778 8267 17781
rect 10080 17778 10880 17808
rect 8201 17776 10880 17778
rect 8201 17720 8206 17776
rect 8262 17720 10880 17776
rect 8201 17718 10880 17720
rect 8201 17715 8267 17718
rect 10080 17688 10880 17718
rect 2389 17440 2709 17441
rect 2389 17376 2397 17440
rect 2461 17376 2477 17440
rect 2541 17376 2557 17440
rect 2621 17376 2637 17440
rect 2701 17376 2709 17440
rect 2389 17375 2709 17376
rect 5280 17440 5600 17441
rect 5280 17376 5288 17440
rect 5352 17376 5368 17440
rect 5432 17376 5448 17440
rect 5512 17376 5528 17440
rect 5592 17376 5600 17440
rect 5280 17375 5600 17376
rect 8170 17440 8490 17441
rect 8170 17376 8178 17440
rect 8242 17376 8258 17440
rect 8322 17376 8338 17440
rect 8402 17376 8418 17440
rect 8482 17376 8490 17440
rect 8170 17375 8490 17376
rect 3834 16896 4154 16897
rect 3834 16832 3842 16896
rect 3906 16832 3922 16896
rect 3986 16832 4002 16896
rect 4066 16832 4082 16896
rect 4146 16832 4154 16896
rect 3834 16831 4154 16832
rect 6725 16896 7045 16897
rect 6725 16832 6733 16896
rect 6797 16832 6813 16896
rect 6877 16832 6893 16896
rect 6957 16832 6973 16896
rect 7037 16832 7045 16896
rect 6725 16831 7045 16832
rect 2389 16352 2709 16353
rect 2389 16288 2397 16352
rect 2461 16288 2477 16352
rect 2541 16288 2557 16352
rect 2621 16288 2637 16352
rect 2701 16288 2709 16352
rect 2389 16287 2709 16288
rect 5280 16352 5600 16353
rect 5280 16288 5288 16352
rect 5352 16288 5368 16352
rect 5432 16288 5448 16352
rect 5512 16288 5528 16352
rect 5592 16288 5600 16352
rect 5280 16287 5600 16288
rect 8170 16352 8490 16353
rect 8170 16288 8178 16352
rect 8242 16288 8258 16352
rect 8322 16288 8338 16352
rect 8402 16288 8418 16352
rect 8482 16288 8490 16352
rect 8170 16287 8490 16288
rect 10080 15874 10880 15904
rect 8158 15814 10880 15874
rect 3834 15808 4154 15809
rect 3834 15744 3842 15808
rect 3906 15744 3922 15808
rect 3986 15744 4002 15808
rect 4066 15744 4082 15808
rect 4146 15744 4154 15808
rect 3834 15743 4154 15744
rect 6725 15808 7045 15809
rect 6725 15744 6733 15808
rect 6797 15744 6813 15808
rect 6877 15744 6893 15808
rect 6957 15744 6973 15808
rect 7037 15744 7045 15808
rect 6725 15743 7045 15744
rect 6453 15602 6519 15605
rect 8158 15602 8218 15814
rect 10080 15784 10880 15814
rect 6453 15600 8218 15602
rect 6453 15544 6458 15600
rect 6514 15544 8218 15600
rect 6453 15542 8218 15544
rect 6453 15539 6519 15542
rect 2389 15264 2709 15265
rect 2389 15200 2397 15264
rect 2461 15200 2477 15264
rect 2541 15200 2557 15264
rect 2621 15200 2637 15264
rect 2701 15200 2709 15264
rect 2389 15199 2709 15200
rect 5280 15264 5600 15265
rect 5280 15200 5288 15264
rect 5352 15200 5368 15264
rect 5432 15200 5448 15264
rect 5512 15200 5528 15264
rect 5592 15200 5600 15264
rect 5280 15199 5600 15200
rect 8170 15264 8490 15265
rect 8170 15200 8178 15264
rect 8242 15200 8258 15264
rect 8322 15200 8338 15264
rect 8402 15200 8418 15264
rect 8482 15200 8490 15264
rect 8170 15199 8490 15200
rect 3834 14720 4154 14721
rect 3834 14656 3842 14720
rect 3906 14656 3922 14720
rect 3986 14656 4002 14720
rect 4066 14656 4082 14720
rect 4146 14656 4154 14720
rect 3834 14655 4154 14656
rect 6725 14720 7045 14721
rect 6725 14656 6733 14720
rect 6797 14656 6813 14720
rect 6877 14656 6893 14720
rect 6957 14656 6973 14720
rect 7037 14656 7045 14720
rect 6725 14655 7045 14656
rect 2389 14176 2709 14177
rect 2389 14112 2397 14176
rect 2461 14112 2477 14176
rect 2541 14112 2557 14176
rect 2621 14112 2637 14176
rect 2701 14112 2709 14176
rect 2389 14111 2709 14112
rect 5280 14176 5600 14177
rect 5280 14112 5288 14176
rect 5352 14112 5368 14176
rect 5432 14112 5448 14176
rect 5512 14112 5528 14176
rect 5592 14112 5600 14176
rect 5280 14111 5600 14112
rect 8170 14176 8490 14177
rect 8170 14112 8178 14176
rect 8242 14112 8258 14176
rect 8322 14112 8338 14176
rect 8402 14112 8418 14176
rect 8482 14112 8490 14176
rect 8170 14111 8490 14112
rect 5625 13970 5691 13973
rect 10080 13970 10880 14000
rect 5625 13968 10880 13970
rect 5625 13912 5630 13968
rect 5686 13912 10880 13968
rect 5625 13910 10880 13912
rect 5625 13907 5691 13910
rect 10080 13880 10880 13910
rect 3834 13632 4154 13633
rect 3834 13568 3842 13632
rect 3906 13568 3922 13632
rect 3986 13568 4002 13632
rect 4066 13568 4082 13632
rect 4146 13568 4154 13632
rect 3834 13567 4154 13568
rect 6725 13632 7045 13633
rect 6725 13568 6733 13632
rect 6797 13568 6813 13632
rect 6877 13568 6893 13632
rect 6957 13568 6973 13632
rect 7037 13568 7045 13632
rect 6725 13567 7045 13568
rect 2389 13088 2709 13089
rect 2389 13024 2397 13088
rect 2461 13024 2477 13088
rect 2541 13024 2557 13088
rect 2621 13024 2637 13088
rect 2701 13024 2709 13088
rect 2389 13023 2709 13024
rect 5280 13088 5600 13089
rect 5280 13024 5288 13088
rect 5352 13024 5368 13088
rect 5432 13024 5448 13088
rect 5512 13024 5528 13088
rect 5592 13024 5600 13088
rect 5280 13023 5600 13024
rect 8170 13088 8490 13089
rect 8170 13024 8178 13088
rect 8242 13024 8258 13088
rect 8322 13024 8338 13088
rect 8402 13024 8418 13088
rect 8482 13024 8490 13088
rect 8170 13023 8490 13024
rect 3834 12544 4154 12545
rect 3834 12480 3842 12544
rect 3906 12480 3922 12544
rect 3986 12480 4002 12544
rect 4066 12480 4082 12544
rect 4146 12480 4154 12544
rect 3834 12479 4154 12480
rect 6725 12544 7045 12545
rect 6725 12480 6733 12544
rect 6797 12480 6813 12544
rect 6877 12480 6893 12544
rect 6957 12480 6973 12544
rect 7037 12480 7045 12544
rect 6725 12479 7045 12480
rect 0 12338 800 12368
rect 2865 12338 2931 12341
rect 0 12336 2931 12338
rect 0 12280 2870 12336
rect 2926 12280 2931 12336
rect 0 12278 2931 12280
rect 0 12248 800 12278
rect 2865 12275 2931 12278
rect 5625 12202 5691 12205
rect 10080 12202 10880 12232
rect 5625 12200 10880 12202
rect 5625 12144 5630 12200
rect 5686 12144 10880 12200
rect 5625 12142 10880 12144
rect 5625 12139 5691 12142
rect 10080 12112 10880 12142
rect 2389 12000 2709 12001
rect 2389 11936 2397 12000
rect 2461 11936 2477 12000
rect 2541 11936 2557 12000
rect 2621 11936 2637 12000
rect 2701 11936 2709 12000
rect 2389 11935 2709 11936
rect 5280 12000 5600 12001
rect 5280 11936 5288 12000
rect 5352 11936 5368 12000
rect 5432 11936 5448 12000
rect 5512 11936 5528 12000
rect 5592 11936 5600 12000
rect 5280 11935 5600 11936
rect 8170 12000 8490 12001
rect 8170 11936 8178 12000
rect 8242 11936 8258 12000
rect 8322 11936 8338 12000
rect 8402 11936 8418 12000
rect 8482 11936 8490 12000
rect 8170 11935 8490 11936
rect 3834 11456 4154 11457
rect 3834 11392 3842 11456
rect 3906 11392 3922 11456
rect 3986 11392 4002 11456
rect 4066 11392 4082 11456
rect 4146 11392 4154 11456
rect 3834 11391 4154 11392
rect 6725 11456 7045 11457
rect 6725 11392 6733 11456
rect 6797 11392 6813 11456
rect 6877 11392 6893 11456
rect 6957 11392 6973 11456
rect 7037 11392 7045 11456
rect 6725 11391 7045 11392
rect 2389 10912 2709 10913
rect 2389 10848 2397 10912
rect 2461 10848 2477 10912
rect 2541 10848 2557 10912
rect 2621 10848 2637 10912
rect 2701 10848 2709 10912
rect 2389 10847 2709 10848
rect 5280 10912 5600 10913
rect 5280 10848 5288 10912
rect 5352 10848 5368 10912
rect 5432 10848 5448 10912
rect 5512 10848 5528 10912
rect 5592 10848 5600 10912
rect 5280 10847 5600 10848
rect 8170 10912 8490 10913
rect 8170 10848 8178 10912
rect 8242 10848 8258 10912
rect 8322 10848 8338 10912
rect 8402 10848 8418 10912
rect 8482 10848 8490 10912
rect 8170 10847 8490 10848
rect 6545 10570 6611 10573
rect 6545 10568 8218 10570
rect 6545 10512 6550 10568
rect 6606 10512 8218 10568
rect 6545 10510 8218 10512
rect 6545 10507 6611 10510
rect 3834 10368 4154 10369
rect 3834 10304 3842 10368
rect 3906 10304 3922 10368
rect 3986 10304 4002 10368
rect 4066 10304 4082 10368
rect 4146 10304 4154 10368
rect 3834 10303 4154 10304
rect 6725 10368 7045 10369
rect 6725 10304 6733 10368
rect 6797 10304 6813 10368
rect 6877 10304 6893 10368
rect 6957 10304 6973 10368
rect 7037 10304 7045 10368
rect 6725 10303 7045 10304
rect 8158 10298 8218 10510
rect 10080 10298 10880 10328
rect 8158 10238 10880 10298
rect 10080 10208 10880 10238
rect 2389 9824 2709 9825
rect 2389 9760 2397 9824
rect 2461 9760 2477 9824
rect 2541 9760 2557 9824
rect 2621 9760 2637 9824
rect 2701 9760 2709 9824
rect 2389 9759 2709 9760
rect 5280 9824 5600 9825
rect 5280 9760 5288 9824
rect 5352 9760 5368 9824
rect 5432 9760 5448 9824
rect 5512 9760 5528 9824
rect 5592 9760 5600 9824
rect 5280 9759 5600 9760
rect 8170 9824 8490 9825
rect 8170 9760 8178 9824
rect 8242 9760 8258 9824
rect 8322 9760 8338 9824
rect 8402 9760 8418 9824
rect 8482 9760 8490 9824
rect 8170 9759 8490 9760
rect 3834 9280 4154 9281
rect 3834 9216 3842 9280
rect 3906 9216 3922 9280
rect 3986 9216 4002 9280
rect 4066 9216 4082 9280
rect 4146 9216 4154 9280
rect 3834 9215 4154 9216
rect 6725 9280 7045 9281
rect 6725 9216 6733 9280
rect 6797 9216 6813 9280
rect 6877 9216 6893 9280
rect 6957 9216 6973 9280
rect 7037 9216 7045 9280
rect 6725 9215 7045 9216
rect 2389 8736 2709 8737
rect 2389 8672 2397 8736
rect 2461 8672 2477 8736
rect 2541 8672 2557 8736
rect 2621 8672 2637 8736
rect 2701 8672 2709 8736
rect 2389 8671 2709 8672
rect 5280 8736 5600 8737
rect 5280 8672 5288 8736
rect 5352 8672 5368 8736
rect 5432 8672 5448 8736
rect 5512 8672 5528 8736
rect 5592 8672 5600 8736
rect 5280 8671 5600 8672
rect 8170 8736 8490 8737
rect 8170 8672 8178 8736
rect 8242 8672 8258 8736
rect 8322 8672 8338 8736
rect 8402 8672 8418 8736
rect 8482 8672 8490 8736
rect 8170 8671 8490 8672
rect 6637 8394 6703 8397
rect 10080 8394 10880 8424
rect 6637 8392 10880 8394
rect 6637 8336 6642 8392
rect 6698 8336 10880 8392
rect 6637 8334 10880 8336
rect 6637 8331 6703 8334
rect 10080 8304 10880 8334
rect 3834 8192 4154 8193
rect 3834 8128 3842 8192
rect 3906 8128 3922 8192
rect 3986 8128 4002 8192
rect 4066 8128 4082 8192
rect 4146 8128 4154 8192
rect 3834 8127 4154 8128
rect 6725 8192 7045 8193
rect 6725 8128 6733 8192
rect 6797 8128 6813 8192
rect 6877 8128 6893 8192
rect 6957 8128 6973 8192
rect 7037 8128 7045 8192
rect 6725 8127 7045 8128
rect 2389 7648 2709 7649
rect 2389 7584 2397 7648
rect 2461 7584 2477 7648
rect 2541 7584 2557 7648
rect 2621 7584 2637 7648
rect 2701 7584 2709 7648
rect 2389 7583 2709 7584
rect 5280 7648 5600 7649
rect 5280 7584 5288 7648
rect 5352 7584 5368 7648
rect 5432 7584 5448 7648
rect 5512 7584 5528 7648
rect 5592 7584 5600 7648
rect 5280 7583 5600 7584
rect 8170 7648 8490 7649
rect 8170 7584 8178 7648
rect 8242 7584 8258 7648
rect 8322 7584 8338 7648
rect 8402 7584 8418 7648
rect 8482 7584 8490 7648
rect 8170 7583 8490 7584
rect 3834 7104 4154 7105
rect 3834 7040 3842 7104
rect 3906 7040 3922 7104
rect 3986 7040 4002 7104
rect 4066 7040 4082 7104
rect 4146 7040 4154 7104
rect 3834 7039 4154 7040
rect 6725 7104 7045 7105
rect 6725 7040 6733 7104
rect 6797 7040 6813 7104
rect 6877 7040 6893 7104
rect 6957 7040 6973 7104
rect 7037 7040 7045 7104
rect 6725 7039 7045 7040
rect 6177 6762 6243 6765
rect 6177 6760 8770 6762
rect 6177 6704 6182 6760
rect 6238 6704 8770 6760
rect 6177 6702 8770 6704
rect 6177 6699 6243 6702
rect 2389 6560 2709 6561
rect 2389 6496 2397 6560
rect 2461 6496 2477 6560
rect 2541 6496 2557 6560
rect 2621 6496 2637 6560
rect 2701 6496 2709 6560
rect 2389 6495 2709 6496
rect 5280 6560 5600 6561
rect 5280 6496 5288 6560
rect 5352 6496 5368 6560
rect 5432 6496 5448 6560
rect 5512 6496 5528 6560
rect 5592 6496 5600 6560
rect 5280 6495 5600 6496
rect 8170 6560 8490 6561
rect 8170 6496 8178 6560
rect 8242 6496 8258 6560
rect 8322 6496 8338 6560
rect 8402 6496 8418 6560
rect 8482 6496 8490 6560
rect 8170 6495 8490 6496
rect 8710 6490 8770 6702
rect 10080 6490 10880 6520
rect 8710 6430 10880 6490
rect 10080 6400 10880 6430
rect 3834 6016 4154 6017
rect 3834 5952 3842 6016
rect 3906 5952 3922 6016
rect 3986 5952 4002 6016
rect 4066 5952 4082 6016
rect 4146 5952 4154 6016
rect 3834 5951 4154 5952
rect 6725 6016 7045 6017
rect 6725 5952 6733 6016
rect 6797 5952 6813 6016
rect 6877 5952 6893 6016
rect 6957 5952 6973 6016
rect 7037 5952 7045 6016
rect 6725 5951 7045 5952
rect 2389 5472 2709 5473
rect 2389 5408 2397 5472
rect 2461 5408 2477 5472
rect 2541 5408 2557 5472
rect 2621 5408 2637 5472
rect 2701 5408 2709 5472
rect 2389 5407 2709 5408
rect 5280 5472 5600 5473
rect 5280 5408 5288 5472
rect 5352 5408 5368 5472
rect 5432 5408 5448 5472
rect 5512 5408 5528 5472
rect 5592 5408 5600 5472
rect 5280 5407 5600 5408
rect 8170 5472 8490 5473
rect 8170 5408 8178 5472
rect 8242 5408 8258 5472
rect 8322 5408 8338 5472
rect 8402 5408 8418 5472
rect 8482 5408 8490 5472
rect 8170 5407 8490 5408
rect 3834 4928 4154 4929
rect 3834 4864 3842 4928
rect 3906 4864 3922 4928
rect 3986 4864 4002 4928
rect 4066 4864 4082 4928
rect 4146 4864 4154 4928
rect 3834 4863 4154 4864
rect 6725 4928 7045 4929
rect 6725 4864 6733 4928
rect 6797 4864 6813 4928
rect 6877 4864 6893 4928
rect 6957 4864 6973 4928
rect 7037 4864 7045 4928
rect 6725 4863 7045 4864
rect 5625 4586 5691 4589
rect 10080 4586 10880 4616
rect 5625 4584 10880 4586
rect 5625 4528 5630 4584
rect 5686 4528 10880 4584
rect 5625 4526 10880 4528
rect 5625 4523 5691 4526
rect 10080 4496 10880 4526
rect 2389 4384 2709 4385
rect 2389 4320 2397 4384
rect 2461 4320 2477 4384
rect 2541 4320 2557 4384
rect 2621 4320 2637 4384
rect 2701 4320 2709 4384
rect 2389 4319 2709 4320
rect 5280 4384 5600 4385
rect 5280 4320 5288 4384
rect 5352 4320 5368 4384
rect 5432 4320 5448 4384
rect 5512 4320 5528 4384
rect 5592 4320 5600 4384
rect 5280 4319 5600 4320
rect 8170 4384 8490 4385
rect 8170 4320 8178 4384
rect 8242 4320 8258 4384
rect 8322 4320 8338 4384
rect 8402 4320 8418 4384
rect 8482 4320 8490 4384
rect 8170 4319 8490 4320
rect 0 4178 800 4208
rect 3325 4178 3391 4181
rect 0 4176 3391 4178
rect 0 4120 3330 4176
rect 3386 4120 3391 4176
rect 0 4118 3391 4120
rect 0 4088 800 4118
rect 3325 4115 3391 4118
rect 3834 3840 4154 3841
rect 3834 3776 3842 3840
rect 3906 3776 3922 3840
rect 3986 3776 4002 3840
rect 4066 3776 4082 3840
rect 4146 3776 4154 3840
rect 3834 3775 4154 3776
rect 6725 3840 7045 3841
rect 6725 3776 6733 3840
rect 6797 3776 6813 3840
rect 6877 3776 6893 3840
rect 6957 3776 6973 3840
rect 7037 3776 7045 3840
rect 6725 3775 7045 3776
rect 2389 3296 2709 3297
rect 2389 3232 2397 3296
rect 2461 3232 2477 3296
rect 2541 3232 2557 3296
rect 2621 3232 2637 3296
rect 2701 3232 2709 3296
rect 2389 3231 2709 3232
rect 5280 3296 5600 3297
rect 5280 3232 5288 3296
rect 5352 3232 5368 3296
rect 5432 3232 5448 3296
rect 5512 3232 5528 3296
rect 5592 3232 5600 3296
rect 5280 3231 5600 3232
rect 8170 3296 8490 3297
rect 8170 3232 8178 3296
rect 8242 3232 8258 3296
rect 8322 3232 8338 3296
rect 8402 3232 8418 3296
rect 8482 3232 8490 3296
rect 8170 3231 8490 3232
rect 3834 2752 4154 2753
rect 3834 2688 3842 2752
rect 3906 2688 3922 2752
rect 3986 2688 4002 2752
rect 4066 2688 4082 2752
rect 4146 2688 4154 2752
rect 3834 2687 4154 2688
rect 6725 2752 7045 2753
rect 6725 2688 6733 2752
rect 6797 2688 6813 2752
rect 6877 2688 6893 2752
rect 6957 2688 6973 2752
rect 7037 2688 7045 2752
rect 6725 2687 7045 2688
rect 8569 2682 8635 2685
rect 10080 2682 10880 2712
rect 8569 2680 10880 2682
rect 8569 2624 8574 2680
rect 8630 2624 10880 2680
rect 8569 2622 10880 2624
rect 8569 2619 8635 2622
rect 10080 2592 10880 2622
rect 2389 2208 2709 2209
rect 2389 2144 2397 2208
rect 2461 2144 2477 2208
rect 2541 2144 2557 2208
rect 2621 2144 2637 2208
rect 2701 2144 2709 2208
rect 2389 2143 2709 2144
rect 5280 2208 5600 2209
rect 5280 2144 5288 2208
rect 5352 2144 5368 2208
rect 5432 2144 5448 2208
rect 5512 2144 5528 2208
rect 5592 2144 5600 2208
rect 5280 2143 5600 2144
rect 8170 2208 8490 2209
rect 8170 2144 8178 2208
rect 8242 2144 8258 2208
rect 8322 2144 8338 2208
rect 8402 2144 8418 2208
rect 8482 2144 8490 2208
rect 8170 2143 8490 2144
rect 5073 914 5139 917
rect 10080 914 10880 944
rect 5073 912 10880 914
rect 5073 856 5078 912
rect 5134 856 10880 912
rect 5073 854 10880 856
rect 5073 851 5139 854
rect 10080 824 10880 854
<< via3 >>
rect 3842 22332 3906 22336
rect 3842 22276 3846 22332
rect 3846 22276 3902 22332
rect 3902 22276 3906 22332
rect 3842 22272 3906 22276
rect 3922 22332 3986 22336
rect 3922 22276 3926 22332
rect 3926 22276 3982 22332
rect 3982 22276 3986 22332
rect 3922 22272 3986 22276
rect 4002 22332 4066 22336
rect 4002 22276 4006 22332
rect 4006 22276 4062 22332
rect 4062 22276 4066 22332
rect 4002 22272 4066 22276
rect 4082 22332 4146 22336
rect 4082 22276 4086 22332
rect 4086 22276 4142 22332
rect 4142 22276 4146 22332
rect 4082 22272 4146 22276
rect 6733 22332 6797 22336
rect 6733 22276 6737 22332
rect 6737 22276 6793 22332
rect 6793 22276 6797 22332
rect 6733 22272 6797 22276
rect 6813 22332 6877 22336
rect 6813 22276 6817 22332
rect 6817 22276 6873 22332
rect 6873 22276 6877 22332
rect 6813 22272 6877 22276
rect 6893 22332 6957 22336
rect 6893 22276 6897 22332
rect 6897 22276 6953 22332
rect 6953 22276 6957 22332
rect 6893 22272 6957 22276
rect 6973 22332 7037 22336
rect 6973 22276 6977 22332
rect 6977 22276 7033 22332
rect 7033 22276 7037 22332
rect 6973 22272 7037 22276
rect 2397 21788 2461 21792
rect 2397 21732 2401 21788
rect 2401 21732 2457 21788
rect 2457 21732 2461 21788
rect 2397 21728 2461 21732
rect 2477 21788 2541 21792
rect 2477 21732 2481 21788
rect 2481 21732 2537 21788
rect 2537 21732 2541 21788
rect 2477 21728 2541 21732
rect 2557 21788 2621 21792
rect 2557 21732 2561 21788
rect 2561 21732 2617 21788
rect 2617 21732 2621 21788
rect 2557 21728 2621 21732
rect 2637 21788 2701 21792
rect 2637 21732 2641 21788
rect 2641 21732 2697 21788
rect 2697 21732 2701 21788
rect 2637 21728 2701 21732
rect 5288 21788 5352 21792
rect 5288 21732 5292 21788
rect 5292 21732 5348 21788
rect 5348 21732 5352 21788
rect 5288 21728 5352 21732
rect 5368 21788 5432 21792
rect 5368 21732 5372 21788
rect 5372 21732 5428 21788
rect 5428 21732 5432 21788
rect 5368 21728 5432 21732
rect 5448 21788 5512 21792
rect 5448 21732 5452 21788
rect 5452 21732 5508 21788
rect 5508 21732 5512 21788
rect 5448 21728 5512 21732
rect 5528 21788 5592 21792
rect 5528 21732 5532 21788
rect 5532 21732 5588 21788
rect 5588 21732 5592 21788
rect 5528 21728 5592 21732
rect 8178 21788 8242 21792
rect 8178 21732 8182 21788
rect 8182 21732 8238 21788
rect 8238 21732 8242 21788
rect 8178 21728 8242 21732
rect 8258 21788 8322 21792
rect 8258 21732 8262 21788
rect 8262 21732 8318 21788
rect 8318 21732 8322 21788
rect 8258 21728 8322 21732
rect 8338 21788 8402 21792
rect 8338 21732 8342 21788
rect 8342 21732 8398 21788
rect 8398 21732 8402 21788
rect 8338 21728 8402 21732
rect 8418 21788 8482 21792
rect 8418 21732 8422 21788
rect 8422 21732 8478 21788
rect 8478 21732 8482 21788
rect 8418 21728 8482 21732
rect 3842 21244 3906 21248
rect 3842 21188 3846 21244
rect 3846 21188 3902 21244
rect 3902 21188 3906 21244
rect 3842 21184 3906 21188
rect 3922 21244 3986 21248
rect 3922 21188 3926 21244
rect 3926 21188 3982 21244
rect 3982 21188 3986 21244
rect 3922 21184 3986 21188
rect 4002 21244 4066 21248
rect 4002 21188 4006 21244
rect 4006 21188 4062 21244
rect 4062 21188 4066 21244
rect 4002 21184 4066 21188
rect 4082 21244 4146 21248
rect 4082 21188 4086 21244
rect 4086 21188 4142 21244
rect 4142 21188 4146 21244
rect 4082 21184 4146 21188
rect 6733 21244 6797 21248
rect 6733 21188 6737 21244
rect 6737 21188 6793 21244
rect 6793 21188 6797 21244
rect 6733 21184 6797 21188
rect 6813 21244 6877 21248
rect 6813 21188 6817 21244
rect 6817 21188 6873 21244
rect 6873 21188 6877 21244
rect 6813 21184 6877 21188
rect 6893 21244 6957 21248
rect 6893 21188 6897 21244
rect 6897 21188 6953 21244
rect 6953 21188 6957 21244
rect 6893 21184 6957 21188
rect 6973 21244 7037 21248
rect 6973 21188 6977 21244
rect 6977 21188 7033 21244
rect 7033 21188 7037 21244
rect 6973 21184 7037 21188
rect 2397 20700 2461 20704
rect 2397 20644 2401 20700
rect 2401 20644 2457 20700
rect 2457 20644 2461 20700
rect 2397 20640 2461 20644
rect 2477 20700 2541 20704
rect 2477 20644 2481 20700
rect 2481 20644 2537 20700
rect 2537 20644 2541 20700
rect 2477 20640 2541 20644
rect 2557 20700 2621 20704
rect 2557 20644 2561 20700
rect 2561 20644 2617 20700
rect 2617 20644 2621 20700
rect 2557 20640 2621 20644
rect 2637 20700 2701 20704
rect 2637 20644 2641 20700
rect 2641 20644 2697 20700
rect 2697 20644 2701 20700
rect 2637 20640 2701 20644
rect 5288 20700 5352 20704
rect 5288 20644 5292 20700
rect 5292 20644 5348 20700
rect 5348 20644 5352 20700
rect 5288 20640 5352 20644
rect 5368 20700 5432 20704
rect 5368 20644 5372 20700
rect 5372 20644 5428 20700
rect 5428 20644 5432 20700
rect 5368 20640 5432 20644
rect 5448 20700 5512 20704
rect 5448 20644 5452 20700
rect 5452 20644 5508 20700
rect 5508 20644 5512 20700
rect 5448 20640 5512 20644
rect 5528 20700 5592 20704
rect 5528 20644 5532 20700
rect 5532 20644 5588 20700
rect 5588 20644 5592 20700
rect 5528 20640 5592 20644
rect 8178 20700 8242 20704
rect 8178 20644 8182 20700
rect 8182 20644 8238 20700
rect 8238 20644 8242 20700
rect 8178 20640 8242 20644
rect 8258 20700 8322 20704
rect 8258 20644 8262 20700
rect 8262 20644 8318 20700
rect 8318 20644 8322 20700
rect 8258 20640 8322 20644
rect 8338 20700 8402 20704
rect 8338 20644 8342 20700
rect 8342 20644 8398 20700
rect 8398 20644 8402 20700
rect 8338 20640 8402 20644
rect 8418 20700 8482 20704
rect 8418 20644 8422 20700
rect 8422 20644 8478 20700
rect 8478 20644 8482 20700
rect 8418 20640 8482 20644
rect 3842 20156 3906 20160
rect 3842 20100 3846 20156
rect 3846 20100 3902 20156
rect 3902 20100 3906 20156
rect 3842 20096 3906 20100
rect 3922 20156 3986 20160
rect 3922 20100 3926 20156
rect 3926 20100 3982 20156
rect 3982 20100 3986 20156
rect 3922 20096 3986 20100
rect 4002 20156 4066 20160
rect 4002 20100 4006 20156
rect 4006 20100 4062 20156
rect 4062 20100 4066 20156
rect 4002 20096 4066 20100
rect 4082 20156 4146 20160
rect 4082 20100 4086 20156
rect 4086 20100 4142 20156
rect 4142 20100 4146 20156
rect 4082 20096 4146 20100
rect 6733 20156 6797 20160
rect 6733 20100 6737 20156
rect 6737 20100 6793 20156
rect 6793 20100 6797 20156
rect 6733 20096 6797 20100
rect 6813 20156 6877 20160
rect 6813 20100 6817 20156
rect 6817 20100 6873 20156
rect 6873 20100 6877 20156
rect 6813 20096 6877 20100
rect 6893 20156 6957 20160
rect 6893 20100 6897 20156
rect 6897 20100 6953 20156
rect 6953 20100 6957 20156
rect 6893 20096 6957 20100
rect 6973 20156 7037 20160
rect 6973 20100 6977 20156
rect 6977 20100 7033 20156
rect 7033 20100 7037 20156
rect 6973 20096 7037 20100
rect 2397 19612 2461 19616
rect 2397 19556 2401 19612
rect 2401 19556 2457 19612
rect 2457 19556 2461 19612
rect 2397 19552 2461 19556
rect 2477 19612 2541 19616
rect 2477 19556 2481 19612
rect 2481 19556 2537 19612
rect 2537 19556 2541 19612
rect 2477 19552 2541 19556
rect 2557 19612 2621 19616
rect 2557 19556 2561 19612
rect 2561 19556 2617 19612
rect 2617 19556 2621 19612
rect 2557 19552 2621 19556
rect 2637 19612 2701 19616
rect 2637 19556 2641 19612
rect 2641 19556 2697 19612
rect 2697 19556 2701 19612
rect 2637 19552 2701 19556
rect 5288 19612 5352 19616
rect 5288 19556 5292 19612
rect 5292 19556 5348 19612
rect 5348 19556 5352 19612
rect 5288 19552 5352 19556
rect 5368 19612 5432 19616
rect 5368 19556 5372 19612
rect 5372 19556 5428 19612
rect 5428 19556 5432 19612
rect 5368 19552 5432 19556
rect 5448 19612 5512 19616
rect 5448 19556 5452 19612
rect 5452 19556 5508 19612
rect 5508 19556 5512 19612
rect 5448 19552 5512 19556
rect 5528 19612 5592 19616
rect 5528 19556 5532 19612
rect 5532 19556 5588 19612
rect 5588 19556 5592 19612
rect 5528 19552 5592 19556
rect 8178 19612 8242 19616
rect 8178 19556 8182 19612
rect 8182 19556 8238 19612
rect 8238 19556 8242 19612
rect 8178 19552 8242 19556
rect 8258 19612 8322 19616
rect 8258 19556 8262 19612
rect 8262 19556 8318 19612
rect 8318 19556 8322 19612
rect 8258 19552 8322 19556
rect 8338 19612 8402 19616
rect 8338 19556 8342 19612
rect 8342 19556 8398 19612
rect 8398 19556 8402 19612
rect 8338 19552 8402 19556
rect 8418 19612 8482 19616
rect 8418 19556 8422 19612
rect 8422 19556 8478 19612
rect 8478 19556 8482 19612
rect 8418 19552 8482 19556
rect 3842 19068 3906 19072
rect 3842 19012 3846 19068
rect 3846 19012 3902 19068
rect 3902 19012 3906 19068
rect 3842 19008 3906 19012
rect 3922 19068 3986 19072
rect 3922 19012 3926 19068
rect 3926 19012 3982 19068
rect 3982 19012 3986 19068
rect 3922 19008 3986 19012
rect 4002 19068 4066 19072
rect 4002 19012 4006 19068
rect 4006 19012 4062 19068
rect 4062 19012 4066 19068
rect 4002 19008 4066 19012
rect 4082 19068 4146 19072
rect 4082 19012 4086 19068
rect 4086 19012 4142 19068
rect 4142 19012 4146 19068
rect 4082 19008 4146 19012
rect 6733 19068 6797 19072
rect 6733 19012 6737 19068
rect 6737 19012 6793 19068
rect 6793 19012 6797 19068
rect 6733 19008 6797 19012
rect 6813 19068 6877 19072
rect 6813 19012 6817 19068
rect 6817 19012 6873 19068
rect 6873 19012 6877 19068
rect 6813 19008 6877 19012
rect 6893 19068 6957 19072
rect 6893 19012 6897 19068
rect 6897 19012 6953 19068
rect 6953 19012 6957 19068
rect 6893 19008 6957 19012
rect 6973 19068 7037 19072
rect 6973 19012 6977 19068
rect 6977 19012 7033 19068
rect 7033 19012 7037 19068
rect 6973 19008 7037 19012
rect 2397 18524 2461 18528
rect 2397 18468 2401 18524
rect 2401 18468 2457 18524
rect 2457 18468 2461 18524
rect 2397 18464 2461 18468
rect 2477 18524 2541 18528
rect 2477 18468 2481 18524
rect 2481 18468 2537 18524
rect 2537 18468 2541 18524
rect 2477 18464 2541 18468
rect 2557 18524 2621 18528
rect 2557 18468 2561 18524
rect 2561 18468 2617 18524
rect 2617 18468 2621 18524
rect 2557 18464 2621 18468
rect 2637 18524 2701 18528
rect 2637 18468 2641 18524
rect 2641 18468 2697 18524
rect 2697 18468 2701 18524
rect 2637 18464 2701 18468
rect 5288 18524 5352 18528
rect 5288 18468 5292 18524
rect 5292 18468 5348 18524
rect 5348 18468 5352 18524
rect 5288 18464 5352 18468
rect 5368 18524 5432 18528
rect 5368 18468 5372 18524
rect 5372 18468 5428 18524
rect 5428 18468 5432 18524
rect 5368 18464 5432 18468
rect 5448 18524 5512 18528
rect 5448 18468 5452 18524
rect 5452 18468 5508 18524
rect 5508 18468 5512 18524
rect 5448 18464 5512 18468
rect 5528 18524 5592 18528
rect 5528 18468 5532 18524
rect 5532 18468 5588 18524
rect 5588 18468 5592 18524
rect 5528 18464 5592 18468
rect 8178 18524 8242 18528
rect 8178 18468 8182 18524
rect 8182 18468 8238 18524
rect 8238 18468 8242 18524
rect 8178 18464 8242 18468
rect 8258 18524 8322 18528
rect 8258 18468 8262 18524
rect 8262 18468 8318 18524
rect 8318 18468 8322 18524
rect 8258 18464 8322 18468
rect 8338 18524 8402 18528
rect 8338 18468 8342 18524
rect 8342 18468 8398 18524
rect 8398 18468 8402 18524
rect 8338 18464 8402 18468
rect 8418 18524 8482 18528
rect 8418 18468 8422 18524
rect 8422 18468 8478 18524
rect 8478 18468 8482 18524
rect 8418 18464 8482 18468
rect 3842 17980 3906 17984
rect 3842 17924 3846 17980
rect 3846 17924 3902 17980
rect 3902 17924 3906 17980
rect 3842 17920 3906 17924
rect 3922 17980 3986 17984
rect 3922 17924 3926 17980
rect 3926 17924 3982 17980
rect 3982 17924 3986 17980
rect 3922 17920 3986 17924
rect 4002 17980 4066 17984
rect 4002 17924 4006 17980
rect 4006 17924 4062 17980
rect 4062 17924 4066 17980
rect 4002 17920 4066 17924
rect 4082 17980 4146 17984
rect 4082 17924 4086 17980
rect 4086 17924 4142 17980
rect 4142 17924 4146 17980
rect 4082 17920 4146 17924
rect 6733 17980 6797 17984
rect 6733 17924 6737 17980
rect 6737 17924 6793 17980
rect 6793 17924 6797 17980
rect 6733 17920 6797 17924
rect 6813 17980 6877 17984
rect 6813 17924 6817 17980
rect 6817 17924 6873 17980
rect 6873 17924 6877 17980
rect 6813 17920 6877 17924
rect 6893 17980 6957 17984
rect 6893 17924 6897 17980
rect 6897 17924 6953 17980
rect 6953 17924 6957 17980
rect 6893 17920 6957 17924
rect 6973 17980 7037 17984
rect 6973 17924 6977 17980
rect 6977 17924 7033 17980
rect 7033 17924 7037 17980
rect 6973 17920 7037 17924
rect 2397 17436 2461 17440
rect 2397 17380 2401 17436
rect 2401 17380 2457 17436
rect 2457 17380 2461 17436
rect 2397 17376 2461 17380
rect 2477 17436 2541 17440
rect 2477 17380 2481 17436
rect 2481 17380 2537 17436
rect 2537 17380 2541 17436
rect 2477 17376 2541 17380
rect 2557 17436 2621 17440
rect 2557 17380 2561 17436
rect 2561 17380 2617 17436
rect 2617 17380 2621 17436
rect 2557 17376 2621 17380
rect 2637 17436 2701 17440
rect 2637 17380 2641 17436
rect 2641 17380 2697 17436
rect 2697 17380 2701 17436
rect 2637 17376 2701 17380
rect 5288 17436 5352 17440
rect 5288 17380 5292 17436
rect 5292 17380 5348 17436
rect 5348 17380 5352 17436
rect 5288 17376 5352 17380
rect 5368 17436 5432 17440
rect 5368 17380 5372 17436
rect 5372 17380 5428 17436
rect 5428 17380 5432 17436
rect 5368 17376 5432 17380
rect 5448 17436 5512 17440
rect 5448 17380 5452 17436
rect 5452 17380 5508 17436
rect 5508 17380 5512 17436
rect 5448 17376 5512 17380
rect 5528 17436 5592 17440
rect 5528 17380 5532 17436
rect 5532 17380 5588 17436
rect 5588 17380 5592 17436
rect 5528 17376 5592 17380
rect 8178 17436 8242 17440
rect 8178 17380 8182 17436
rect 8182 17380 8238 17436
rect 8238 17380 8242 17436
rect 8178 17376 8242 17380
rect 8258 17436 8322 17440
rect 8258 17380 8262 17436
rect 8262 17380 8318 17436
rect 8318 17380 8322 17436
rect 8258 17376 8322 17380
rect 8338 17436 8402 17440
rect 8338 17380 8342 17436
rect 8342 17380 8398 17436
rect 8398 17380 8402 17436
rect 8338 17376 8402 17380
rect 8418 17436 8482 17440
rect 8418 17380 8422 17436
rect 8422 17380 8478 17436
rect 8478 17380 8482 17436
rect 8418 17376 8482 17380
rect 3842 16892 3906 16896
rect 3842 16836 3846 16892
rect 3846 16836 3902 16892
rect 3902 16836 3906 16892
rect 3842 16832 3906 16836
rect 3922 16892 3986 16896
rect 3922 16836 3926 16892
rect 3926 16836 3982 16892
rect 3982 16836 3986 16892
rect 3922 16832 3986 16836
rect 4002 16892 4066 16896
rect 4002 16836 4006 16892
rect 4006 16836 4062 16892
rect 4062 16836 4066 16892
rect 4002 16832 4066 16836
rect 4082 16892 4146 16896
rect 4082 16836 4086 16892
rect 4086 16836 4142 16892
rect 4142 16836 4146 16892
rect 4082 16832 4146 16836
rect 6733 16892 6797 16896
rect 6733 16836 6737 16892
rect 6737 16836 6793 16892
rect 6793 16836 6797 16892
rect 6733 16832 6797 16836
rect 6813 16892 6877 16896
rect 6813 16836 6817 16892
rect 6817 16836 6873 16892
rect 6873 16836 6877 16892
rect 6813 16832 6877 16836
rect 6893 16892 6957 16896
rect 6893 16836 6897 16892
rect 6897 16836 6953 16892
rect 6953 16836 6957 16892
rect 6893 16832 6957 16836
rect 6973 16892 7037 16896
rect 6973 16836 6977 16892
rect 6977 16836 7033 16892
rect 7033 16836 7037 16892
rect 6973 16832 7037 16836
rect 2397 16348 2461 16352
rect 2397 16292 2401 16348
rect 2401 16292 2457 16348
rect 2457 16292 2461 16348
rect 2397 16288 2461 16292
rect 2477 16348 2541 16352
rect 2477 16292 2481 16348
rect 2481 16292 2537 16348
rect 2537 16292 2541 16348
rect 2477 16288 2541 16292
rect 2557 16348 2621 16352
rect 2557 16292 2561 16348
rect 2561 16292 2617 16348
rect 2617 16292 2621 16348
rect 2557 16288 2621 16292
rect 2637 16348 2701 16352
rect 2637 16292 2641 16348
rect 2641 16292 2697 16348
rect 2697 16292 2701 16348
rect 2637 16288 2701 16292
rect 5288 16348 5352 16352
rect 5288 16292 5292 16348
rect 5292 16292 5348 16348
rect 5348 16292 5352 16348
rect 5288 16288 5352 16292
rect 5368 16348 5432 16352
rect 5368 16292 5372 16348
rect 5372 16292 5428 16348
rect 5428 16292 5432 16348
rect 5368 16288 5432 16292
rect 5448 16348 5512 16352
rect 5448 16292 5452 16348
rect 5452 16292 5508 16348
rect 5508 16292 5512 16348
rect 5448 16288 5512 16292
rect 5528 16348 5592 16352
rect 5528 16292 5532 16348
rect 5532 16292 5588 16348
rect 5588 16292 5592 16348
rect 5528 16288 5592 16292
rect 8178 16348 8242 16352
rect 8178 16292 8182 16348
rect 8182 16292 8238 16348
rect 8238 16292 8242 16348
rect 8178 16288 8242 16292
rect 8258 16348 8322 16352
rect 8258 16292 8262 16348
rect 8262 16292 8318 16348
rect 8318 16292 8322 16348
rect 8258 16288 8322 16292
rect 8338 16348 8402 16352
rect 8338 16292 8342 16348
rect 8342 16292 8398 16348
rect 8398 16292 8402 16348
rect 8338 16288 8402 16292
rect 8418 16348 8482 16352
rect 8418 16292 8422 16348
rect 8422 16292 8478 16348
rect 8478 16292 8482 16348
rect 8418 16288 8482 16292
rect 3842 15804 3906 15808
rect 3842 15748 3846 15804
rect 3846 15748 3902 15804
rect 3902 15748 3906 15804
rect 3842 15744 3906 15748
rect 3922 15804 3986 15808
rect 3922 15748 3926 15804
rect 3926 15748 3982 15804
rect 3982 15748 3986 15804
rect 3922 15744 3986 15748
rect 4002 15804 4066 15808
rect 4002 15748 4006 15804
rect 4006 15748 4062 15804
rect 4062 15748 4066 15804
rect 4002 15744 4066 15748
rect 4082 15804 4146 15808
rect 4082 15748 4086 15804
rect 4086 15748 4142 15804
rect 4142 15748 4146 15804
rect 4082 15744 4146 15748
rect 6733 15804 6797 15808
rect 6733 15748 6737 15804
rect 6737 15748 6793 15804
rect 6793 15748 6797 15804
rect 6733 15744 6797 15748
rect 6813 15804 6877 15808
rect 6813 15748 6817 15804
rect 6817 15748 6873 15804
rect 6873 15748 6877 15804
rect 6813 15744 6877 15748
rect 6893 15804 6957 15808
rect 6893 15748 6897 15804
rect 6897 15748 6953 15804
rect 6953 15748 6957 15804
rect 6893 15744 6957 15748
rect 6973 15804 7037 15808
rect 6973 15748 6977 15804
rect 6977 15748 7033 15804
rect 7033 15748 7037 15804
rect 6973 15744 7037 15748
rect 2397 15260 2461 15264
rect 2397 15204 2401 15260
rect 2401 15204 2457 15260
rect 2457 15204 2461 15260
rect 2397 15200 2461 15204
rect 2477 15260 2541 15264
rect 2477 15204 2481 15260
rect 2481 15204 2537 15260
rect 2537 15204 2541 15260
rect 2477 15200 2541 15204
rect 2557 15260 2621 15264
rect 2557 15204 2561 15260
rect 2561 15204 2617 15260
rect 2617 15204 2621 15260
rect 2557 15200 2621 15204
rect 2637 15260 2701 15264
rect 2637 15204 2641 15260
rect 2641 15204 2697 15260
rect 2697 15204 2701 15260
rect 2637 15200 2701 15204
rect 5288 15260 5352 15264
rect 5288 15204 5292 15260
rect 5292 15204 5348 15260
rect 5348 15204 5352 15260
rect 5288 15200 5352 15204
rect 5368 15260 5432 15264
rect 5368 15204 5372 15260
rect 5372 15204 5428 15260
rect 5428 15204 5432 15260
rect 5368 15200 5432 15204
rect 5448 15260 5512 15264
rect 5448 15204 5452 15260
rect 5452 15204 5508 15260
rect 5508 15204 5512 15260
rect 5448 15200 5512 15204
rect 5528 15260 5592 15264
rect 5528 15204 5532 15260
rect 5532 15204 5588 15260
rect 5588 15204 5592 15260
rect 5528 15200 5592 15204
rect 8178 15260 8242 15264
rect 8178 15204 8182 15260
rect 8182 15204 8238 15260
rect 8238 15204 8242 15260
rect 8178 15200 8242 15204
rect 8258 15260 8322 15264
rect 8258 15204 8262 15260
rect 8262 15204 8318 15260
rect 8318 15204 8322 15260
rect 8258 15200 8322 15204
rect 8338 15260 8402 15264
rect 8338 15204 8342 15260
rect 8342 15204 8398 15260
rect 8398 15204 8402 15260
rect 8338 15200 8402 15204
rect 8418 15260 8482 15264
rect 8418 15204 8422 15260
rect 8422 15204 8478 15260
rect 8478 15204 8482 15260
rect 8418 15200 8482 15204
rect 3842 14716 3906 14720
rect 3842 14660 3846 14716
rect 3846 14660 3902 14716
rect 3902 14660 3906 14716
rect 3842 14656 3906 14660
rect 3922 14716 3986 14720
rect 3922 14660 3926 14716
rect 3926 14660 3982 14716
rect 3982 14660 3986 14716
rect 3922 14656 3986 14660
rect 4002 14716 4066 14720
rect 4002 14660 4006 14716
rect 4006 14660 4062 14716
rect 4062 14660 4066 14716
rect 4002 14656 4066 14660
rect 4082 14716 4146 14720
rect 4082 14660 4086 14716
rect 4086 14660 4142 14716
rect 4142 14660 4146 14716
rect 4082 14656 4146 14660
rect 6733 14716 6797 14720
rect 6733 14660 6737 14716
rect 6737 14660 6793 14716
rect 6793 14660 6797 14716
rect 6733 14656 6797 14660
rect 6813 14716 6877 14720
rect 6813 14660 6817 14716
rect 6817 14660 6873 14716
rect 6873 14660 6877 14716
rect 6813 14656 6877 14660
rect 6893 14716 6957 14720
rect 6893 14660 6897 14716
rect 6897 14660 6953 14716
rect 6953 14660 6957 14716
rect 6893 14656 6957 14660
rect 6973 14716 7037 14720
rect 6973 14660 6977 14716
rect 6977 14660 7033 14716
rect 7033 14660 7037 14716
rect 6973 14656 7037 14660
rect 2397 14172 2461 14176
rect 2397 14116 2401 14172
rect 2401 14116 2457 14172
rect 2457 14116 2461 14172
rect 2397 14112 2461 14116
rect 2477 14172 2541 14176
rect 2477 14116 2481 14172
rect 2481 14116 2537 14172
rect 2537 14116 2541 14172
rect 2477 14112 2541 14116
rect 2557 14172 2621 14176
rect 2557 14116 2561 14172
rect 2561 14116 2617 14172
rect 2617 14116 2621 14172
rect 2557 14112 2621 14116
rect 2637 14172 2701 14176
rect 2637 14116 2641 14172
rect 2641 14116 2697 14172
rect 2697 14116 2701 14172
rect 2637 14112 2701 14116
rect 5288 14172 5352 14176
rect 5288 14116 5292 14172
rect 5292 14116 5348 14172
rect 5348 14116 5352 14172
rect 5288 14112 5352 14116
rect 5368 14172 5432 14176
rect 5368 14116 5372 14172
rect 5372 14116 5428 14172
rect 5428 14116 5432 14172
rect 5368 14112 5432 14116
rect 5448 14172 5512 14176
rect 5448 14116 5452 14172
rect 5452 14116 5508 14172
rect 5508 14116 5512 14172
rect 5448 14112 5512 14116
rect 5528 14172 5592 14176
rect 5528 14116 5532 14172
rect 5532 14116 5588 14172
rect 5588 14116 5592 14172
rect 5528 14112 5592 14116
rect 8178 14172 8242 14176
rect 8178 14116 8182 14172
rect 8182 14116 8238 14172
rect 8238 14116 8242 14172
rect 8178 14112 8242 14116
rect 8258 14172 8322 14176
rect 8258 14116 8262 14172
rect 8262 14116 8318 14172
rect 8318 14116 8322 14172
rect 8258 14112 8322 14116
rect 8338 14172 8402 14176
rect 8338 14116 8342 14172
rect 8342 14116 8398 14172
rect 8398 14116 8402 14172
rect 8338 14112 8402 14116
rect 8418 14172 8482 14176
rect 8418 14116 8422 14172
rect 8422 14116 8478 14172
rect 8478 14116 8482 14172
rect 8418 14112 8482 14116
rect 3842 13628 3906 13632
rect 3842 13572 3846 13628
rect 3846 13572 3902 13628
rect 3902 13572 3906 13628
rect 3842 13568 3906 13572
rect 3922 13628 3986 13632
rect 3922 13572 3926 13628
rect 3926 13572 3982 13628
rect 3982 13572 3986 13628
rect 3922 13568 3986 13572
rect 4002 13628 4066 13632
rect 4002 13572 4006 13628
rect 4006 13572 4062 13628
rect 4062 13572 4066 13628
rect 4002 13568 4066 13572
rect 4082 13628 4146 13632
rect 4082 13572 4086 13628
rect 4086 13572 4142 13628
rect 4142 13572 4146 13628
rect 4082 13568 4146 13572
rect 6733 13628 6797 13632
rect 6733 13572 6737 13628
rect 6737 13572 6793 13628
rect 6793 13572 6797 13628
rect 6733 13568 6797 13572
rect 6813 13628 6877 13632
rect 6813 13572 6817 13628
rect 6817 13572 6873 13628
rect 6873 13572 6877 13628
rect 6813 13568 6877 13572
rect 6893 13628 6957 13632
rect 6893 13572 6897 13628
rect 6897 13572 6953 13628
rect 6953 13572 6957 13628
rect 6893 13568 6957 13572
rect 6973 13628 7037 13632
rect 6973 13572 6977 13628
rect 6977 13572 7033 13628
rect 7033 13572 7037 13628
rect 6973 13568 7037 13572
rect 2397 13084 2461 13088
rect 2397 13028 2401 13084
rect 2401 13028 2457 13084
rect 2457 13028 2461 13084
rect 2397 13024 2461 13028
rect 2477 13084 2541 13088
rect 2477 13028 2481 13084
rect 2481 13028 2537 13084
rect 2537 13028 2541 13084
rect 2477 13024 2541 13028
rect 2557 13084 2621 13088
rect 2557 13028 2561 13084
rect 2561 13028 2617 13084
rect 2617 13028 2621 13084
rect 2557 13024 2621 13028
rect 2637 13084 2701 13088
rect 2637 13028 2641 13084
rect 2641 13028 2697 13084
rect 2697 13028 2701 13084
rect 2637 13024 2701 13028
rect 5288 13084 5352 13088
rect 5288 13028 5292 13084
rect 5292 13028 5348 13084
rect 5348 13028 5352 13084
rect 5288 13024 5352 13028
rect 5368 13084 5432 13088
rect 5368 13028 5372 13084
rect 5372 13028 5428 13084
rect 5428 13028 5432 13084
rect 5368 13024 5432 13028
rect 5448 13084 5512 13088
rect 5448 13028 5452 13084
rect 5452 13028 5508 13084
rect 5508 13028 5512 13084
rect 5448 13024 5512 13028
rect 5528 13084 5592 13088
rect 5528 13028 5532 13084
rect 5532 13028 5588 13084
rect 5588 13028 5592 13084
rect 5528 13024 5592 13028
rect 8178 13084 8242 13088
rect 8178 13028 8182 13084
rect 8182 13028 8238 13084
rect 8238 13028 8242 13084
rect 8178 13024 8242 13028
rect 8258 13084 8322 13088
rect 8258 13028 8262 13084
rect 8262 13028 8318 13084
rect 8318 13028 8322 13084
rect 8258 13024 8322 13028
rect 8338 13084 8402 13088
rect 8338 13028 8342 13084
rect 8342 13028 8398 13084
rect 8398 13028 8402 13084
rect 8338 13024 8402 13028
rect 8418 13084 8482 13088
rect 8418 13028 8422 13084
rect 8422 13028 8478 13084
rect 8478 13028 8482 13084
rect 8418 13024 8482 13028
rect 3842 12540 3906 12544
rect 3842 12484 3846 12540
rect 3846 12484 3902 12540
rect 3902 12484 3906 12540
rect 3842 12480 3906 12484
rect 3922 12540 3986 12544
rect 3922 12484 3926 12540
rect 3926 12484 3982 12540
rect 3982 12484 3986 12540
rect 3922 12480 3986 12484
rect 4002 12540 4066 12544
rect 4002 12484 4006 12540
rect 4006 12484 4062 12540
rect 4062 12484 4066 12540
rect 4002 12480 4066 12484
rect 4082 12540 4146 12544
rect 4082 12484 4086 12540
rect 4086 12484 4142 12540
rect 4142 12484 4146 12540
rect 4082 12480 4146 12484
rect 6733 12540 6797 12544
rect 6733 12484 6737 12540
rect 6737 12484 6793 12540
rect 6793 12484 6797 12540
rect 6733 12480 6797 12484
rect 6813 12540 6877 12544
rect 6813 12484 6817 12540
rect 6817 12484 6873 12540
rect 6873 12484 6877 12540
rect 6813 12480 6877 12484
rect 6893 12540 6957 12544
rect 6893 12484 6897 12540
rect 6897 12484 6953 12540
rect 6953 12484 6957 12540
rect 6893 12480 6957 12484
rect 6973 12540 7037 12544
rect 6973 12484 6977 12540
rect 6977 12484 7033 12540
rect 7033 12484 7037 12540
rect 6973 12480 7037 12484
rect 2397 11996 2461 12000
rect 2397 11940 2401 11996
rect 2401 11940 2457 11996
rect 2457 11940 2461 11996
rect 2397 11936 2461 11940
rect 2477 11996 2541 12000
rect 2477 11940 2481 11996
rect 2481 11940 2537 11996
rect 2537 11940 2541 11996
rect 2477 11936 2541 11940
rect 2557 11996 2621 12000
rect 2557 11940 2561 11996
rect 2561 11940 2617 11996
rect 2617 11940 2621 11996
rect 2557 11936 2621 11940
rect 2637 11996 2701 12000
rect 2637 11940 2641 11996
rect 2641 11940 2697 11996
rect 2697 11940 2701 11996
rect 2637 11936 2701 11940
rect 5288 11996 5352 12000
rect 5288 11940 5292 11996
rect 5292 11940 5348 11996
rect 5348 11940 5352 11996
rect 5288 11936 5352 11940
rect 5368 11996 5432 12000
rect 5368 11940 5372 11996
rect 5372 11940 5428 11996
rect 5428 11940 5432 11996
rect 5368 11936 5432 11940
rect 5448 11996 5512 12000
rect 5448 11940 5452 11996
rect 5452 11940 5508 11996
rect 5508 11940 5512 11996
rect 5448 11936 5512 11940
rect 5528 11996 5592 12000
rect 5528 11940 5532 11996
rect 5532 11940 5588 11996
rect 5588 11940 5592 11996
rect 5528 11936 5592 11940
rect 8178 11996 8242 12000
rect 8178 11940 8182 11996
rect 8182 11940 8238 11996
rect 8238 11940 8242 11996
rect 8178 11936 8242 11940
rect 8258 11996 8322 12000
rect 8258 11940 8262 11996
rect 8262 11940 8318 11996
rect 8318 11940 8322 11996
rect 8258 11936 8322 11940
rect 8338 11996 8402 12000
rect 8338 11940 8342 11996
rect 8342 11940 8398 11996
rect 8398 11940 8402 11996
rect 8338 11936 8402 11940
rect 8418 11996 8482 12000
rect 8418 11940 8422 11996
rect 8422 11940 8478 11996
rect 8478 11940 8482 11996
rect 8418 11936 8482 11940
rect 3842 11452 3906 11456
rect 3842 11396 3846 11452
rect 3846 11396 3902 11452
rect 3902 11396 3906 11452
rect 3842 11392 3906 11396
rect 3922 11452 3986 11456
rect 3922 11396 3926 11452
rect 3926 11396 3982 11452
rect 3982 11396 3986 11452
rect 3922 11392 3986 11396
rect 4002 11452 4066 11456
rect 4002 11396 4006 11452
rect 4006 11396 4062 11452
rect 4062 11396 4066 11452
rect 4002 11392 4066 11396
rect 4082 11452 4146 11456
rect 4082 11396 4086 11452
rect 4086 11396 4142 11452
rect 4142 11396 4146 11452
rect 4082 11392 4146 11396
rect 6733 11452 6797 11456
rect 6733 11396 6737 11452
rect 6737 11396 6793 11452
rect 6793 11396 6797 11452
rect 6733 11392 6797 11396
rect 6813 11452 6877 11456
rect 6813 11396 6817 11452
rect 6817 11396 6873 11452
rect 6873 11396 6877 11452
rect 6813 11392 6877 11396
rect 6893 11452 6957 11456
rect 6893 11396 6897 11452
rect 6897 11396 6953 11452
rect 6953 11396 6957 11452
rect 6893 11392 6957 11396
rect 6973 11452 7037 11456
rect 6973 11396 6977 11452
rect 6977 11396 7033 11452
rect 7033 11396 7037 11452
rect 6973 11392 7037 11396
rect 2397 10908 2461 10912
rect 2397 10852 2401 10908
rect 2401 10852 2457 10908
rect 2457 10852 2461 10908
rect 2397 10848 2461 10852
rect 2477 10908 2541 10912
rect 2477 10852 2481 10908
rect 2481 10852 2537 10908
rect 2537 10852 2541 10908
rect 2477 10848 2541 10852
rect 2557 10908 2621 10912
rect 2557 10852 2561 10908
rect 2561 10852 2617 10908
rect 2617 10852 2621 10908
rect 2557 10848 2621 10852
rect 2637 10908 2701 10912
rect 2637 10852 2641 10908
rect 2641 10852 2697 10908
rect 2697 10852 2701 10908
rect 2637 10848 2701 10852
rect 5288 10908 5352 10912
rect 5288 10852 5292 10908
rect 5292 10852 5348 10908
rect 5348 10852 5352 10908
rect 5288 10848 5352 10852
rect 5368 10908 5432 10912
rect 5368 10852 5372 10908
rect 5372 10852 5428 10908
rect 5428 10852 5432 10908
rect 5368 10848 5432 10852
rect 5448 10908 5512 10912
rect 5448 10852 5452 10908
rect 5452 10852 5508 10908
rect 5508 10852 5512 10908
rect 5448 10848 5512 10852
rect 5528 10908 5592 10912
rect 5528 10852 5532 10908
rect 5532 10852 5588 10908
rect 5588 10852 5592 10908
rect 5528 10848 5592 10852
rect 8178 10908 8242 10912
rect 8178 10852 8182 10908
rect 8182 10852 8238 10908
rect 8238 10852 8242 10908
rect 8178 10848 8242 10852
rect 8258 10908 8322 10912
rect 8258 10852 8262 10908
rect 8262 10852 8318 10908
rect 8318 10852 8322 10908
rect 8258 10848 8322 10852
rect 8338 10908 8402 10912
rect 8338 10852 8342 10908
rect 8342 10852 8398 10908
rect 8398 10852 8402 10908
rect 8338 10848 8402 10852
rect 8418 10908 8482 10912
rect 8418 10852 8422 10908
rect 8422 10852 8478 10908
rect 8478 10852 8482 10908
rect 8418 10848 8482 10852
rect 3842 10364 3906 10368
rect 3842 10308 3846 10364
rect 3846 10308 3902 10364
rect 3902 10308 3906 10364
rect 3842 10304 3906 10308
rect 3922 10364 3986 10368
rect 3922 10308 3926 10364
rect 3926 10308 3982 10364
rect 3982 10308 3986 10364
rect 3922 10304 3986 10308
rect 4002 10364 4066 10368
rect 4002 10308 4006 10364
rect 4006 10308 4062 10364
rect 4062 10308 4066 10364
rect 4002 10304 4066 10308
rect 4082 10364 4146 10368
rect 4082 10308 4086 10364
rect 4086 10308 4142 10364
rect 4142 10308 4146 10364
rect 4082 10304 4146 10308
rect 6733 10364 6797 10368
rect 6733 10308 6737 10364
rect 6737 10308 6793 10364
rect 6793 10308 6797 10364
rect 6733 10304 6797 10308
rect 6813 10364 6877 10368
rect 6813 10308 6817 10364
rect 6817 10308 6873 10364
rect 6873 10308 6877 10364
rect 6813 10304 6877 10308
rect 6893 10364 6957 10368
rect 6893 10308 6897 10364
rect 6897 10308 6953 10364
rect 6953 10308 6957 10364
rect 6893 10304 6957 10308
rect 6973 10364 7037 10368
rect 6973 10308 6977 10364
rect 6977 10308 7033 10364
rect 7033 10308 7037 10364
rect 6973 10304 7037 10308
rect 2397 9820 2461 9824
rect 2397 9764 2401 9820
rect 2401 9764 2457 9820
rect 2457 9764 2461 9820
rect 2397 9760 2461 9764
rect 2477 9820 2541 9824
rect 2477 9764 2481 9820
rect 2481 9764 2537 9820
rect 2537 9764 2541 9820
rect 2477 9760 2541 9764
rect 2557 9820 2621 9824
rect 2557 9764 2561 9820
rect 2561 9764 2617 9820
rect 2617 9764 2621 9820
rect 2557 9760 2621 9764
rect 2637 9820 2701 9824
rect 2637 9764 2641 9820
rect 2641 9764 2697 9820
rect 2697 9764 2701 9820
rect 2637 9760 2701 9764
rect 5288 9820 5352 9824
rect 5288 9764 5292 9820
rect 5292 9764 5348 9820
rect 5348 9764 5352 9820
rect 5288 9760 5352 9764
rect 5368 9820 5432 9824
rect 5368 9764 5372 9820
rect 5372 9764 5428 9820
rect 5428 9764 5432 9820
rect 5368 9760 5432 9764
rect 5448 9820 5512 9824
rect 5448 9764 5452 9820
rect 5452 9764 5508 9820
rect 5508 9764 5512 9820
rect 5448 9760 5512 9764
rect 5528 9820 5592 9824
rect 5528 9764 5532 9820
rect 5532 9764 5588 9820
rect 5588 9764 5592 9820
rect 5528 9760 5592 9764
rect 8178 9820 8242 9824
rect 8178 9764 8182 9820
rect 8182 9764 8238 9820
rect 8238 9764 8242 9820
rect 8178 9760 8242 9764
rect 8258 9820 8322 9824
rect 8258 9764 8262 9820
rect 8262 9764 8318 9820
rect 8318 9764 8322 9820
rect 8258 9760 8322 9764
rect 8338 9820 8402 9824
rect 8338 9764 8342 9820
rect 8342 9764 8398 9820
rect 8398 9764 8402 9820
rect 8338 9760 8402 9764
rect 8418 9820 8482 9824
rect 8418 9764 8422 9820
rect 8422 9764 8478 9820
rect 8478 9764 8482 9820
rect 8418 9760 8482 9764
rect 3842 9276 3906 9280
rect 3842 9220 3846 9276
rect 3846 9220 3902 9276
rect 3902 9220 3906 9276
rect 3842 9216 3906 9220
rect 3922 9276 3986 9280
rect 3922 9220 3926 9276
rect 3926 9220 3982 9276
rect 3982 9220 3986 9276
rect 3922 9216 3986 9220
rect 4002 9276 4066 9280
rect 4002 9220 4006 9276
rect 4006 9220 4062 9276
rect 4062 9220 4066 9276
rect 4002 9216 4066 9220
rect 4082 9276 4146 9280
rect 4082 9220 4086 9276
rect 4086 9220 4142 9276
rect 4142 9220 4146 9276
rect 4082 9216 4146 9220
rect 6733 9276 6797 9280
rect 6733 9220 6737 9276
rect 6737 9220 6793 9276
rect 6793 9220 6797 9276
rect 6733 9216 6797 9220
rect 6813 9276 6877 9280
rect 6813 9220 6817 9276
rect 6817 9220 6873 9276
rect 6873 9220 6877 9276
rect 6813 9216 6877 9220
rect 6893 9276 6957 9280
rect 6893 9220 6897 9276
rect 6897 9220 6953 9276
rect 6953 9220 6957 9276
rect 6893 9216 6957 9220
rect 6973 9276 7037 9280
rect 6973 9220 6977 9276
rect 6977 9220 7033 9276
rect 7033 9220 7037 9276
rect 6973 9216 7037 9220
rect 2397 8732 2461 8736
rect 2397 8676 2401 8732
rect 2401 8676 2457 8732
rect 2457 8676 2461 8732
rect 2397 8672 2461 8676
rect 2477 8732 2541 8736
rect 2477 8676 2481 8732
rect 2481 8676 2537 8732
rect 2537 8676 2541 8732
rect 2477 8672 2541 8676
rect 2557 8732 2621 8736
rect 2557 8676 2561 8732
rect 2561 8676 2617 8732
rect 2617 8676 2621 8732
rect 2557 8672 2621 8676
rect 2637 8732 2701 8736
rect 2637 8676 2641 8732
rect 2641 8676 2697 8732
rect 2697 8676 2701 8732
rect 2637 8672 2701 8676
rect 5288 8732 5352 8736
rect 5288 8676 5292 8732
rect 5292 8676 5348 8732
rect 5348 8676 5352 8732
rect 5288 8672 5352 8676
rect 5368 8732 5432 8736
rect 5368 8676 5372 8732
rect 5372 8676 5428 8732
rect 5428 8676 5432 8732
rect 5368 8672 5432 8676
rect 5448 8732 5512 8736
rect 5448 8676 5452 8732
rect 5452 8676 5508 8732
rect 5508 8676 5512 8732
rect 5448 8672 5512 8676
rect 5528 8732 5592 8736
rect 5528 8676 5532 8732
rect 5532 8676 5588 8732
rect 5588 8676 5592 8732
rect 5528 8672 5592 8676
rect 8178 8732 8242 8736
rect 8178 8676 8182 8732
rect 8182 8676 8238 8732
rect 8238 8676 8242 8732
rect 8178 8672 8242 8676
rect 8258 8732 8322 8736
rect 8258 8676 8262 8732
rect 8262 8676 8318 8732
rect 8318 8676 8322 8732
rect 8258 8672 8322 8676
rect 8338 8732 8402 8736
rect 8338 8676 8342 8732
rect 8342 8676 8398 8732
rect 8398 8676 8402 8732
rect 8338 8672 8402 8676
rect 8418 8732 8482 8736
rect 8418 8676 8422 8732
rect 8422 8676 8478 8732
rect 8478 8676 8482 8732
rect 8418 8672 8482 8676
rect 3842 8188 3906 8192
rect 3842 8132 3846 8188
rect 3846 8132 3902 8188
rect 3902 8132 3906 8188
rect 3842 8128 3906 8132
rect 3922 8188 3986 8192
rect 3922 8132 3926 8188
rect 3926 8132 3982 8188
rect 3982 8132 3986 8188
rect 3922 8128 3986 8132
rect 4002 8188 4066 8192
rect 4002 8132 4006 8188
rect 4006 8132 4062 8188
rect 4062 8132 4066 8188
rect 4002 8128 4066 8132
rect 4082 8188 4146 8192
rect 4082 8132 4086 8188
rect 4086 8132 4142 8188
rect 4142 8132 4146 8188
rect 4082 8128 4146 8132
rect 6733 8188 6797 8192
rect 6733 8132 6737 8188
rect 6737 8132 6793 8188
rect 6793 8132 6797 8188
rect 6733 8128 6797 8132
rect 6813 8188 6877 8192
rect 6813 8132 6817 8188
rect 6817 8132 6873 8188
rect 6873 8132 6877 8188
rect 6813 8128 6877 8132
rect 6893 8188 6957 8192
rect 6893 8132 6897 8188
rect 6897 8132 6953 8188
rect 6953 8132 6957 8188
rect 6893 8128 6957 8132
rect 6973 8188 7037 8192
rect 6973 8132 6977 8188
rect 6977 8132 7033 8188
rect 7033 8132 7037 8188
rect 6973 8128 7037 8132
rect 2397 7644 2461 7648
rect 2397 7588 2401 7644
rect 2401 7588 2457 7644
rect 2457 7588 2461 7644
rect 2397 7584 2461 7588
rect 2477 7644 2541 7648
rect 2477 7588 2481 7644
rect 2481 7588 2537 7644
rect 2537 7588 2541 7644
rect 2477 7584 2541 7588
rect 2557 7644 2621 7648
rect 2557 7588 2561 7644
rect 2561 7588 2617 7644
rect 2617 7588 2621 7644
rect 2557 7584 2621 7588
rect 2637 7644 2701 7648
rect 2637 7588 2641 7644
rect 2641 7588 2697 7644
rect 2697 7588 2701 7644
rect 2637 7584 2701 7588
rect 5288 7644 5352 7648
rect 5288 7588 5292 7644
rect 5292 7588 5348 7644
rect 5348 7588 5352 7644
rect 5288 7584 5352 7588
rect 5368 7644 5432 7648
rect 5368 7588 5372 7644
rect 5372 7588 5428 7644
rect 5428 7588 5432 7644
rect 5368 7584 5432 7588
rect 5448 7644 5512 7648
rect 5448 7588 5452 7644
rect 5452 7588 5508 7644
rect 5508 7588 5512 7644
rect 5448 7584 5512 7588
rect 5528 7644 5592 7648
rect 5528 7588 5532 7644
rect 5532 7588 5588 7644
rect 5588 7588 5592 7644
rect 5528 7584 5592 7588
rect 8178 7644 8242 7648
rect 8178 7588 8182 7644
rect 8182 7588 8238 7644
rect 8238 7588 8242 7644
rect 8178 7584 8242 7588
rect 8258 7644 8322 7648
rect 8258 7588 8262 7644
rect 8262 7588 8318 7644
rect 8318 7588 8322 7644
rect 8258 7584 8322 7588
rect 8338 7644 8402 7648
rect 8338 7588 8342 7644
rect 8342 7588 8398 7644
rect 8398 7588 8402 7644
rect 8338 7584 8402 7588
rect 8418 7644 8482 7648
rect 8418 7588 8422 7644
rect 8422 7588 8478 7644
rect 8478 7588 8482 7644
rect 8418 7584 8482 7588
rect 3842 7100 3906 7104
rect 3842 7044 3846 7100
rect 3846 7044 3902 7100
rect 3902 7044 3906 7100
rect 3842 7040 3906 7044
rect 3922 7100 3986 7104
rect 3922 7044 3926 7100
rect 3926 7044 3982 7100
rect 3982 7044 3986 7100
rect 3922 7040 3986 7044
rect 4002 7100 4066 7104
rect 4002 7044 4006 7100
rect 4006 7044 4062 7100
rect 4062 7044 4066 7100
rect 4002 7040 4066 7044
rect 4082 7100 4146 7104
rect 4082 7044 4086 7100
rect 4086 7044 4142 7100
rect 4142 7044 4146 7100
rect 4082 7040 4146 7044
rect 6733 7100 6797 7104
rect 6733 7044 6737 7100
rect 6737 7044 6793 7100
rect 6793 7044 6797 7100
rect 6733 7040 6797 7044
rect 6813 7100 6877 7104
rect 6813 7044 6817 7100
rect 6817 7044 6873 7100
rect 6873 7044 6877 7100
rect 6813 7040 6877 7044
rect 6893 7100 6957 7104
rect 6893 7044 6897 7100
rect 6897 7044 6953 7100
rect 6953 7044 6957 7100
rect 6893 7040 6957 7044
rect 6973 7100 7037 7104
rect 6973 7044 6977 7100
rect 6977 7044 7033 7100
rect 7033 7044 7037 7100
rect 6973 7040 7037 7044
rect 2397 6556 2461 6560
rect 2397 6500 2401 6556
rect 2401 6500 2457 6556
rect 2457 6500 2461 6556
rect 2397 6496 2461 6500
rect 2477 6556 2541 6560
rect 2477 6500 2481 6556
rect 2481 6500 2537 6556
rect 2537 6500 2541 6556
rect 2477 6496 2541 6500
rect 2557 6556 2621 6560
rect 2557 6500 2561 6556
rect 2561 6500 2617 6556
rect 2617 6500 2621 6556
rect 2557 6496 2621 6500
rect 2637 6556 2701 6560
rect 2637 6500 2641 6556
rect 2641 6500 2697 6556
rect 2697 6500 2701 6556
rect 2637 6496 2701 6500
rect 5288 6556 5352 6560
rect 5288 6500 5292 6556
rect 5292 6500 5348 6556
rect 5348 6500 5352 6556
rect 5288 6496 5352 6500
rect 5368 6556 5432 6560
rect 5368 6500 5372 6556
rect 5372 6500 5428 6556
rect 5428 6500 5432 6556
rect 5368 6496 5432 6500
rect 5448 6556 5512 6560
rect 5448 6500 5452 6556
rect 5452 6500 5508 6556
rect 5508 6500 5512 6556
rect 5448 6496 5512 6500
rect 5528 6556 5592 6560
rect 5528 6500 5532 6556
rect 5532 6500 5588 6556
rect 5588 6500 5592 6556
rect 5528 6496 5592 6500
rect 8178 6556 8242 6560
rect 8178 6500 8182 6556
rect 8182 6500 8238 6556
rect 8238 6500 8242 6556
rect 8178 6496 8242 6500
rect 8258 6556 8322 6560
rect 8258 6500 8262 6556
rect 8262 6500 8318 6556
rect 8318 6500 8322 6556
rect 8258 6496 8322 6500
rect 8338 6556 8402 6560
rect 8338 6500 8342 6556
rect 8342 6500 8398 6556
rect 8398 6500 8402 6556
rect 8338 6496 8402 6500
rect 8418 6556 8482 6560
rect 8418 6500 8422 6556
rect 8422 6500 8478 6556
rect 8478 6500 8482 6556
rect 8418 6496 8482 6500
rect 3842 6012 3906 6016
rect 3842 5956 3846 6012
rect 3846 5956 3902 6012
rect 3902 5956 3906 6012
rect 3842 5952 3906 5956
rect 3922 6012 3986 6016
rect 3922 5956 3926 6012
rect 3926 5956 3982 6012
rect 3982 5956 3986 6012
rect 3922 5952 3986 5956
rect 4002 6012 4066 6016
rect 4002 5956 4006 6012
rect 4006 5956 4062 6012
rect 4062 5956 4066 6012
rect 4002 5952 4066 5956
rect 4082 6012 4146 6016
rect 4082 5956 4086 6012
rect 4086 5956 4142 6012
rect 4142 5956 4146 6012
rect 4082 5952 4146 5956
rect 6733 6012 6797 6016
rect 6733 5956 6737 6012
rect 6737 5956 6793 6012
rect 6793 5956 6797 6012
rect 6733 5952 6797 5956
rect 6813 6012 6877 6016
rect 6813 5956 6817 6012
rect 6817 5956 6873 6012
rect 6873 5956 6877 6012
rect 6813 5952 6877 5956
rect 6893 6012 6957 6016
rect 6893 5956 6897 6012
rect 6897 5956 6953 6012
rect 6953 5956 6957 6012
rect 6893 5952 6957 5956
rect 6973 6012 7037 6016
rect 6973 5956 6977 6012
rect 6977 5956 7033 6012
rect 7033 5956 7037 6012
rect 6973 5952 7037 5956
rect 2397 5468 2461 5472
rect 2397 5412 2401 5468
rect 2401 5412 2457 5468
rect 2457 5412 2461 5468
rect 2397 5408 2461 5412
rect 2477 5468 2541 5472
rect 2477 5412 2481 5468
rect 2481 5412 2537 5468
rect 2537 5412 2541 5468
rect 2477 5408 2541 5412
rect 2557 5468 2621 5472
rect 2557 5412 2561 5468
rect 2561 5412 2617 5468
rect 2617 5412 2621 5468
rect 2557 5408 2621 5412
rect 2637 5468 2701 5472
rect 2637 5412 2641 5468
rect 2641 5412 2697 5468
rect 2697 5412 2701 5468
rect 2637 5408 2701 5412
rect 5288 5468 5352 5472
rect 5288 5412 5292 5468
rect 5292 5412 5348 5468
rect 5348 5412 5352 5468
rect 5288 5408 5352 5412
rect 5368 5468 5432 5472
rect 5368 5412 5372 5468
rect 5372 5412 5428 5468
rect 5428 5412 5432 5468
rect 5368 5408 5432 5412
rect 5448 5468 5512 5472
rect 5448 5412 5452 5468
rect 5452 5412 5508 5468
rect 5508 5412 5512 5468
rect 5448 5408 5512 5412
rect 5528 5468 5592 5472
rect 5528 5412 5532 5468
rect 5532 5412 5588 5468
rect 5588 5412 5592 5468
rect 5528 5408 5592 5412
rect 8178 5468 8242 5472
rect 8178 5412 8182 5468
rect 8182 5412 8238 5468
rect 8238 5412 8242 5468
rect 8178 5408 8242 5412
rect 8258 5468 8322 5472
rect 8258 5412 8262 5468
rect 8262 5412 8318 5468
rect 8318 5412 8322 5468
rect 8258 5408 8322 5412
rect 8338 5468 8402 5472
rect 8338 5412 8342 5468
rect 8342 5412 8398 5468
rect 8398 5412 8402 5468
rect 8338 5408 8402 5412
rect 8418 5468 8482 5472
rect 8418 5412 8422 5468
rect 8422 5412 8478 5468
rect 8478 5412 8482 5468
rect 8418 5408 8482 5412
rect 3842 4924 3906 4928
rect 3842 4868 3846 4924
rect 3846 4868 3902 4924
rect 3902 4868 3906 4924
rect 3842 4864 3906 4868
rect 3922 4924 3986 4928
rect 3922 4868 3926 4924
rect 3926 4868 3982 4924
rect 3982 4868 3986 4924
rect 3922 4864 3986 4868
rect 4002 4924 4066 4928
rect 4002 4868 4006 4924
rect 4006 4868 4062 4924
rect 4062 4868 4066 4924
rect 4002 4864 4066 4868
rect 4082 4924 4146 4928
rect 4082 4868 4086 4924
rect 4086 4868 4142 4924
rect 4142 4868 4146 4924
rect 4082 4864 4146 4868
rect 6733 4924 6797 4928
rect 6733 4868 6737 4924
rect 6737 4868 6793 4924
rect 6793 4868 6797 4924
rect 6733 4864 6797 4868
rect 6813 4924 6877 4928
rect 6813 4868 6817 4924
rect 6817 4868 6873 4924
rect 6873 4868 6877 4924
rect 6813 4864 6877 4868
rect 6893 4924 6957 4928
rect 6893 4868 6897 4924
rect 6897 4868 6953 4924
rect 6953 4868 6957 4924
rect 6893 4864 6957 4868
rect 6973 4924 7037 4928
rect 6973 4868 6977 4924
rect 6977 4868 7033 4924
rect 7033 4868 7037 4924
rect 6973 4864 7037 4868
rect 2397 4380 2461 4384
rect 2397 4324 2401 4380
rect 2401 4324 2457 4380
rect 2457 4324 2461 4380
rect 2397 4320 2461 4324
rect 2477 4380 2541 4384
rect 2477 4324 2481 4380
rect 2481 4324 2537 4380
rect 2537 4324 2541 4380
rect 2477 4320 2541 4324
rect 2557 4380 2621 4384
rect 2557 4324 2561 4380
rect 2561 4324 2617 4380
rect 2617 4324 2621 4380
rect 2557 4320 2621 4324
rect 2637 4380 2701 4384
rect 2637 4324 2641 4380
rect 2641 4324 2697 4380
rect 2697 4324 2701 4380
rect 2637 4320 2701 4324
rect 5288 4380 5352 4384
rect 5288 4324 5292 4380
rect 5292 4324 5348 4380
rect 5348 4324 5352 4380
rect 5288 4320 5352 4324
rect 5368 4380 5432 4384
rect 5368 4324 5372 4380
rect 5372 4324 5428 4380
rect 5428 4324 5432 4380
rect 5368 4320 5432 4324
rect 5448 4380 5512 4384
rect 5448 4324 5452 4380
rect 5452 4324 5508 4380
rect 5508 4324 5512 4380
rect 5448 4320 5512 4324
rect 5528 4380 5592 4384
rect 5528 4324 5532 4380
rect 5532 4324 5588 4380
rect 5588 4324 5592 4380
rect 5528 4320 5592 4324
rect 8178 4380 8242 4384
rect 8178 4324 8182 4380
rect 8182 4324 8238 4380
rect 8238 4324 8242 4380
rect 8178 4320 8242 4324
rect 8258 4380 8322 4384
rect 8258 4324 8262 4380
rect 8262 4324 8318 4380
rect 8318 4324 8322 4380
rect 8258 4320 8322 4324
rect 8338 4380 8402 4384
rect 8338 4324 8342 4380
rect 8342 4324 8398 4380
rect 8398 4324 8402 4380
rect 8338 4320 8402 4324
rect 8418 4380 8482 4384
rect 8418 4324 8422 4380
rect 8422 4324 8478 4380
rect 8478 4324 8482 4380
rect 8418 4320 8482 4324
rect 3842 3836 3906 3840
rect 3842 3780 3846 3836
rect 3846 3780 3902 3836
rect 3902 3780 3906 3836
rect 3842 3776 3906 3780
rect 3922 3836 3986 3840
rect 3922 3780 3926 3836
rect 3926 3780 3982 3836
rect 3982 3780 3986 3836
rect 3922 3776 3986 3780
rect 4002 3836 4066 3840
rect 4002 3780 4006 3836
rect 4006 3780 4062 3836
rect 4062 3780 4066 3836
rect 4002 3776 4066 3780
rect 4082 3836 4146 3840
rect 4082 3780 4086 3836
rect 4086 3780 4142 3836
rect 4142 3780 4146 3836
rect 4082 3776 4146 3780
rect 6733 3836 6797 3840
rect 6733 3780 6737 3836
rect 6737 3780 6793 3836
rect 6793 3780 6797 3836
rect 6733 3776 6797 3780
rect 6813 3836 6877 3840
rect 6813 3780 6817 3836
rect 6817 3780 6873 3836
rect 6873 3780 6877 3836
rect 6813 3776 6877 3780
rect 6893 3836 6957 3840
rect 6893 3780 6897 3836
rect 6897 3780 6953 3836
rect 6953 3780 6957 3836
rect 6893 3776 6957 3780
rect 6973 3836 7037 3840
rect 6973 3780 6977 3836
rect 6977 3780 7033 3836
rect 7033 3780 7037 3836
rect 6973 3776 7037 3780
rect 2397 3292 2461 3296
rect 2397 3236 2401 3292
rect 2401 3236 2457 3292
rect 2457 3236 2461 3292
rect 2397 3232 2461 3236
rect 2477 3292 2541 3296
rect 2477 3236 2481 3292
rect 2481 3236 2537 3292
rect 2537 3236 2541 3292
rect 2477 3232 2541 3236
rect 2557 3292 2621 3296
rect 2557 3236 2561 3292
rect 2561 3236 2617 3292
rect 2617 3236 2621 3292
rect 2557 3232 2621 3236
rect 2637 3292 2701 3296
rect 2637 3236 2641 3292
rect 2641 3236 2697 3292
rect 2697 3236 2701 3292
rect 2637 3232 2701 3236
rect 5288 3292 5352 3296
rect 5288 3236 5292 3292
rect 5292 3236 5348 3292
rect 5348 3236 5352 3292
rect 5288 3232 5352 3236
rect 5368 3292 5432 3296
rect 5368 3236 5372 3292
rect 5372 3236 5428 3292
rect 5428 3236 5432 3292
rect 5368 3232 5432 3236
rect 5448 3292 5512 3296
rect 5448 3236 5452 3292
rect 5452 3236 5508 3292
rect 5508 3236 5512 3292
rect 5448 3232 5512 3236
rect 5528 3292 5592 3296
rect 5528 3236 5532 3292
rect 5532 3236 5588 3292
rect 5588 3236 5592 3292
rect 5528 3232 5592 3236
rect 8178 3292 8242 3296
rect 8178 3236 8182 3292
rect 8182 3236 8238 3292
rect 8238 3236 8242 3292
rect 8178 3232 8242 3236
rect 8258 3292 8322 3296
rect 8258 3236 8262 3292
rect 8262 3236 8318 3292
rect 8318 3236 8322 3292
rect 8258 3232 8322 3236
rect 8338 3292 8402 3296
rect 8338 3236 8342 3292
rect 8342 3236 8398 3292
rect 8398 3236 8402 3292
rect 8338 3232 8402 3236
rect 8418 3292 8482 3296
rect 8418 3236 8422 3292
rect 8422 3236 8478 3292
rect 8478 3236 8482 3292
rect 8418 3232 8482 3236
rect 3842 2748 3906 2752
rect 3842 2692 3846 2748
rect 3846 2692 3902 2748
rect 3902 2692 3906 2748
rect 3842 2688 3906 2692
rect 3922 2748 3986 2752
rect 3922 2692 3926 2748
rect 3926 2692 3982 2748
rect 3982 2692 3986 2748
rect 3922 2688 3986 2692
rect 4002 2748 4066 2752
rect 4002 2692 4006 2748
rect 4006 2692 4062 2748
rect 4062 2692 4066 2748
rect 4002 2688 4066 2692
rect 4082 2748 4146 2752
rect 4082 2692 4086 2748
rect 4086 2692 4142 2748
rect 4142 2692 4146 2748
rect 4082 2688 4146 2692
rect 6733 2748 6797 2752
rect 6733 2692 6737 2748
rect 6737 2692 6793 2748
rect 6793 2692 6797 2748
rect 6733 2688 6797 2692
rect 6813 2748 6877 2752
rect 6813 2692 6817 2748
rect 6817 2692 6873 2748
rect 6873 2692 6877 2748
rect 6813 2688 6877 2692
rect 6893 2748 6957 2752
rect 6893 2692 6897 2748
rect 6897 2692 6953 2748
rect 6953 2692 6957 2748
rect 6893 2688 6957 2692
rect 6973 2748 7037 2752
rect 6973 2692 6977 2748
rect 6977 2692 7033 2748
rect 7033 2692 7037 2748
rect 6973 2688 7037 2692
rect 2397 2204 2461 2208
rect 2397 2148 2401 2204
rect 2401 2148 2457 2204
rect 2457 2148 2461 2204
rect 2397 2144 2461 2148
rect 2477 2204 2541 2208
rect 2477 2148 2481 2204
rect 2481 2148 2537 2204
rect 2537 2148 2541 2204
rect 2477 2144 2541 2148
rect 2557 2204 2621 2208
rect 2557 2148 2561 2204
rect 2561 2148 2617 2204
rect 2617 2148 2621 2204
rect 2557 2144 2621 2148
rect 2637 2204 2701 2208
rect 2637 2148 2641 2204
rect 2641 2148 2697 2204
rect 2697 2148 2701 2204
rect 2637 2144 2701 2148
rect 5288 2204 5352 2208
rect 5288 2148 5292 2204
rect 5292 2148 5348 2204
rect 5348 2148 5352 2204
rect 5288 2144 5352 2148
rect 5368 2204 5432 2208
rect 5368 2148 5372 2204
rect 5372 2148 5428 2204
rect 5428 2148 5432 2204
rect 5368 2144 5432 2148
rect 5448 2204 5512 2208
rect 5448 2148 5452 2204
rect 5452 2148 5508 2204
rect 5508 2148 5512 2204
rect 5448 2144 5512 2148
rect 5528 2204 5592 2208
rect 5528 2148 5532 2204
rect 5532 2148 5588 2204
rect 5588 2148 5592 2204
rect 5528 2144 5592 2148
rect 8178 2204 8242 2208
rect 8178 2148 8182 2204
rect 8182 2148 8238 2204
rect 8238 2148 8242 2204
rect 8178 2144 8242 2148
rect 8258 2204 8322 2208
rect 8258 2148 8262 2204
rect 8262 2148 8318 2204
rect 8318 2148 8322 2204
rect 8258 2144 8322 2148
rect 8338 2204 8402 2208
rect 8338 2148 8342 2204
rect 8342 2148 8398 2204
rect 8398 2148 8402 2204
rect 8338 2144 8402 2148
rect 8418 2204 8482 2208
rect 8418 2148 8422 2204
rect 8422 2148 8478 2204
rect 8478 2148 8482 2204
rect 8418 2144 8482 2148
<< metal4 >>
rect 2389 21792 2709 22352
rect 2389 21728 2397 21792
rect 2461 21728 2477 21792
rect 2541 21728 2557 21792
rect 2621 21728 2637 21792
rect 2701 21728 2709 21792
rect 2389 20704 2709 21728
rect 2389 20640 2397 20704
rect 2461 20640 2477 20704
rect 2541 20640 2557 20704
rect 2621 20640 2637 20704
rect 2701 20640 2709 20704
rect 2389 19616 2709 20640
rect 2389 19552 2397 19616
rect 2461 19552 2477 19616
rect 2541 19552 2557 19616
rect 2621 19552 2637 19616
rect 2701 19552 2709 19616
rect 2389 18528 2709 19552
rect 2389 18464 2397 18528
rect 2461 18464 2477 18528
rect 2541 18464 2557 18528
rect 2621 18464 2637 18528
rect 2701 18464 2709 18528
rect 2389 17440 2709 18464
rect 2389 17376 2397 17440
rect 2461 17376 2477 17440
rect 2541 17376 2557 17440
rect 2621 17376 2637 17440
rect 2701 17376 2709 17440
rect 2389 16352 2709 17376
rect 2389 16288 2397 16352
rect 2461 16288 2477 16352
rect 2541 16288 2557 16352
rect 2621 16288 2637 16352
rect 2701 16288 2709 16352
rect 2389 15264 2709 16288
rect 2389 15200 2397 15264
rect 2461 15200 2477 15264
rect 2541 15200 2557 15264
rect 2621 15200 2637 15264
rect 2701 15200 2709 15264
rect 2389 14176 2709 15200
rect 2389 14112 2397 14176
rect 2461 14112 2477 14176
rect 2541 14112 2557 14176
rect 2621 14112 2637 14176
rect 2701 14112 2709 14176
rect 2389 13088 2709 14112
rect 2389 13024 2397 13088
rect 2461 13024 2477 13088
rect 2541 13024 2557 13088
rect 2621 13024 2637 13088
rect 2701 13024 2709 13088
rect 2389 12000 2709 13024
rect 2389 11936 2397 12000
rect 2461 11936 2477 12000
rect 2541 11936 2557 12000
rect 2621 11936 2637 12000
rect 2701 11936 2709 12000
rect 2389 10912 2709 11936
rect 2389 10848 2397 10912
rect 2461 10848 2477 10912
rect 2541 10848 2557 10912
rect 2621 10848 2637 10912
rect 2701 10848 2709 10912
rect 2389 9824 2709 10848
rect 2389 9760 2397 9824
rect 2461 9760 2477 9824
rect 2541 9760 2557 9824
rect 2621 9760 2637 9824
rect 2701 9760 2709 9824
rect 2389 8736 2709 9760
rect 2389 8672 2397 8736
rect 2461 8672 2477 8736
rect 2541 8672 2557 8736
rect 2621 8672 2637 8736
rect 2701 8672 2709 8736
rect 2389 7648 2709 8672
rect 2389 7584 2397 7648
rect 2461 7584 2477 7648
rect 2541 7584 2557 7648
rect 2621 7584 2637 7648
rect 2701 7584 2709 7648
rect 2389 6560 2709 7584
rect 2389 6496 2397 6560
rect 2461 6496 2477 6560
rect 2541 6496 2557 6560
rect 2621 6496 2637 6560
rect 2701 6496 2709 6560
rect 2389 5472 2709 6496
rect 2389 5408 2397 5472
rect 2461 5408 2477 5472
rect 2541 5408 2557 5472
rect 2621 5408 2637 5472
rect 2701 5408 2709 5472
rect 2389 4384 2709 5408
rect 2389 4320 2397 4384
rect 2461 4320 2477 4384
rect 2541 4320 2557 4384
rect 2621 4320 2637 4384
rect 2701 4320 2709 4384
rect 2389 3296 2709 4320
rect 2389 3232 2397 3296
rect 2461 3232 2477 3296
rect 2541 3232 2557 3296
rect 2621 3232 2637 3296
rect 2701 3232 2709 3296
rect 2389 2208 2709 3232
rect 2389 2144 2397 2208
rect 2461 2144 2477 2208
rect 2541 2144 2557 2208
rect 2621 2144 2637 2208
rect 2701 2144 2709 2208
rect 2389 2128 2709 2144
rect 3834 22336 4155 22352
rect 3834 22272 3842 22336
rect 3906 22272 3922 22336
rect 3986 22272 4002 22336
rect 4066 22272 4082 22336
rect 4146 22272 4155 22336
rect 3834 21248 4155 22272
rect 3834 21184 3842 21248
rect 3906 21184 3922 21248
rect 3986 21184 4002 21248
rect 4066 21184 4082 21248
rect 4146 21184 4155 21248
rect 3834 20160 4155 21184
rect 3834 20096 3842 20160
rect 3906 20096 3922 20160
rect 3986 20096 4002 20160
rect 4066 20096 4082 20160
rect 4146 20096 4155 20160
rect 3834 19072 4155 20096
rect 3834 19008 3842 19072
rect 3906 19008 3922 19072
rect 3986 19008 4002 19072
rect 4066 19008 4082 19072
rect 4146 19008 4155 19072
rect 3834 17984 4155 19008
rect 3834 17920 3842 17984
rect 3906 17920 3922 17984
rect 3986 17920 4002 17984
rect 4066 17920 4082 17984
rect 4146 17920 4155 17984
rect 3834 16896 4155 17920
rect 3834 16832 3842 16896
rect 3906 16832 3922 16896
rect 3986 16832 4002 16896
rect 4066 16832 4082 16896
rect 4146 16832 4155 16896
rect 3834 15808 4155 16832
rect 3834 15744 3842 15808
rect 3906 15744 3922 15808
rect 3986 15744 4002 15808
rect 4066 15744 4082 15808
rect 4146 15744 4155 15808
rect 3834 14720 4155 15744
rect 3834 14656 3842 14720
rect 3906 14656 3922 14720
rect 3986 14656 4002 14720
rect 4066 14656 4082 14720
rect 4146 14656 4155 14720
rect 3834 13632 4155 14656
rect 3834 13568 3842 13632
rect 3906 13568 3922 13632
rect 3986 13568 4002 13632
rect 4066 13568 4082 13632
rect 4146 13568 4155 13632
rect 3834 12544 4155 13568
rect 3834 12480 3842 12544
rect 3906 12480 3922 12544
rect 3986 12480 4002 12544
rect 4066 12480 4082 12544
rect 4146 12480 4155 12544
rect 3834 11456 4155 12480
rect 3834 11392 3842 11456
rect 3906 11392 3922 11456
rect 3986 11392 4002 11456
rect 4066 11392 4082 11456
rect 4146 11392 4155 11456
rect 3834 10368 4155 11392
rect 3834 10304 3842 10368
rect 3906 10304 3922 10368
rect 3986 10304 4002 10368
rect 4066 10304 4082 10368
rect 4146 10304 4155 10368
rect 3834 9280 4155 10304
rect 3834 9216 3842 9280
rect 3906 9216 3922 9280
rect 3986 9216 4002 9280
rect 4066 9216 4082 9280
rect 4146 9216 4155 9280
rect 3834 8192 4155 9216
rect 3834 8128 3842 8192
rect 3906 8128 3922 8192
rect 3986 8128 4002 8192
rect 4066 8128 4082 8192
rect 4146 8128 4155 8192
rect 3834 7104 4155 8128
rect 3834 7040 3842 7104
rect 3906 7040 3922 7104
rect 3986 7040 4002 7104
rect 4066 7040 4082 7104
rect 4146 7040 4155 7104
rect 3834 6016 4155 7040
rect 3834 5952 3842 6016
rect 3906 5952 3922 6016
rect 3986 5952 4002 6016
rect 4066 5952 4082 6016
rect 4146 5952 4155 6016
rect 3834 4928 4155 5952
rect 3834 4864 3842 4928
rect 3906 4864 3922 4928
rect 3986 4864 4002 4928
rect 4066 4864 4082 4928
rect 4146 4864 4155 4928
rect 3834 3840 4155 4864
rect 3834 3776 3842 3840
rect 3906 3776 3922 3840
rect 3986 3776 4002 3840
rect 4066 3776 4082 3840
rect 4146 3776 4155 3840
rect 3834 2752 4155 3776
rect 3834 2688 3842 2752
rect 3906 2688 3922 2752
rect 3986 2688 4002 2752
rect 4066 2688 4082 2752
rect 4146 2688 4155 2752
rect 3834 2128 4155 2688
rect 5280 21792 5600 22352
rect 5280 21728 5288 21792
rect 5352 21728 5368 21792
rect 5432 21728 5448 21792
rect 5512 21728 5528 21792
rect 5592 21728 5600 21792
rect 5280 20704 5600 21728
rect 5280 20640 5288 20704
rect 5352 20640 5368 20704
rect 5432 20640 5448 20704
rect 5512 20640 5528 20704
rect 5592 20640 5600 20704
rect 5280 19616 5600 20640
rect 5280 19552 5288 19616
rect 5352 19552 5368 19616
rect 5432 19552 5448 19616
rect 5512 19552 5528 19616
rect 5592 19552 5600 19616
rect 5280 18528 5600 19552
rect 5280 18464 5288 18528
rect 5352 18464 5368 18528
rect 5432 18464 5448 18528
rect 5512 18464 5528 18528
rect 5592 18464 5600 18528
rect 5280 17440 5600 18464
rect 5280 17376 5288 17440
rect 5352 17376 5368 17440
rect 5432 17376 5448 17440
rect 5512 17376 5528 17440
rect 5592 17376 5600 17440
rect 5280 16352 5600 17376
rect 5280 16288 5288 16352
rect 5352 16288 5368 16352
rect 5432 16288 5448 16352
rect 5512 16288 5528 16352
rect 5592 16288 5600 16352
rect 5280 15264 5600 16288
rect 5280 15200 5288 15264
rect 5352 15200 5368 15264
rect 5432 15200 5448 15264
rect 5512 15200 5528 15264
rect 5592 15200 5600 15264
rect 5280 14176 5600 15200
rect 5280 14112 5288 14176
rect 5352 14112 5368 14176
rect 5432 14112 5448 14176
rect 5512 14112 5528 14176
rect 5592 14112 5600 14176
rect 5280 13088 5600 14112
rect 5280 13024 5288 13088
rect 5352 13024 5368 13088
rect 5432 13024 5448 13088
rect 5512 13024 5528 13088
rect 5592 13024 5600 13088
rect 5280 12000 5600 13024
rect 5280 11936 5288 12000
rect 5352 11936 5368 12000
rect 5432 11936 5448 12000
rect 5512 11936 5528 12000
rect 5592 11936 5600 12000
rect 5280 10912 5600 11936
rect 5280 10848 5288 10912
rect 5352 10848 5368 10912
rect 5432 10848 5448 10912
rect 5512 10848 5528 10912
rect 5592 10848 5600 10912
rect 5280 9824 5600 10848
rect 5280 9760 5288 9824
rect 5352 9760 5368 9824
rect 5432 9760 5448 9824
rect 5512 9760 5528 9824
rect 5592 9760 5600 9824
rect 5280 8736 5600 9760
rect 5280 8672 5288 8736
rect 5352 8672 5368 8736
rect 5432 8672 5448 8736
rect 5512 8672 5528 8736
rect 5592 8672 5600 8736
rect 5280 7648 5600 8672
rect 5280 7584 5288 7648
rect 5352 7584 5368 7648
rect 5432 7584 5448 7648
rect 5512 7584 5528 7648
rect 5592 7584 5600 7648
rect 5280 6560 5600 7584
rect 5280 6496 5288 6560
rect 5352 6496 5368 6560
rect 5432 6496 5448 6560
rect 5512 6496 5528 6560
rect 5592 6496 5600 6560
rect 5280 5472 5600 6496
rect 5280 5408 5288 5472
rect 5352 5408 5368 5472
rect 5432 5408 5448 5472
rect 5512 5408 5528 5472
rect 5592 5408 5600 5472
rect 5280 4384 5600 5408
rect 5280 4320 5288 4384
rect 5352 4320 5368 4384
rect 5432 4320 5448 4384
rect 5512 4320 5528 4384
rect 5592 4320 5600 4384
rect 5280 3296 5600 4320
rect 5280 3232 5288 3296
rect 5352 3232 5368 3296
rect 5432 3232 5448 3296
rect 5512 3232 5528 3296
rect 5592 3232 5600 3296
rect 5280 2208 5600 3232
rect 5280 2144 5288 2208
rect 5352 2144 5368 2208
rect 5432 2144 5448 2208
rect 5512 2144 5528 2208
rect 5592 2144 5600 2208
rect 5280 2128 5600 2144
rect 6725 22336 7045 22352
rect 6725 22272 6733 22336
rect 6797 22272 6813 22336
rect 6877 22272 6893 22336
rect 6957 22272 6973 22336
rect 7037 22272 7045 22336
rect 6725 21248 7045 22272
rect 6725 21184 6733 21248
rect 6797 21184 6813 21248
rect 6877 21184 6893 21248
rect 6957 21184 6973 21248
rect 7037 21184 7045 21248
rect 6725 20160 7045 21184
rect 6725 20096 6733 20160
rect 6797 20096 6813 20160
rect 6877 20096 6893 20160
rect 6957 20096 6973 20160
rect 7037 20096 7045 20160
rect 6725 19072 7045 20096
rect 6725 19008 6733 19072
rect 6797 19008 6813 19072
rect 6877 19008 6893 19072
rect 6957 19008 6973 19072
rect 7037 19008 7045 19072
rect 6725 17984 7045 19008
rect 6725 17920 6733 17984
rect 6797 17920 6813 17984
rect 6877 17920 6893 17984
rect 6957 17920 6973 17984
rect 7037 17920 7045 17984
rect 6725 16896 7045 17920
rect 6725 16832 6733 16896
rect 6797 16832 6813 16896
rect 6877 16832 6893 16896
rect 6957 16832 6973 16896
rect 7037 16832 7045 16896
rect 6725 15808 7045 16832
rect 6725 15744 6733 15808
rect 6797 15744 6813 15808
rect 6877 15744 6893 15808
rect 6957 15744 6973 15808
rect 7037 15744 7045 15808
rect 6725 14720 7045 15744
rect 6725 14656 6733 14720
rect 6797 14656 6813 14720
rect 6877 14656 6893 14720
rect 6957 14656 6973 14720
rect 7037 14656 7045 14720
rect 6725 13632 7045 14656
rect 6725 13568 6733 13632
rect 6797 13568 6813 13632
rect 6877 13568 6893 13632
rect 6957 13568 6973 13632
rect 7037 13568 7045 13632
rect 6725 12544 7045 13568
rect 6725 12480 6733 12544
rect 6797 12480 6813 12544
rect 6877 12480 6893 12544
rect 6957 12480 6973 12544
rect 7037 12480 7045 12544
rect 6725 11456 7045 12480
rect 6725 11392 6733 11456
rect 6797 11392 6813 11456
rect 6877 11392 6893 11456
rect 6957 11392 6973 11456
rect 7037 11392 7045 11456
rect 6725 10368 7045 11392
rect 6725 10304 6733 10368
rect 6797 10304 6813 10368
rect 6877 10304 6893 10368
rect 6957 10304 6973 10368
rect 7037 10304 7045 10368
rect 6725 9280 7045 10304
rect 6725 9216 6733 9280
rect 6797 9216 6813 9280
rect 6877 9216 6893 9280
rect 6957 9216 6973 9280
rect 7037 9216 7045 9280
rect 6725 8192 7045 9216
rect 6725 8128 6733 8192
rect 6797 8128 6813 8192
rect 6877 8128 6893 8192
rect 6957 8128 6973 8192
rect 7037 8128 7045 8192
rect 6725 7104 7045 8128
rect 6725 7040 6733 7104
rect 6797 7040 6813 7104
rect 6877 7040 6893 7104
rect 6957 7040 6973 7104
rect 7037 7040 7045 7104
rect 6725 6016 7045 7040
rect 6725 5952 6733 6016
rect 6797 5952 6813 6016
rect 6877 5952 6893 6016
rect 6957 5952 6973 6016
rect 7037 5952 7045 6016
rect 6725 4928 7045 5952
rect 6725 4864 6733 4928
rect 6797 4864 6813 4928
rect 6877 4864 6893 4928
rect 6957 4864 6973 4928
rect 7037 4864 7045 4928
rect 6725 3840 7045 4864
rect 6725 3776 6733 3840
rect 6797 3776 6813 3840
rect 6877 3776 6893 3840
rect 6957 3776 6973 3840
rect 7037 3776 7045 3840
rect 6725 2752 7045 3776
rect 6725 2688 6733 2752
rect 6797 2688 6813 2752
rect 6877 2688 6893 2752
rect 6957 2688 6973 2752
rect 7037 2688 7045 2752
rect 6725 2128 7045 2688
rect 8170 21792 8490 22352
rect 8170 21728 8178 21792
rect 8242 21728 8258 21792
rect 8322 21728 8338 21792
rect 8402 21728 8418 21792
rect 8482 21728 8490 21792
rect 8170 20704 8490 21728
rect 8170 20640 8178 20704
rect 8242 20640 8258 20704
rect 8322 20640 8338 20704
rect 8402 20640 8418 20704
rect 8482 20640 8490 20704
rect 8170 19616 8490 20640
rect 8170 19552 8178 19616
rect 8242 19552 8258 19616
rect 8322 19552 8338 19616
rect 8402 19552 8418 19616
rect 8482 19552 8490 19616
rect 8170 18528 8490 19552
rect 8170 18464 8178 18528
rect 8242 18464 8258 18528
rect 8322 18464 8338 18528
rect 8402 18464 8418 18528
rect 8482 18464 8490 18528
rect 8170 17440 8490 18464
rect 8170 17376 8178 17440
rect 8242 17376 8258 17440
rect 8322 17376 8338 17440
rect 8402 17376 8418 17440
rect 8482 17376 8490 17440
rect 8170 16352 8490 17376
rect 8170 16288 8178 16352
rect 8242 16288 8258 16352
rect 8322 16288 8338 16352
rect 8402 16288 8418 16352
rect 8482 16288 8490 16352
rect 8170 15264 8490 16288
rect 8170 15200 8178 15264
rect 8242 15200 8258 15264
rect 8322 15200 8338 15264
rect 8402 15200 8418 15264
rect 8482 15200 8490 15264
rect 8170 14176 8490 15200
rect 8170 14112 8178 14176
rect 8242 14112 8258 14176
rect 8322 14112 8338 14176
rect 8402 14112 8418 14176
rect 8482 14112 8490 14176
rect 8170 13088 8490 14112
rect 8170 13024 8178 13088
rect 8242 13024 8258 13088
rect 8322 13024 8338 13088
rect 8402 13024 8418 13088
rect 8482 13024 8490 13088
rect 8170 12000 8490 13024
rect 8170 11936 8178 12000
rect 8242 11936 8258 12000
rect 8322 11936 8338 12000
rect 8402 11936 8418 12000
rect 8482 11936 8490 12000
rect 8170 10912 8490 11936
rect 8170 10848 8178 10912
rect 8242 10848 8258 10912
rect 8322 10848 8338 10912
rect 8402 10848 8418 10912
rect 8482 10848 8490 10912
rect 8170 9824 8490 10848
rect 8170 9760 8178 9824
rect 8242 9760 8258 9824
rect 8322 9760 8338 9824
rect 8402 9760 8418 9824
rect 8482 9760 8490 9824
rect 8170 8736 8490 9760
rect 8170 8672 8178 8736
rect 8242 8672 8258 8736
rect 8322 8672 8338 8736
rect 8402 8672 8418 8736
rect 8482 8672 8490 8736
rect 8170 7648 8490 8672
rect 8170 7584 8178 7648
rect 8242 7584 8258 7648
rect 8322 7584 8338 7648
rect 8402 7584 8418 7648
rect 8482 7584 8490 7648
rect 8170 6560 8490 7584
rect 8170 6496 8178 6560
rect 8242 6496 8258 6560
rect 8322 6496 8338 6560
rect 8402 6496 8418 6560
rect 8482 6496 8490 6560
rect 8170 5472 8490 6496
rect 8170 5408 8178 5472
rect 8242 5408 8258 5472
rect 8322 5408 8338 5472
rect 8402 5408 8418 5472
rect 8482 5408 8490 5472
rect 8170 4384 8490 5408
rect 8170 4320 8178 4384
rect 8242 4320 8258 4384
rect 8322 4320 8338 4384
rect 8402 4320 8418 4384
rect 8482 4320 8490 4384
rect 8170 3296 8490 4320
rect 8170 3232 8178 3296
rect 8242 3232 8258 3296
rect 8322 3232 8338 3296
rect 8402 3232 8418 3296
rect 8482 3232 8490 3296
rect 8170 2208 8490 3232
rect 8170 2144 8178 2208
rect 8242 2144 8258 2208
rect 8322 2144 8338 2208
rect 8402 2144 8418 2208
rect 8482 2144 8490 2208
rect 8170 2128 8490 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607194113
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607194113
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607194113
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607194113
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1607194113
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607194113
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607194113
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607194113
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607194113
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1607194113
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1607194113
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1607194113
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1607194113
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607194113
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 9384 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1607194113
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87
timestamp 1607194113
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607194113
transform -1 0 9752 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607194113
transform -1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607194113
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607194113
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607194113
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607194113
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607194113
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1607194113
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607194113
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607194113
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_80
timestamp 1607194113
transform 1 0 8464 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607194113
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp 1607194113
transform 1 0 9200 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607194113
transform -1 0 9752 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1607194113
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1607194113
transform 1 0 2484 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1607194113
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1607194113
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_LEFT1a_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607194113
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[1\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2576 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  LEFT1a
timestamp 1607194113
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_36
timestamp 1607194113
transform 1 0 4416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_24
timestamp 1607194113
transform 1 0 3312 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[1\]_A
timestamp 1607194113
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1607194113
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1607194113
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_48
timestamp 1607194113
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1607194113
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1607194113
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1607194113
transform 1 0 7912 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  LEFT2a
timestamp 1607194113
transform 1 0 8280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_90
timestamp 1607194113
transform 1 0 9384 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1607194113
transform 1 0 9016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_LEFT2a_A
timestamp 1607194113
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607194113
transform -1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607194113
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607194113
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607194113
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607194113
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607194113
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1607194113
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1607194113
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1607194113
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_80
timestamp 1607194113
transform 1 0 8464 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1607194113
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp 1607194113
transform 1 0 9200 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607194113
transform -1 0 9752 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1607194113
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607194113
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607194113
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1607194113
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1607194113
transform 1 0 4140 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_27
timestamp 1607194113
transform 1 0 3588 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[9\]_A
timestamp 1607194113
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[9\]
timestamp 1607194113
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1607194113
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1607194113
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_54
timestamp 1607194113
transform 1 0 6072 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1607194113
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1607194113
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp 1607194113
transform 1 0 8556 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_78
timestamp 1607194113
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1607194113
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[7\]_A
timestamp 1607194113
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1607194113
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607194113
transform -1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1607194113
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607194113
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607194113
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607194113
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607194113
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607194113
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1607194113
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1607194113
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1607194113
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607194113
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1607194113
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1607194113
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1607194113
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1607194113
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1607194113
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1607194113
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[10\]
timestamp 1607194113
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_82
timestamp 1607194113
transform 1 0 8648 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1607194113
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_66
timestamp 1607194113
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_83
timestamp 1607194113
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_76
timestamp 1607194113
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_68
timestamp 1607194113
transform 1 0 7360 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[10\]_A
timestamp 1607194113
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[7\]
timestamp 1607194113
transform 1 0 8372 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_90
timestamp 1607194113
transform 1 0 9384 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607194113
transform -1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607194113
transform -1 0 9752 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607194113
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607194113
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607194113
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607194113
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607194113
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1607194113
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1607194113
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1607194113
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_80
timestamp 1607194113
transform 1 0 8464 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1607194113
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp 1607194113
transform 1 0 9200 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607194113
transform -1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_14
timestamp 1607194113
transform 1 0 2392 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1607194113
transform 1 0 2116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1607194113
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[5\]_A
timestamp 1607194113
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607194113
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_38
timestamp 1607194113
transform 1 0 4600 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_26
timestamp 1607194113
transform 1 0 3496 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1607194113
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1607194113
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_52
timestamp 1607194113
transform 1 0 5888 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_CLKBUF_0_A
timestamp 1607194113
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1607194113
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1607194113
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_90
timestamp 1607194113
transform 1 0 9384 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1607194113
transform 1 0 9016 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607194113
transform -1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_16
timestamp 1607194113
transform 1 0 2576 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1607194113
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1607194113
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607194113
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[5\]
timestamp 1607194113
transform 1 0 2208 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1607194113
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1607194113
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1607194113
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_44
timestamp 1607194113
transform 1 0 5152 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  CLKBUF_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5704 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_10_82
timestamp 1607194113
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_70
timestamp 1607194113
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_90
timestamp 1607194113
transform 1 0 9384 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607194113
transform -1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1607194113
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607194113
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607194113
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1607194113
transform 1 0 4692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1607194113
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1607194113
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1607194113
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1607194113
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 1607194113
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_CLKBUF_3_A
timestamp 1607194113
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1607194113
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1607194113
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_90
timestamp 1607194113
transform 1 0 9384 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1607194113
transform 1 0 9016 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607194113
transform -1 0 9752 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607194113
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607194113
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607194113
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1607194113
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607194113
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1607194113
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_44
timestamp 1607194113
transform 1 0 5152 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  CLKBUF_3
timestamp 1607194113
transform 1 0 5704 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_12_82
timestamp 1607194113
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_70
timestamp 1607194113
transform 1 0 7544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_90
timestamp 1607194113
transform 1 0 9384 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607194113
transform -1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607194113
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607194113
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1607194113
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607194113
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607194113
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607194113
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607194113
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607194113
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1607194113
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1607194113
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1607194113
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1607194113
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1607194113
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1607194113
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1607194113
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1607194113
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1607194113
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_80
timestamp 1607194113
transform 1 0 8464 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1607194113
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1607194113
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_88
timestamp 1607194113
transform 1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_90
timestamp 1607194113
transform 1 0 9384 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1607194113
transform 1 0 9016 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607194113
transform -1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607194113
transform -1 0 9752 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1607194113
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607194113
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607194113
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1607194113
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1607194113
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1607194113
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1607194113
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1607194113
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1607194113
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1607194113
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_78
timestamp 1607194113
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1607194113
transform 1 0 7912 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1607194113
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1607194113
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[3\]_A
timestamp 1607194113
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_CLKBUF_A
timestamp 1607194113
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[11\]
timestamp 1607194113
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  CLKBUF $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1607194113
transform 1 0 9108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[11\]_A
timestamp 1607194113
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607194113
transform -1 0 9752 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607194113
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607194113
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607194113
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607194113
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607194113
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1607194113
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1607194113
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1607194113
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1607194113
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_79
timestamp 1607194113
transform 1 0 8372 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_67
timestamp 1607194113
transform 1 0 7268 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[3\]
timestamp 1607194113
transform 1 0 6900 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607194113
transform -1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1607194113
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607194113
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607194113
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_31
timestamp 1607194113
transform 1 0 3956 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1607194113
transform 1 0 3588 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  ZEROA $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_4  LEFT2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 4416 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  LEFT1
timestamp 1607194113
transform 1 0 4048 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1607194113
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1607194113
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1607194113
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1607194113
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  RIGHT2
timestamp 1607194113
transform 1 0 5428 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  RIGHT1
timestamp 1607194113
transform 1 0 5060 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1607194113
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_90
timestamp 1607194113
transform 1 0 9384 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1607194113
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607194113
transform -1 0 9752 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607194113
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607194113
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607194113
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607194113
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607194113
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1607194113
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1607194113
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1607194113
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_80
timestamp 1607194113
transform 1 0 8464 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1607194113
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_88
timestamp 1607194113
transform 1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607194113
transform -1 0 9752 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607194113
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607194113
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1607194113
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607194113
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607194113
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607194113
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607194113
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607194113
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1607194113
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1607194113
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1607194113
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1607194113
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1607194113
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1607194113
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1607194113
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1607194113
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[4\]
timestamp 1607194113
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_80
timestamp 1607194113
transform 1 0 8464 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1607194113
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_83
timestamp 1607194113
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_78
timestamp 1607194113
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_70
timestamp 1607194113
transform 1 0 7544 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1607194113
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[4\]_A
timestamp 1607194113
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[0\]
timestamp 1607194113
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_88
timestamp 1607194113
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_87
timestamp 1607194113
transform 1 0 9108 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[0\]_A
timestamp 1607194113
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607194113
transform -1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607194113
transform -1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1607194113
transform 1 0 2852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_7
timestamp 1607194113
transform 1 0 1748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1607194113
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[6\]_A
timestamp 1607194113
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607194113
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1607194113
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1607194113
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1607194113
transform 1 0 5060 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1607194113
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  CLKBUF_2
timestamp 1607194113
transform 1 0 6808 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_21_82
timestamp 1607194113
transform 1 0 8648 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_90
timestamp 1607194113
transform 1 0 9384 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607194113
transform -1 0 9752 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_19
timestamp 1607194113
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_7
timestamp 1607194113
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607194113
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[6\]
timestamp 1607194113
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607194113
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1607194113
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1607194113
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1607194113
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_CLKBUF_2_A
timestamp 1607194113
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_76
timestamp 1607194113
transform 1 0 8096 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_64
timestamp 1607194113
transform 1 0 6992 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_88
timestamp 1607194113
transform 1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607194113
transform -1 0 9752 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_20
timestamp 1607194113
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1607194113
transform 1 0 2484 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607194113
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607194113
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[2\]
timestamp 1607194113
transform 1 0 2576 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1607194113
transform 1 0 4416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_24
timestamp 1607194113
transform 1 0 3312 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[2\]_A
timestamp 1607194113
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1607194113
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1607194113
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_48
timestamp 1607194113
transform 1 0 5520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1607194113
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1607194113
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_90
timestamp 1607194113
transform 1 0 9384 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_86
timestamp 1607194113
transform 1 0 9016 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607194113
transform -1 0 9752 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607194113
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607194113
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607194113
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1607194113
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607194113
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1607194113
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1607194113
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1607194113
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_80
timestamp 1607194113
transform 1 0 8464 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1607194113
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_88
timestamp 1607194113
transform 1 0 9200 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607194113
transform -1 0 9752 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1607194113
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607194113
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607194113
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1607194113
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1607194113
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1607194113
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607194113
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1607194113
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1607194113
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1607194113
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_90
timestamp 1607194113
transform 1 0 9384 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1607194113
transform 1 0 9016 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607194113
transform -1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1607194113
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607194113
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607194113
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607194113
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607194113
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607194113
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1607194113
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1607194113
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607194113
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607194113
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1607194113
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1607194113
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1607194113
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1607194113
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1607194113
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607194113
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1607194113
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1607194113
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_80
timestamp 1607194113
transform 1 0 8464 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1607194113
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_90
timestamp 1607194113
transform 1 0 9384 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_86
timestamp 1607194113
transform 1 0 9016 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_88
timestamp 1607194113
transform 1 0 9200 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607194113
transform -1 0 9752 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607194113
transform -1 0 9752 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1607194113
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607194113
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607194113
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1607194113
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1607194113
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1607194113
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1607194113
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1607194113
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_80
timestamp 1607194113
transform 1 0 8464 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1607194113
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_88
timestamp 1607194113
transform 1 0 9200 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607194113
transform -1 0 9752 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1607194113
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1607194113
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607194113
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_27
timestamp 1607194113
transform 1 0 3588 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  CLKBUF_1
timestamp 1607194113
transform 1 0 4140 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1607194113
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1607194113
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1607194113
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1607194113
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_78
timestamp 1607194113
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 1607194113
transform 1 0 7912 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  RIGHT2a\[8\]
timestamp 1607194113
transform 1 0 8372 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 1607194113
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT2a\[8\]_A
timestamp 1607194113
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607194113
transform -1 0 9752 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607194113
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607194113
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607194113
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_36
timestamp 1607194113
transform 1 0 4416 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1607194113
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607194113
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_CLKBUF_1_A
timestamp 1607194113
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1607194113
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_60
timestamp 1607194113
transform 1 0 6624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_48
timestamp 1607194113
transform 1 0 5520 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1607194113
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_90
timestamp 1607194113
transform 1 0 9384 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_84
timestamp 1607194113
transform 1 0 8832 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607194113
transform -1 0 9752 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1607194113
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607194113
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607194113
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1607194113
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1607194113
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1607194113
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1607194113
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1607194113
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1607194113
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1607194113
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_90
timestamp 1607194113
transform 1 0 9384 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_86
timestamp 1607194113
transform 1 0 9016 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607194113
transform -1 0 9752 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1607194113
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607194113
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607194113
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1607194113
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1607194113
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1607194113
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1607194113
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1607194113
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_80
timestamp 1607194113
transform 1 0 8464 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1607194113
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_88
timestamp 1607194113
transform 1 0 9200 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607194113
transform -1 0 9752 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607194113
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607194113
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1607194113
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607194113
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607194113
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607194113
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1607194113
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607194113
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1607194113
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1607194113
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1607194113
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1607194113
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1607194113
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_62
timestamp 1607194113
transform 1 0 6808 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1607194113
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1607194113
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1607194113
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_80
timestamp 1607194113
transform 1 0 8464 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1607194113
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_76
timestamp 1607194113
transform 1 0 8096 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_72
timestamp 1607194113
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_RIGHT1a_A
timestamp 1607194113
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  RIGHT1a
timestamp 1607194113
transform 1 0 7360 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_88
timestamp 1607194113
transform 1 0 9200 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_88
timestamp 1607194113
transform 1 0 9200 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607194113
transform -1 0 9752 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607194113
transform -1 0 9752 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1607194113
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1607194113
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607194113
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1607194113
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1607194113
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1607194113
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1607194113
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1607194113
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1607194113
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1607194113
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_90
timestamp 1607194113
transform 1 0 9384 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1607194113
transform 1 0 9016 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607194113
transform -1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1607194113
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607194113
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607194113
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1607194113
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1607194113
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1607194113
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_56
timestamp 1607194113
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1607194113
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1607194113
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_75
timestamp 1607194113
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_63
timestamp 1607194113
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1607194113
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607194113
transform -1 0 9752 0 -1 22304
box -38 -48 314 592
<< labels >>
rlabel metal2 s 8942 0 8998 800 6 clk_i
port 0 nsew default input
rlabel metal2 s 1766 0 1822 800 6 clk_o[0]
port 1 nsew default tristate
rlabel metal3 s 10080 824 10880 944 6 clk_o[1]
port 2 nsew default tristate
rlabel metal2 s 2686 23680 2742 24480 6 clk_o[2]
port 3 nsew default tristate
rlabel metal3 s 0 4088 800 4208 6 clk_o[3]
port 4 nsew default tristate
rlabel metal3 s 10080 2592 10880 2712 6 e_o[0]
port 5 nsew default tristate
rlabel metal3 s 10080 21496 10880 21616 6 e_o[10]
port 6 nsew default tristate
rlabel metal3 s 10080 23400 10880 23520 6 e_o[11]
port 7 nsew default tristate
rlabel metal3 s 10080 4496 10880 4616 6 e_o[1]
port 8 nsew default tristate
rlabel metal3 s 10080 6400 10880 6520 6 e_o[2]
port 9 nsew default tristate
rlabel metal3 s 10080 8304 10880 8424 6 e_o[3]
port 10 nsew default tristate
rlabel metal3 s 10080 10208 10880 10328 6 e_o[4]
port 11 nsew default tristate
rlabel metal3 s 10080 12112 10880 12232 6 e_o[5]
port 12 nsew default tristate
rlabel metal3 s 10080 13880 10880 14000 6 e_o[6]
port 13 nsew default tristate
rlabel metal3 s 10080 15784 10880 15904 6 e_o[7]
port 14 nsew default tristate
rlabel metal3 s 10080 17688 10880 17808 6 e_o[8]
port 15 nsew default tristate
rlabel metal3 s 10080 19592 10880 19712 6 e_o[9]
port 16 nsew default tristate
rlabel metal3 s 0 20408 800 20528 6 n1_o
port 17 nsew default tristate
rlabel metal2 s 8114 23680 8170 24480 6 n_o
port 18 nsew default tristate
rlabel metal2 s 5354 0 5410 800 6 s_o
port 19 nsew default tristate
rlabel metal3 s 0 12248 800 12368 6 w_o
port 20 nsew default tristate
rlabel metal4 s 2389 2128 2709 22352 6 VPWR
port 21 nsew default input
rlabel metal4 s 3835 2128 4155 22352 6 VGND
port 22 nsew default input
<< properties >>
string FIXED_BBOX 0 0 10880 24480
<< end >>
