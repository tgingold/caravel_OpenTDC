magic
tech sky130A
magscale 1 2
timestamp 1607276172
<< locali >>
rect 31953 45815 31987 46121
rect 45937 44183 45971 44285
rect 51549 42211 51583 42313
rect 12449 41055 12483 41157
rect 29377 41123 29411 41225
rect 9873 40919 9907 41021
rect 40049 40987 40083 41225
rect 9505 40443 9539 40545
rect 14657 38879 14691 39049
rect 26525 38199 26559 38301
rect 40693 38199 40727 38369
rect 16129 37655 16163 37757
rect 20361 37655 20395 37757
rect 23673 37723 23707 37961
rect 16957 35139 16991 35241
rect 43177 34935 43211 35037
rect 48789 34935 48823 35241
rect 55321 35071 55355 35241
rect 55321 34935 55355 35037
rect 40325 34595 40359 34697
rect 67741 34527 67775 34697
rect 21649 33847 21683 34017
rect 37565 33847 37599 33949
rect 31493 32759 31527 32861
rect 54401 31875 54435 31977
rect 12173 31263 12207 31433
rect 23765 31263 23799 31365
rect 57161 31331 57195 31433
rect 36921 30651 36955 30889
rect 51273 29495 51307 29665
rect 71237 29563 71271 29665
rect 13553 28407 13587 28713
rect 15301 28407 15335 28645
rect 14105 26843 14139 27013
rect 9505 22967 9539 23205
rect 12817 19159 12851 19261
rect 23949 18819 23983 18921
<< viali >>
rect 8401 47617 8435 47651
rect 7941 47549 7975 47583
rect 8493 47549 8527 47583
rect 7757 47209 7791 47243
rect 22477 47209 22511 47243
rect 4537 47073 4571 47107
rect 7941 47073 7975 47107
rect 8217 47073 8251 47107
rect 8585 47073 8619 47107
rect 12449 47073 12483 47107
rect 13001 47073 13035 47107
rect 13185 47073 13219 47107
rect 22661 47073 22695 47107
rect 22845 47073 22879 47107
rect 23397 47073 23431 47107
rect 23581 47073 23615 47107
rect 25421 47073 25455 47107
rect 34345 47073 34379 47107
rect 43361 47073 43395 47107
rect 45569 47073 45603 47107
rect 45937 47073 45971 47107
rect 46949 47073 46983 47107
rect 47133 47073 47167 47107
rect 49433 47073 49467 47107
rect 50813 47073 50847 47107
rect 50905 47073 50939 47107
rect 52193 47073 52227 47107
rect 56701 47073 56735 47107
rect 56793 47073 56827 47107
rect 61209 47073 61243 47107
rect 4261 47005 4295 47039
rect 5641 47005 5675 47039
rect 12265 47005 12299 47039
rect 13921 47005 13955 47039
rect 17141 47005 17175 47039
rect 17417 47005 17451 47039
rect 32597 47005 32631 47039
rect 32873 47005 32907 47039
rect 38945 47005 38979 47039
rect 39221 47005 39255 47039
rect 44925 47005 44959 47039
rect 45477 47005 45511 47039
rect 46029 47005 46063 47039
rect 46305 47005 46339 47039
rect 47501 47005 47535 47039
rect 51365 47005 51399 47039
rect 57253 47005 57287 47039
rect 61485 47005 61519 47039
rect 6101 46937 6135 46971
rect 12081 46937 12115 46971
rect 13369 46937 13403 46971
rect 13829 46937 13863 46971
rect 14197 46937 14231 46971
rect 24225 46937 24259 46971
rect 25513 46937 25547 46971
rect 38761 46937 38795 46971
rect 50629 46937 50663 46971
rect 51457 46937 51491 46971
rect 56517 46937 56551 46971
rect 57345 46937 57379 46971
rect 16957 46869 16991 46903
rect 18705 46869 18739 46903
rect 23857 46869 23891 46903
rect 33977 46869 34011 46903
rect 40325 46869 40359 46903
rect 43453 46869 43487 46903
rect 46489 46869 46523 46903
rect 47593 46869 47627 46903
rect 49525 46869 49559 46903
rect 52377 46869 52411 46903
rect 62589 46869 62623 46903
rect 62957 46869 62991 46903
rect 2513 46665 2547 46699
rect 25329 46665 25363 46699
rect 37289 46665 37323 46699
rect 37473 46665 37507 46699
rect 40601 46665 40635 46699
rect 47593 46665 47627 46699
rect 48789 46665 48823 46699
rect 54953 46665 54987 46699
rect 62129 46665 62163 46699
rect 19993 46597 20027 46631
rect 2881 46529 2915 46563
rect 7573 46529 7607 46563
rect 9137 46529 9171 46563
rect 12449 46529 12483 46563
rect 12725 46529 12759 46563
rect 20085 46529 20119 46563
rect 20821 46529 20855 46563
rect 31125 46529 31159 46563
rect 37657 46529 37691 46563
rect 42533 46529 42567 46563
rect 46673 46529 46707 46563
rect 50537 46529 50571 46563
rect 52009 46529 52043 46563
rect 56425 46529 56459 46563
rect 57621 46529 57655 46563
rect 2605 46461 2639 46495
rect 7297 46461 7331 46495
rect 14197 46461 14231 46495
rect 18061 46461 18095 46495
rect 19073 46461 19107 46495
rect 20729 46461 20763 46495
rect 21097 46461 21131 46495
rect 21281 46461 21315 46495
rect 21465 46461 21499 46495
rect 23949 46461 23983 46495
rect 24225 46461 24259 46495
rect 26433 46461 26467 46495
rect 26709 46461 26743 46495
rect 31309 46461 31343 46495
rect 31861 46461 31895 46495
rect 32045 46461 32079 46495
rect 33793 46461 33827 46495
rect 34897 46461 34931 46495
rect 37841 46461 37875 46495
rect 38301 46461 38335 46495
rect 38393 46461 38427 46495
rect 40509 46461 40543 46495
rect 42257 46461 42291 46495
rect 46305 46461 46339 46495
rect 46765 46461 46799 46495
rect 47501 46461 47535 46495
rect 48513 46461 48547 46495
rect 48697 46461 48731 46495
rect 50169 46461 50203 46495
rect 51733 46461 51767 46495
rect 54861 46461 54895 46495
rect 55873 46461 55907 46495
rect 56057 46461 56091 46495
rect 57345 46461 57379 46495
rect 61761 46461 61795 46495
rect 32689 46393 32723 46427
rect 38945 46393 38979 46427
rect 42073 46393 42107 46427
rect 43913 46393 43947 46427
rect 46121 46393 46155 46427
rect 49985 46393 50019 46427
rect 4169 46325 4203 46359
rect 4445 46325 4479 46359
rect 8677 46325 8711 46359
rect 14013 46325 14047 46359
rect 18153 46325 18187 46359
rect 19165 46325 19199 46359
rect 23765 46325 23799 46359
rect 26249 46325 26283 46359
rect 27813 46325 27847 46359
rect 30941 46325 30975 46359
rect 32321 46325 32355 46359
rect 33885 46325 33919 46359
rect 34989 46325 35023 46359
rect 39221 46325 39255 46359
rect 39405 46325 39439 46359
rect 51457 46325 51491 46359
rect 53113 46325 53147 46359
rect 56609 46325 56643 46359
rect 58725 46325 58759 46359
rect 59185 46325 59219 46359
rect 61853 46325 61887 46359
rect 8033 46121 8067 46155
rect 14013 46121 14047 46155
rect 18613 46121 18647 46155
rect 18797 46121 18831 46155
rect 24961 46121 24995 46155
rect 31953 46121 31987 46155
rect 34437 46121 34471 46155
rect 39221 46121 39255 46155
rect 39405 46121 39439 46155
rect 46857 46121 46891 46155
rect 29469 46053 29503 46087
rect 8033 45985 8067 46019
rect 8401 45985 8435 46019
rect 13921 45985 13955 46019
rect 17049 45985 17083 46019
rect 17601 45985 17635 46019
rect 17785 45985 17819 46019
rect 18337 45985 18371 46019
rect 20637 45985 20671 46019
rect 21557 45985 21591 46019
rect 21925 45985 21959 46019
rect 22109 45985 22143 46019
rect 23949 45985 23983 46019
rect 24501 45985 24535 46019
rect 24685 45985 24719 46019
rect 27077 45985 27111 46019
rect 28733 45985 28767 46019
rect 29101 45985 29135 46019
rect 29285 45985 29319 46019
rect 16957 45917 16991 45951
rect 18061 45917 18095 45951
rect 21373 45917 21407 45951
rect 23765 45917 23799 45951
rect 28089 45917 28123 45951
rect 28825 45917 28859 45951
rect 16773 45849 16807 45883
rect 23581 45849 23615 45883
rect 37289 46053 37323 46087
rect 37473 46053 37507 46087
rect 39037 46053 39071 46087
rect 44373 46053 44407 46087
rect 45661 46053 45695 46087
rect 55689 46053 55723 46087
rect 56241 46053 56275 46087
rect 61761 46053 61795 46087
rect 33149 45985 33183 46019
rect 37749 45985 37783 46019
rect 37933 45985 37967 46019
rect 38485 45985 38519 46019
rect 38669 45985 38703 46019
rect 45017 45985 45051 46019
rect 45385 45985 45419 46019
rect 45569 45985 45603 46019
rect 46397 45985 46431 46019
rect 46673 45985 46707 46019
rect 51181 45985 51215 46019
rect 51733 45985 51767 46019
rect 51917 45985 51951 46019
rect 55873 45985 55907 46019
rect 62589 45985 62623 46019
rect 32873 45917 32907 45951
rect 34621 45917 34655 45951
rect 45109 45917 45143 45951
rect 46489 45917 46523 45951
rect 50997 45917 51031 45951
rect 62313 45917 62347 45951
rect 62773 45917 62807 45951
rect 50629 45849 50663 45883
rect 50813 45849 50847 45883
rect 21189 45781 21223 45815
rect 22293 45781 22327 45815
rect 25329 45781 25363 45815
rect 27169 45781 27203 45815
rect 29653 45781 29687 45815
rect 31953 45781 31987 45815
rect 45937 45781 45971 45815
rect 47317 45781 47351 45815
rect 52193 45781 52227 45815
rect 46213 45577 46247 45611
rect 15025 45509 15059 45543
rect 2881 45441 2915 45475
rect 13461 45441 13495 45475
rect 15209 45441 15243 45475
rect 31033 45441 31067 45475
rect 32321 45441 32355 45475
rect 2605 45373 2639 45407
rect 13737 45373 13771 45407
rect 30665 45373 30699 45407
rect 31217 45373 31251 45407
rect 31769 45373 31803 45407
rect 31953 45373 31987 45407
rect 44465 45373 44499 45407
rect 46121 45373 46155 45407
rect 51917 45373 51951 45407
rect 52009 45373 52043 45407
rect 52377 45373 52411 45407
rect 52469 45373 52503 45407
rect 56057 45373 56091 45407
rect 58081 45373 58115 45407
rect 51365 45305 51399 45339
rect 51549 45305 51583 45339
rect 53021 45305 53055 45339
rect 3985 45237 4019 45271
rect 4445 45237 4479 45271
rect 30849 45237 30883 45271
rect 32597 45237 32631 45271
rect 44557 45237 44591 45271
rect 56149 45237 56183 45271
rect 56425 45237 56459 45271
rect 58173 45237 58207 45271
rect 7205 45033 7239 45067
rect 24409 45033 24443 45067
rect 29193 45033 29227 45067
rect 44557 45033 44591 45067
rect 44741 45033 44775 45067
rect 62497 45033 62531 45067
rect 46121 44965 46155 44999
rect 52285 44965 52319 44999
rect 60197 44965 60231 44999
rect 63601 44965 63635 44999
rect 5365 44897 5399 44931
rect 24225 44897 24259 44931
rect 29009 44897 29043 44931
rect 29377 44897 29411 44931
rect 44833 44897 44867 44931
rect 45002 44897 45036 44931
rect 45477 44897 45511 44931
rect 45569 44897 45603 44931
rect 57713 44897 57747 44931
rect 60381 44897 60415 44931
rect 61761 44897 61795 44931
rect 62589 44897 62623 44931
rect 62957 44897 62991 44931
rect 5641 44829 5675 44863
rect 38945 44829 38979 44863
rect 39221 44829 39255 44863
rect 46397 44829 46431 44863
rect 52653 44829 52687 44863
rect 57437 44829 57471 44863
rect 63233 44829 63267 44863
rect 66637 44829 66671 44863
rect 66729 44829 66763 44863
rect 67005 44829 67039 44863
rect 59277 44761 59311 44795
rect 61577 44761 61611 44795
rect 6929 44693 6963 44727
rect 24041 44693 24075 44727
rect 38761 44693 38795 44727
rect 40509 44693 40543 44727
rect 52450 44693 52484 44727
rect 52561 44693 52595 44727
rect 52929 44693 52963 44727
rect 59001 44693 59035 44727
rect 60473 44693 60507 44727
rect 68293 44693 68327 44727
rect 4445 44489 4479 44523
rect 27445 44489 27479 44523
rect 33701 44489 33735 44523
rect 41521 44489 41555 44523
rect 58541 44489 58575 44523
rect 60611 44489 60645 44523
rect 60749 44489 60783 44523
rect 60933 44489 60967 44523
rect 65257 44489 65291 44523
rect 65993 44489 66027 44523
rect 15301 44421 15335 44455
rect 15485 44421 15519 44455
rect 32321 44421 32355 44455
rect 45753 44421 45787 44455
rect 47685 44421 47719 44455
rect 59829 44421 59863 44455
rect 27905 44353 27939 44387
rect 28733 44353 28767 44387
rect 32505 44353 32539 44387
rect 34069 44353 34103 44387
rect 46121 44353 46155 44387
rect 51733 44353 51767 44387
rect 59001 44353 59035 44387
rect 60841 44353 60875 44387
rect 2605 44285 2639 44319
rect 2881 44285 2915 44319
rect 7665 44285 7699 44319
rect 7941 44285 7975 44319
rect 13737 44285 13771 44319
rect 14013 44285 14047 44319
rect 18705 44285 18739 44319
rect 18981 44285 19015 44319
rect 27813 44285 27847 44319
rect 28181 44285 28215 44319
rect 28365 44285 28399 44319
rect 32689 44285 32723 44319
rect 33241 44285 33275 44319
rect 33425 44285 33459 44319
rect 41429 44285 41463 44319
rect 45937 44285 45971 44319
rect 46305 44285 46339 44319
rect 46765 44285 46799 44319
rect 46857 44285 46891 44319
rect 51917 44285 51951 44319
rect 52377 44285 52411 44319
rect 52469 44285 52503 44319
rect 59093 44285 59127 44319
rect 59461 44285 59495 44319
rect 59645 44285 59679 44319
rect 65073 44285 65107 44319
rect 65441 44285 65475 44319
rect 66177 44285 66211 44319
rect 66729 44285 66763 44319
rect 67005 44285 67039 44319
rect 68569 44285 68603 44319
rect 71421 44285 71455 44319
rect 71697 44285 71731 44319
rect 9321 44217 9355 44251
rect 20361 44217 20395 44251
rect 28549 44217 28583 44251
rect 47409 44217 47443 44251
rect 53021 44217 53055 44251
rect 60473 44217 60507 44251
rect 67373 44217 67407 44251
rect 73169 44217 73203 44251
rect 3985 44149 4019 44183
rect 9413 44149 9447 44183
rect 20545 44149 20579 44183
rect 45569 44149 45603 44183
rect 45937 44149 45971 44183
rect 53297 44149 53331 44183
rect 66269 44149 66303 44183
rect 68661 44149 68695 44183
rect 72985 44149 73019 44183
rect 6929 43945 6963 43979
rect 7757 43945 7791 43979
rect 14013 43945 14047 43979
rect 15669 43945 15703 43979
rect 27353 43945 27387 43979
rect 31953 43945 31987 43979
rect 38577 43945 38611 43979
rect 46581 43945 46615 43979
rect 55229 43945 55263 43979
rect 59001 43945 59035 43979
rect 72893 43945 72927 43979
rect 77401 43945 77435 43979
rect 15393 43877 15427 43911
rect 33517 43877 33551 43911
rect 52377 43877 52411 43911
rect 54585 43877 54619 43911
rect 59185 43877 59219 43911
rect 65993 43877 66027 43911
rect 66177 43877 66211 43911
rect 71421 43877 71455 43911
rect 7021 43809 7055 43843
rect 7389 43809 7423 43843
rect 9689 43809 9723 43843
rect 13001 43809 13035 43843
rect 13553 43809 13587 43843
rect 13737 43809 13771 43843
rect 15301 43809 15335 43843
rect 17233 43809 17267 43843
rect 20913 43809 20947 43843
rect 27905 43809 27939 43843
rect 28273 43809 28307 43843
rect 28457 43809 28491 43843
rect 32229 43809 32263 43843
rect 32413 43809 32447 43843
rect 32965 43809 32999 43843
rect 33149 43809 33183 43843
rect 37013 43809 37047 43843
rect 38485 43809 38519 43843
rect 39957 43809 39991 43843
rect 41337 43809 41371 43843
rect 42165 43809 42199 43843
rect 44741 43809 44775 43843
rect 45293 43809 45327 43843
rect 45845 43809 45879 43843
rect 46029 43809 46063 43843
rect 51089 43809 51123 43843
rect 51273 43809 51307 43843
rect 51825 43809 51859 43843
rect 52009 43809 52043 43843
rect 54732 43809 54766 43843
rect 58909 43809 58943 43843
rect 60197 43809 60231 43843
rect 60381 43809 60415 43843
rect 61577 43809 61611 43843
rect 61761 43809 61795 43843
rect 66729 43809 66763 43843
rect 67005 43809 67039 43843
rect 71605 43809 71639 43843
rect 72801 43809 72835 43843
rect 77585 43809 77619 43843
rect 12817 43741 12851 43775
rect 17693 43741 17727 43775
rect 21925 43741 21959 43775
rect 22201 43741 22235 43775
rect 27997 43741 28031 43775
rect 39681 43741 39715 43775
rect 45109 43741 45143 43775
rect 54953 43741 54987 43775
rect 67189 43741 67223 43775
rect 71881 43741 71915 43775
rect 77861 43741 77895 43775
rect 12725 43673 12759 43707
rect 33793 43673 33827 43707
rect 46305 43673 46339 43707
rect 52653 43673 52687 43707
rect 9781 43605 9815 43639
rect 17417 43605 17451 43639
rect 21005 43605 21039 43639
rect 21833 43605 21867 43639
rect 23489 43605 23523 43639
rect 28641 43605 28675 43639
rect 28825 43605 28859 43639
rect 36829 43605 36863 43639
rect 39497 43605 39531 43639
rect 42257 43605 42291 43639
rect 44925 43605 44959 43639
rect 46765 43605 46799 43639
rect 54861 43605 54895 43639
rect 60473 43605 60507 43639
rect 61853 43605 61887 43639
rect 79149 43605 79183 43639
rect 3985 43401 4019 43435
rect 4445 43401 4479 43435
rect 12725 43401 12759 43435
rect 14013 43401 14047 43435
rect 15301 43401 15335 43435
rect 21465 43401 21499 43435
rect 22661 43401 22695 43435
rect 25789 43401 25823 43435
rect 37013 43401 37047 43435
rect 52929 43401 52963 43435
rect 53481 43401 53515 43435
rect 60289 43401 60323 43435
rect 4629 43333 4663 43367
rect 8953 43333 8987 43367
rect 19165 43333 19199 43367
rect 19625 43333 19659 43367
rect 24777 43333 24811 43367
rect 37197 43333 37231 43367
rect 37749 43333 37783 43367
rect 72985 43333 73019 43367
rect 2881 43265 2915 43299
rect 12817 43265 12851 43299
rect 35449 43265 35483 43299
rect 53297 43265 53331 43299
rect 71605 43265 71639 43299
rect 77585 43265 77619 43299
rect 2605 43197 2639 43231
rect 7849 43197 7883 43231
rect 8033 43197 8067 43231
rect 8493 43197 8527 43231
rect 8585 43197 8619 43231
rect 13001 43197 13035 43231
rect 13553 43197 13587 43231
rect 13737 43197 13771 43231
rect 15025 43197 15059 43231
rect 18061 43197 18095 43231
rect 18245 43197 18279 43231
rect 18705 43197 18739 43231
rect 18797 43197 18831 43231
rect 20453 43197 20487 43231
rect 20545 43197 20579 43231
rect 20919 43197 20953 43231
rect 21005 43197 21039 43231
rect 22477 43197 22511 43231
rect 23673 43197 23707 43231
rect 24961 43197 24995 43231
rect 25973 43197 26007 43231
rect 26249 43197 26283 43231
rect 32413 43197 32447 43231
rect 32597 43197 32631 43231
rect 33149 43197 33183 43231
rect 33333 43197 33367 43231
rect 35725 43197 35759 43231
rect 37933 43197 37967 43231
rect 38209 43197 38243 43231
rect 51733 43197 51767 43231
rect 51917 43197 51951 43231
rect 52377 43197 52411 43231
rect 52469 43197 52503 43231
rect 58817 43197 58851 43231
rect 59829 43197 59863 43231
rect 60105 43197 60139 43231
rect 61393 43197 61427 43231
rect 61577 43197 61611 43231
rect 66913 43197 66947 43231
rect 71145 43197 71179 43231
rect 71237 43197 71271 43231
rect 71421 43197 71455 43231
rect 72709 43197 72743 43231
rect 78137 43197 78171 43231
rect 78413 43197 78447 43231
rect 78597 43197 78631 43231
rect 15117 43129 15151 43163
rect 20085 43129 20119 43163
rect 21833 43129 21867 43163
rect 33701 43129 33735 43163
rect 51273 43129 51307 43163
rect 60013 43129 60047 43163
rect 66729 43129 66763 43163
rect 71973 43129 72007 43163
rect 7665 43061 7699 43095
rect 9321 43061 9355 43095
rect 17785 43061 17819 43095
rect 22293 43061 22327 43095
rect 23765 43061 23799 43095
rect 25053 43061 25087 43095
rect 27537 43061 27571 43095
rect 32321 43061 32355 43095
rect 33977 43061 34011 43095
rect 39497 43061 39531 43095
rect 51457 43061 51491 43095
rect 58909 43061 58943 43095
rect 60657 43061 60691 43095
rect 61669 43061 61703 43095
rect 67005 43061 67039 43095
rect 72801 43061 72835 43095
rect 77493 43061 77527 43095
rect 32505 42857 32539 42891
rect 39037 42857 39071 42891
rect 44833 42857 44867 42891
rect 46581 42857 46615 42891
rect 51181 42857 51215 42891
rect 53021 42857 53055 42891
rect 53205 42857 53239 42891
rect 77861 42857 77895 42891
rect 7573 42789 7607 42823
rect 66361 42789 66395 42823
rect 7113 42721 7147 42755
rect 7389 42721 7423 42755
rect 7757 42721 7791 42755
rect 13737 42721 13771 42755
rect 14105 42721 14139 42755
rect 14289 42721 14323 42755
rect 20913 42721 20947 42755
rect 21281 42721 21315 42755
rect 30849 42721 30883 42755
rect 30941 42721 30975 42755
rect 32689 42721 32723 42755
rect 32873 42721 32907 42755
rect 33425 42721 33459 42755
rect 33609 42721 33643 42755
rect 34253 42721 34287 42755
rect 38945 42721 38979 42755
rect 44649 42721 44683 42755
rect 45017 42721 45051 42755
rect 45201 42721 45235 42755
rect 45661 42721 45695 42755
rect 45753 42721 45787 42755
rect 46765 42721 46799 42755
rect 51641 42721 51675 42755
rect 52101 42721 52135 42755
rect 52193 42721 52227 42755
rect 58633 42721 58667 42755
rect 58725 42721 58759 42755
rect 58817 42721 58851 42755
rect 59461 42721 59495 42755
rect 60197 42721 60231 42755
rect 60749 42721 60783 42755
rect 66453 42721 66487 42755
rect 68753 42721 68787 42755
rect 68937 42721 68971 42755
rect 69673 42721 69707 42755
rect 72065 42721 72099 42755
rect 72433 42721 72467 42755
rect 72525 42721 72559 42755
rect 77769 42721 77803 42755
rect 78321 42721 78355 42755
rect 79701 42721 79735 42755
rect 13093 42653 13127 42687
rect 13645 42653 13679 42687
rect 33977 42653 34011 42687
rect 51457 42653 51491 42687
rect 69305 42653 69339 42687
rect 71973 42653 72007 42687
rect 72709 42653 72743 42687
rect 77401 42653 77435 42687
rect 78597 42653 78631 42687
rect 46213 42585 46247 42619
rect 51365 42585 51399 42619
rect 52561 42585 52595 42619
rect 60289 42585 60323 42619
rect 66177 42585 66211 42619
rect 69075 42585 69109 42619
rect 71513 42585 71547 42619
rect 21097 42517 21131 42551
rect 31125 42517 31159 42551
rect 59001 42517 59035 42551
rect 66637 42517 66671 42551
rect 67005 42517 67039 42551
rect 69213 42517 69247 42551
rect 77585 42517 77619 42551
rect 79793 42517 79827 42551
rect 3985 42313 4019 42347
rect 4629 42313 4663 42347
rect 7665 42313 7699 42347
rect 16221 42313 16255 42347
rect 19625 42313 19659 42347
rect 25421 42313 25455 42347
rect 27261 42313 27295 42347
rect 51365 42313 51399 42347
rect 51549 42313 51583 42347
rect 53205 42313 53239 42347
rect 60933 42313 60967 42347
rect 64337 42313 64371 42347
rect 67005 42313 67039 42347
rect 70777 42313 70811 42347
rect 78045 42313 78079 42347
rect 15945 42245 15979 42279
rect 19809 42245 19843 42279
rect 31309 42245 31343 42279
rect 60013 42245 60047 42279
rect 2605 42177 2639 42211
rect 18981 42177 19015 42211
rect 45569 42177 45603 42211
rect 46121 42177 46155 42211
rect 51549 42177 51583 42211
rect 51733 42177 51767 42211
rect 58449 42177 58483 42211
rect 64429 42177 64463 42211
rect 64705 42177 64739 42211
rect 69121 42177 69155 42211
rect 72433 42177 72467 42211
rect 77585 42177 77619 42211
rect 78413 42177 78447 42211
rect 2881 42109 2915 42143
rect 4353 42109 4387 42143
rect 7481 42109 7515 42143
rect 15761 42109 15795 42143
rect 18889 42109 18923 42143
rect 19257 42109 19291 42143
rect 19441 42109 19475 42143
rect 24225 42109 24259 42143
rect 24409 42109 24443 42143
rect 24961 42109 24995 42143
rect 25145 42109 25179 42143
rect 26893 42109 26927 42143
rect 31125 42109 31159 42143
rect 46305 42109 46339 42143
rect 46765 42109 46799 42143
rect 46857 42109 46891 42143
rect 51917 42109 51951 42143
rect 52377 42109 52411 42143
rect 52469 42109 52503 42143
rect 58173 42109 58207 42143
rect 60841 42109 60875 42143
rect 67189 42109 67223 42143
rect 67465 42109 67499 42143
rect 68845 42109 68879 42143
rect 70693 42109 70727 42143
rect 72065 42109 72099 42143
rect 72617 42109 72651 42143
rect 77861 42109 77895 42143
rect 18245 42041 18279 42075
rect 47409 42041 47443 42075
rect 53021 42041 53055 42075
rect 60657 42041 60691 42075
rect 68661 42041 68695 42075
rect 71881 42041 71915 42075
rect 77769 42041 77803 42075
rect 24041 41973 24075 42007
rect 26985 41973 27019 42007
rect 30941 41973 30975 42007
rect 45845 41973 45879 42007
rect 47685 41973 47719 42007
rect 51181 41973 51215 42007
rect 59737 41973 59771 42007
rect 65993 41973 66027 42007
rect 6009 41769 6043 41803
rect 12909 41769 12943 41803
rect 16129 41769 16163 41803
rect 16405 41769 16439 41803
rect 27261 41769 27295 41803
rect 29653 41769 29687 41803
rect 29929 41769 29963 41803
rect 34713 41769 34747 41803
rect 53481 41769 53515 41803
rect 60289 41769 60323 41803
rect 34989 41701 35023 41735
rect 39129 41701 39163 41735
rect 66637 41701 66671 41735
rect 77401 41701 77435 41735
rect 6193 41633 6227 41667
rect 6469 41633 6503 41667
rect 7481 41633 7515 41667
rect 11069 41633 11103 41667
rect 15945 41633 15979 41667
rect 26525 41633 26559 41667
rect 26617 41633 26651 41667
rect 27905 41633 27939 41667
rect 29469 41633 29503 41667
rect 33425 41633 33459 41667
rect 39497 41633 39531 41667
rect 40049 41633 40083 41667
rect 40233 41633 40267 41667
rect 45661 41633 45695 41667
rect 45845 41633 45879 41667
rect 46029 41633 46063 41667
rect 46581 41633 46615 41667
rect 46765 41633 46799 41667
rect 47409 41633 47443 41667
rect 52193 41633 52227 41667
rect 52653 41633 52687 41667
rect 52745 41633 52779 41667
rect 60197 41633 60231 41667
rect 60473 41633 60507 41667
rect 66821 41633 66855 41667
rect 72341 41633 72375 41667
rect 72525 41633 72559 41667
rect 75837 41633 75871 41667
rect 77585 41633 77619 41667
rect 77861 41633 77895 41667
rect 11345 41565 11379 41599
rect 33149 41565 33183 41599
rect 39313 41565 39347 41599
rect 47133 41565 47167 41599
rect 52009 41565 52043 41599
rect 53297 41565 53331 41599
rect 76205 41565 76239 41599
rect 83197 41565 83231 41599
rect 83381 41565 83415 41599
rect 83657 41565 83691 41599
rect 7665 41497 7699 41531
rect 27813 41497 27847 41531
rect 51641 41497 51675 41531
rect 76021 41497 76055 41531
rect 12449 41429 12483 41463
rect 26801 41429 26835 41463
rect 27997 41429 28031 41463
rect 40509 41429 40543 41463
rect 40877 41429 40911 41463
rect 45477 41429 45511 41463
rect 51825 41429 51859 41463
rect 66913 41429 66947 41463
rect 72617 41429 72651 41463
rect 78965 41429 78999 41463
rect 84761 41429 84795 41463
rect 11345 41225 11379 41259
rect 27721 41225 27755 41259
rect 29377 41225 29411 41259
rect 39957 41225 39991 41259
rect 40049 41225 40083 41259
rect 40233 41225 40267 41259
rect 42073 41225 42107 41259
rect 53389 41225 53423 41259
rect 72801 41225 72835 41259
rect 4445 41157 4479 41191
rect 12449 41157 12483 41191
rect 3985 41089 4019 41123
rect 11713 41089 11747 41123
rect 18705 41089 18739 41123
rect 19441 41089 19475 41123
rect 23949 41089 23983 41123
rect 25237 41089 25271 41123
rect 26433 41089 26467 41123
rect 29377 41089 29411 41123
rect 29745 41089 29779 41123
rect 39497 41089 39531 41123
rect 2612 41021 2646 41055
rect 2881 41021 2915 41055
rect 5457 41021 5491 41055
rect 5733 41021 5767 41055
rect 6837 41021 6871 41055
rect 7389 41021 7423 41055
rect 9873 41021 9907 41055
rect 10149 41021 10183 41055
rect 10333 41021 10367 41055
rect 10793 41021 10827 41055
rect 10885 41021 10919 41055
rect 12449 41021 12483 41055
rect 12725 41021 12759 41055
rect 13461 41021 13495 41055
rect 13645 41021 13679 41055
rect 14013 41021 14047 41055
rect 14197 41021 14231 41055
rect 19349 41021 19383 41055
rect 19717 41021 19751 41055
rect 19901 41021 19935 41055
rect 24133 41021 24167 41055
rect 24685 41021 24719 41055
rect 24869 41021 24903 41055
rect 26157 41021 26191 41055
rect 29837 41021 29871 41055
rect 30389 41021 30423 41055
rect 30573 41021 30607 41055
rect 31217 41021 31251 41055
rect 38209 41021 38243 41055
rect 38393 41021 38427 41055
rect 38853 41021 38887 41055
rect 39033 41021 39067 41055
rect 46857 41157 46891 41191
rect 60841 41157 60875 41191
rect 61117 41157 61151 41191
rect 65441 41157 65475 41191
rect 72249 41157 72283 41191
rect 83197 41157 83231 41191
rect 41705 41089 41739 41123
rect 47225 41089 47259 41123
rect 48513 41089 48547 41123
rect 53260 41089 53294 41123
rect 53481 41089 53515 41123
rect 59277 41089 59311 41123
rect 59553 41089 59587 41123
rect 66361 41089 66395 41123
rect 72120 41089 72154 41123
rect 72709 41089 72743 41123
rect 76297 41089 76331 41123
rect 77585 41089 77619 41123
rect 40509 41021 40543 41055
rect 40693 41021 40727 41055
rect 41153 41021 41187 41055
rect 41245 41021 41279 41055
rect 47041 41021 47075 41055
rect 47409 41021 47443 41055
rect 47869 41021 47903 41055
rect 47961 41021 47995 41055
rect 53113 41021 53147 41055
rect 58817 41021 58851 41055
rect 59069 41021 59103 41055
rect 65349 41021 65383 41055
rect 65625 41021 65659 41055
rect 66637 41021 66671 41055
rect 71973 41021 72007 41055
rect 72312 41021 72346 41055
rect 76205 41021 76239 41055
rect 76481 41021 76515 41055
rect 77217 41021 77251 41055
rect 77769 41021 77803 41055
rect 83013 41021 83047 41055
rect 12909 40953 12943 40987
rect 30941 40953 30975 40987
rect 40049 40953 40083 40987
rect 48881 40953 48915 40987
rect 66545 40953 66579 40987
rect 67097 40953 67131 40987
rect 83381 40953 83415 40987
rect 5273 40885 5307 40919
rect 6929 40885 6963 40919
rect 9873 40885 9907 40919
rect 9965 40885 9999 40919
rect 13093 40885 13127 40919
rect 23765 40885 23799 40919
rect 27905 40885 27939 40919
rect 29469 40885 29503 40919
rect 38025 40885 38059 40919
rect 39773 40885 39807 40919
rect 48697 40885 48731 40919
rect 53757 40885 53791 40919
rect 58909 40885 58943 40919
rect 67281 40885 67315 40919
rect 71789 40885 71823 40919
rect 7297 40681 7331 40715
rect 12633 40681 12667 40715
rect 27261 40681 27295 40715
rect 58449 40681 58483 40715
rect 77677 40681 77711 40715
rect 84669 40681 84703 40715
rect 15577 40613 15611 40647
rect 20361 40613 20395 40647
rect 27077 40613 27111 40647
rect 40233 40613 40267 40647
rect 40417 40613 40451 40647
rect 40877 40613 40911 40647
rect 58725 40613 58759 40647
rect 60289 40613 60323 40647
rect 82737 40613 82771 40647
rect 5733 40545 5767 40579
rect 6009 40545 6043 40579
rect 7021 40545 7055 40579
rect 7573 40545 7607 40579
rect 9505 40545 9539 40579
rect 10241 40545 10275 40579
rect 12541 40545 12575 40579
rect 15761 40545 15795 40579
rect 18797 40545 18831 40579
rect 19441 40545 19475 40579
rect 19809 40545 19843 40579
rect 19993 40545 20027 40579
rect 20177 40545 20211 40579
rect 26617 40545 26651 40579
rect 29561 40545 29595 40579
rect 30021 40545 30055 40579
rect 30113 40545 30147 40579
rect 38853 40545 38887 40579
rect 39405 40545 39439 40579
rect 39589 40545 39623 40579
rect 44373 40545 44407 40579
rect 44741 40545 44775 40579
rect 45201 40545 45235 40579
rect 45293 40545 45327 40579
rect 52653 40545 52687 40579
rect 58633 40545 58667 40579
rect 60197 40545 60231 40579
rect 66085 40545 66119 40579
rect 77401 40545 77435 40579
rect 77585 40545 77619 40579
rect 83565 40545 83599 40579
rect 83749 40545 83783 40579
rect 83841 40545 83875 40579
rect 84577 40545 84611 40579
rect 5917 40477 5951 40511
rect 16037 40477 16071 40511
rect 17417 40477 17451 40511
rect 19349 40477 19383 40511
rect 22109 40477 22143 40511
rect 22385 40477 22419 40511
rect 26525 40477 26559 40511
rect 29377 40477 29411 40511
rect 30665 40477 30699 40511
rect 33149 40477 33183 40511
rect 33425 40477 33459 40511
rect 38577 40477 38611 40511
rect 38669 40477 38703 40511
rect 39957 40477 39991 40511
rect 41245 40477 41279 40511
rect 44557 40477 44591 40511
rect 46305 40477 46339 40511
rect 53021 40477 53055 40511
rect 65625 40477 65659 40511
rect 65809 40477 65843 40511
rect 67189 40477 67223 40511
rect 71973 40477 72007 40511
rect 72157 40477 72191 40511
rect 72433 40477 72467 40511
rect 83289 40477 83323 40511
rect 9505 40409 9539 40443
rect 30849 40409 30883 40443
rect 41153 40409 41187 40443
rect 52929 40409 52963 40443
rect 10333 40341 10367 40375
rect 21925 40341 21959 40375
rect 23673 40341 23707 40375
rect 29193 40341 29227 40375
rect 32965 40341 32999 40375
rect 34713 40341 34747 40375
rect 41015 40341 41049 40375
rect 41521 40341 41555 40375
rect 45753 40341 45787 40375
rect 46029 40341 46063 40375
rect 46489 40341 46523 40375
rect 52818 40341 52852 40375
rect 53297 40341 53331 40375
rect 73537 40341 73571 40375
rect 10149 40137 10183 40171
rect 29469 40137 29503 40171
rect 57805 40137 57839 40171
rect 58817 40137 58851 40171
rect 72709 40137 72743 40171
rect 74273 40137 74307 40171
rect 83749 40137 83783 40171
rect 40785 40069 40819 40103
rect 48697 40069 48731 40103
rect 54106 40069 54140 40103
rect 54861 40069 54895 40103
rect 82737 40069 82771 40103
rect 16129 40001 16163 40035
rect 18429 40001 18463 40035
rect 40656 40001 40690 40035
rect 40877 40001 40911 40035
rect 48513 40001 48547 40035
rect 54309 40001 54343 40035
rect 58633 40001 58667 40035
rect 83381 40001 83415 40035
rect 8769 39933 8803 39967
rect 9045 39933 9079 39967
rect 15669 39933 15703 39967
rect 16865 39933 16899 39967
rect 18061 39933 18095 39967
rect 23673 39933 23707 39967
rect 29285 39933 29319 39967
rect 47225 39933 47259 39967
rect 47409 39933 47443 39967
rect 47869 39933 47903 39967
rect 47961 39933 47995 39967
rect 53941 39933 53975 39967
rect 54171 39933 54205 39967
rect 57989 39933 58023 39967
rect 58081 39933 58115 39967
rect 59001 39933 59035 39967
rect 59185 39933 59219 39967
rect 59645 39933 59679 39967
rect 59737 39933 59771 39967
rect 71237 39933 71271 39967
rect 72341 39933 72375 39967
rect 72525 39933 72559 39967
rect 74181 39933 74215 39967
rect 77401 39933 77435 39967
rect 82461 39933 82495 39967
rect 83197 39933 83231 39967
rect 18153 39865 18187 39899
rect 23765 39865 23799 39899
rect 40509 39865 40543 39899
rect 47041 39865 47075 39899
rect 48881 39865 48915 39899
rect 60289 39865 60323 39899
rect 72433 39865 72467 39899
rect 10609 39797 10643 39831
rect 15853 39797 15887 39831
rect 17049 39797 17083 39831
rect 17325 39797 17359 39831
rect 29745 39797 29779 39831
rect 41153 39797 41187 39831
rect 46857 39797 46891 39831
rect 54585 39797 54619 39831
rect 60565 39797 60599 39831
rect 71329 39797 71363 39831
rect 73169 39797 73203 39831
rect 77585 39797 77619 39831
rect 82369 39797 82403 39831
rect 22385 39593 22419 39627
rect 22753 39593 22787 39627
rect 45477 39593 45511 39627
rect 45845 39593 45879 39627
rect 48237 39593 48271 39627
rect 59921 39593 59955 39627
rect 72249 39593 72283 39627
rect 73261 39593 73295 39627
rect 77769 39593 77803 39627
rect 84025 39593 84059 39627
rect 32873 39525 32907 39559
rect 46305 39525 46339 39559
rect 48421 39525 48455 39559
rect 54585 39525 54619 39559
rect 65993 39525 66027 39559
rect 71605 39525 71639 39559
rect 72985 39525 73019 39559
rect 78137 39525 78171 39559
rect 4537 39457 4571 39491
rect 16129 39457 16163 39491
rect 17969 39457 18003 39491
rect 21373 39457 21407 39491
rect 21833 39457 21867 39491
rect 21925 39457 21959 39491
rect 27997 39457 28031 39491
rect 29745 39457 29779 39491
rect 33057 39457 33091 39491
rect 39037 39457 39071 39491
rect 39497 39457 39531 39491
rect 39589 39457 39623 39491
rect 40325 39457 40359 39491
rect 44189 39457 44223 39491
rect 44465 39457 44499 39491
rect 44925 39457 44959 39491
rect 45017 39457 45051 39491
rect 46489 39457 46523 39491
rect 46673 39457 46707 39491
rect 47225 39457 47259 39491
rect 47409 39457 47443 39491
rect 52285 39457 52319 39491
rect 52745 39457 52779 39491
rect 52837 39457 52871 39491
rect 60841 39457 60875 39491
rect 61209 39457 61243 39491
rect 61393 39457 61427 39491
rect 65901 39457 65935 39491
rect 67005 39457 67039 39491
rect 67097 39457 67131 39491
rect 71789 39457 71823 39491
rect 72157 39457 72191 39491
rect 73169 39457 73203 39491
rect 77953 39457 77987 39491
rect 78229 39457 78263 39491
rect 84209 39457 84243 39491
rect 16405 39389 16439 39423
rect 17785 39389 17819 39423
rect 21189 39389 21223 39423
rect 28273 39389 28307 39423
rect 33333 39389 33367 39423
rect 38945 39389 38979 39423
rect 44281 39389 44315 39423
rect 46029 39389 46063 39423
rect 52101 39389 52135 39423
rect 53665 39389 53699 39423
rect 53849 39389 53883 39423
rect 54950 39389 54984 39423
rect 60933 39389 60967 39423
rect 67373 39389 67407 39423
rect 84485 39389 84519 39423
rect 47685 39321 47719 39355
rect 54723 39321 54757 39355
rect 72801 39321 72835 39355
rect 4629 39253 4663 39287
rect 21005 39253 21039 39287
rect 29561 39253 29595 39287
rect 34621 39253 34655 39287
rect 40049 39253 40083 39287
rect 40601 39253 40635 39287
rect 44005 39253 44039 39287
rect 47961 39253 47995 39287
rect 51733 39253 51767 39287
rect 51917 39253 51951 39287
rect 53297 39253 53331 39287
rect 54861 39253 54895 39287
rect 55229 39253 55263 39287
rect 60289 39253 60323 39287
rect 68477 39253 68511 39287
rect 71421 39253 71455 39287
rect 78413 39253 78447 39287
rect 85589 39253 85623 39287
rect 4537 39049 4571 39083
rect 4813 39049 4847 39083
rect 9873 39049 9907 39083
rect 13829 39049 13863 39083
rect 14657 39049 14691 39083
rect 23765 39049 23799 39083
rect 28457 39049 28491 39083
rect 54493 39049 54527 39083
rect 54677 39049 54711 39083
rect 72985 39049 73019 39083
rect 78689 39049 78723 39083
rect 84393 39049 84427 39083
rect 86325 39049 86359 39083
rect 9413 38981 9447 39015
rect 2973 38913 3007 38947
rect 16037 38981 16071 39015
rect 28181 38981 28215 39015
rect 46121 38981 46155 39015
rect 54355 38981 54389 39015
rect 58357 38981 58391 39015
rect 60565 38981 60599 39015
rect 62129 38981 62163 39015
rect 68845 38981 68879 39015
rect 77033 38981 77067 39015
rect 46397 38913 46431 38947
rect 48053 38913 48087 38947
rect 48145 38913 48179 38947
rect 54585 38913 54619 38947
rect 58541 38913 58575 38947
rect 59829 38913 59863 38947
rect 61301 38913 61335 38947
rect 64797 38913 64831 38947
rect 72157 38913 72191 38947
rect 72341 38913 72375 38947
rect 77401 38913 77435 38947
rect 80161 38913 80195 38947
rect 87889 38913 87923 38947
rect 3249 38845 3283 38879
rect 8309 38845 8343 38879
rect 8493 38845 8527 38879
rect 8953 38845 8987 38879
rect 9045 38845 9079 38879
rect 14013 38845 14047 38879
rect 14657 38845 14691 38879
rect 14933 38845 14967 38879
rect 15117 38845 15151 38879
rect 15577 38845 15611 38879
rect 15669 38845 15703 38879
rect 23673 38845 23707 38879
rect 27997 38845 28031 38879
rect 36553 38845 36587 38879
rect 36737 38845 36771 38879
rect 46489 38845 46523 38879
rect 47041 38845 47075 38879
rect 47225 38845 47259 38879
rect 52009 38845 52043 38879
rect 52193 38845 52227 38879
rect 52653 38845 52687 38879
rect 52745 38845 52779 38879
rect 53573 38845 53607 38879
rect 53665 38845 53699 38879
rect 54217 38845 54251 38879
rect 58725 38845 58759 38879
rect 59185 38845 59219 38879
rect 59277 38845 59311 38879
rect 61393 38845 61427 38879
rect 61761 38845 61795 38879
rect 61945 38845 61979 38879
rect 64981 38845 65015 38879
rect 65165 38845 65199 38879
rect 65533 38845 65567 38879
rect 65625 38845 65659 38879
rect 66913 38845 66947 38879
rect 67189 38845 67223 38879
rect 68753 38845 68787 38879
rect 71053 38845 71087 38879
rect 71697 38845 71731 38879
rect 71789 38845 71823 38879
rect 72065 38845 72099 38879
rect 73077 38845 73111 38879
rect 77125 38845 77159 38879
rect 79793 38845 79827 38879
rect 83197 38845 83231 38879
rect 83565 38845 83599 38879
rect 84301 38845 84335 38879
rect 85405 38845 85439 38879
rect 86509 38845 86543 38879
rect 86785 38845 86819 38879
rect 47593 38777 47627 38811
rect 51549 38777 51583 38811
rect 51917 38777 51951 38811
rect 60749 38777 60783 38811
rect 64337 38777 64371 38811
rect 85497 38777 85531 38811
rect 8125 38709 8159 38743
rect 14841 38709 14875 38743
rect 36369 38709 36403 38743
rect 47777 38709 47811 38743
rect 53205 38709 53239 38743
rect 58265 38709 58299 38743
rect 60013 38709 60047 38743
rect 65809 38709 65843 38743
rect 67005 38709 67039 38743
rect 70869 38709 70903 38743
rect 72617 38709 72651 38743
rect 73169 38709 73203 38743
rect 79885 38709 79919 38743
rect 83381 38709 83415 38743
rect 28181 38505 28215 38539
rect 40417 38505 40451 38539
rect 53113 38505 53147 38539
rect 72433 38505 72467 38539
rect 76665 38505 76699 38539
rect 79793 38505 79827 38539
rect 84393 38505 84427 38539
rect 17601 38437 17635 38471
rect 17877 38437 17911 38471
rect 21281 38437 21315 38471
rect 23121 38437 23155 38471
rect 27905 38437 27939 38471
rect 64521 38437 64555 38471
rect 79701 38437 79735 38471
rect 83105 38437 83139 38471
rect 10793 38369 10827 38403
rect 12633 38369 12667 38403
rect 15470 38369 15504 38403
rect 16037 38369 16071 38403
rect 16221 38369 16255 38403
rect 17509 38369 17543 38403
rect 21465 38369 21499 38403
rect 26801 38369 26835 38403
rect 27353 38369 27387 38403
rect 27537 38369 27571 38403
rect 38945 38369 38979 38403
rect 39405 38369 39439 38403
rect 39497 38369 39531 38403
rect 40693 38369 40727 38403
rect 40785 38369 40819 38403
rect 40969 38369 41003 38403
rect 52469 38369 52503 38403
rect 52616 38369 52650 38403
rect 60197 38369 60231 38403
rect 60344 38369 60378 38403
rect 64245 38369 64279 38403
rect 64429 38369 64463 38403
rect 65625 38369 65659 38403
rect 72249 38369 72283 38403
rect 73353 38369 73387 38403
rect 76849 38369 76883 38403
rect 77585 38369 77619 38403
rect 77953 38369 77987 38403
rect 78321 38369 78355 38403
rect 78597 38369 78631 38403
rect 78965 38369 78999 38403
rect 80529 38369 80563 38403
rect 80621 38369 80655 38403
rect 83749 38369 83783 38403
rect 84117 38369 84151 38403
rect 11069 38301 11103 38335
rect 15301 38301 15335 38335
rect 21741 38301 21775 38335
rect 26525 38301 26559 38335
rect 26617 38301 26651 38335
rect 33149 38301 33183 38335
rect 33425 38301 33459 38335
rect 38761 38301 38795 38335
rect 16405 38233 16439 38267
rect 34713 38233 34747 38267
rect 39865 38233 39899 38267
rect 41337 38301 41371 38335
rect 52837 38301 52871 38335
rect 60565 38301 60599 38335
rect 77769 38301 77803 38335
rect 79112 38301 79146 38335
rect 79333 38301 79367 38335
rect 83657 38301 83691 38335
rect 84209 38301 84243 38335
rect 52745 38233 52779 38267
rect 59921 38233 59955 38267
rect 60473 38233 60507 38267
rect 65257 38233 65291 38267
rect 73537 38233 73571 38267
rect 79241 38233 79275 38267
rect 82921 38233 82955 38267
rect 12357 38165 12391 38199
rect 15117 38165 15151 38199
rect 16773 38165 16807 38199
rect 26249 38165 26283 38199
rect 26525 38165 26559 38199
rect 32965 38165 32999 38199
rect 40233 38165 40267 38199
rect 40693 38165 40727 38199
rect 41107 38165 41141 38199
rect 41245 38165 41279 38199
rect 41613 38165 41647 38199
rect 60841 38165 60875 38199
rect 65441 38165 65475 38199
rect 78781 38165 78815 38199
rect 4353 37961 4387 37995
rect 4721 37961 4755 37995
rect 4905 37961 4939 37995
rect 5089 37961 5123 37995
rect 10701 37961 10735 37995
rect 22201 37961 22235 37995
rect 23673 37961 23707 37995
rect 52929 37961 52963 37995
rect 58771 37961 58805 37995
rect 58909 37961 58943 37995
rect 72249 37961 72283 37995
rect 77493 37961 77527 37995
rect 77769 37961 77803 37995
rect 86693 37961 86727 37995
rect 16405 37893 16439 37927
rect 21741 37893 21775 37927
rect 3065 37825 3099 37859
rect 3249 37825 3283 37859
rect 11069 37825 11103 37859
rect 12541 37825 12575 37859
rect 3341 37757 3375 37791
rect 3801 37757 3835 37791
rect 3893 37757 3927 37791
rect 5641 37757 5675 37791
rect 9505 37757 9539 37791
rect 9689 37757 9723 37791
rect 10241 37757 10275 37791
rect 10425 37757 10459 37791
rect 12449 37757 12483 37791
rect 16129 37757 16163 37791
rect 16221 37757 16255 37791
rect 20361 37757 20395 37791
rect 20637 37757 20671 37791
rect 20821 37757 20855 37791
rect 21373 37757 21407 37791
rect 21557 37757 21591 37791
rect 5733 37689 5767 37723
rect 38991 37893 39025 37927
rect 39129 37893 39163 37927
rect 58449 37893 58483 37927
rect 81357 37893 81391 37927
rect 25329 37825 25363 37859
rect 25513 37825 25547 37859
rect 39221 37825 39255 37859
rect 53297 37825 53331 37859
rect 58998 37825 59032 37859
rect 65441 37825 65475 37859
rect 23949 37757 23983 37791
rect 25697 37757 25731 37791
rect 26157 37757 26191 37791
rect 26249 37757 26283 37791
rect 33149 37757 33183 37791
rect 33609 37757 33643 37791
rect 34897 37757 34931 37791
rect 46121 37757 46155 37791
rect 51733 37757 51767 37791
rect 51917 37757 51951 37791
rect 52377 37757 52411 37791
rect 52469 37757 52503 37791
rect 53481 37757 53515 37791
rect 61117 37757 61151 37791
rect 63509 37757 63543 37791
rect 64981 37757 65015 37791
rect 65165 37757 65199 37791
rect 65533 37757 65567 37791
rect 72341 37757 72375 37791
rect 74181 37757 74215 37791
rect 77401 37757 77435 37791
rect 79793 37757 79827 37791
rect 79977 37757 80011 37791
rect 80437 37757 80471 37791
rect 81173 37757 81207 37791
rect 86601 37757 86635 37791
rect 23673 37689 23707 37723
rect 23765 37689 23799 37723
rect 26801 37689 26835 37723
rect 38853 37689 38887 37723
rect 39589 37689 39623 37723
rect 58633 37689 58667 37723
rect 63601 37689 63635 37723
rect 64337 37689 64371 37723
rect 80345 37689 80379 37723
rect 9321 37621 9355 37655
rect 16129 37621 16163 37655
rect 16681 37621 16715 37655
rect 20361 37621 20395 37655
rect 20453 37621 20487 37655
rect 24133 37621 24167 37655
rect 26985 37621 27019 37655
rect 32965 37621 32999 37655
rect 33701 37621 33735 37655
rect 34989 37621 35023 37655
rect 46213 37621 46247 37655
rect 59277 37621 59311 37655
rect 60933 37621 60967 37655
rect 63325 37621 63359 37655
rect 64153 37621 64187 37655
rect 64797 37621 64831 37655
rect 72525 37621 72559 37655
rect 74365 37621 74399 37655
rect 5549 37417 5583 37451
rect 10977 37417 11011 37451
rect 11253 37417 11287 37451
rect 63969 37417 64003 37451
rect 66269 37417 66303 37451
rect 72433 37417 72467 37451
rect 73537 37417 73571 37451
rect 78965 37417 78999 37451
rect 86141 37417 86175 37451
rect 5917 37349 5951 37383
rect 20913 37349 20947 37383
rect 22293 37349 22327 37383
rect 28549 37349 28583 37383
rect 33425 37349 33459 37383
rect 33701 37349 33735 37383
rect 38301 37349 38335 37383
rect 46581 37349 46615 37383
rect 53113 37349 53147 37383
rect 53389 37349 53423 37383
rect 53573 37349 53607 37383
rect 60289 37349 60323 37383
rect 79149 37349 79183 37383
rect 79333 37349 79367 37383
rect 80161 37349 80195 37383
rect 80897 37349 80931 37383
rect 85589 37349 85623 37383
rect 4169 37281 4203 37315
rect 9505 37281 9539 37315
rect 10333 37281 10367 37315
rect 10701 37281 10735 37315
rect 10885 37281 10919 37315
rect 15301 37281 15335 37315
rect 15485 37281 15519 37315
rect 16037 37281 16071 37315
rect 20729 37281 20763 37315
rect 21373 37281 21407 37315
rect 21557 37281 21591 37315
rect 21925 37281 21959 37315
rect 22109 37281 22143 37315
rect 22385 37281 22419 37315
rect 27169 37281 27203 37315
rect 32321 37281 32355 37315
rect 32873 37281 32907 37315
rect 33057 37281 33091 37315
rect 34345 37281 34379 37315
rect 40141 37281 40175 37315
rect 40969 37281 41003 37315
rect 44557 37281 44591 37315
rect 44841 37281 44875 37315
rect 51825 37281 51859 37315
rect 52009 37281 52043 37315
rect 52561 37281 52595 37315
rect 52745 37281 52779 37315
rect 60197 37281 60231 37315
rect 64337 37281 64371 37315
rect 64705 37281 64739 37315
rect 64797 37281 64831 37315
rect 65073 37281 65107 37315
rect 65809 37281 65843 37315
rect 66085 37281 66119 37315
rect 70133 37281 70167 37315
rect 70225 37281 70259 37315
rect 72249 37281 72283 37315
rect 73353 37281 73387 37315
rect 79480 37281 79514 37315
rect 81081 37281 81115 37315
rect 81541 37281 81575 37315
rect 85681 37281 85715 37315
rect 85957 37281 85991 37315
rect 88257 37281 88291 37315
rect 88441 37281 88475 37315
rect 88901 37281 88935 37315
rect 4445 37213 4479 37247
rect 9689 37213 9723 37247
rect 10425 37213 10459 37247
rect 22569 37213 22603 37247
rect 26893 37213 26927 37247
rect 28641 37213 28675 37247
rect 32137 37213 32171 37247
rect 38485 37213 38519 37247
rect 38761 37213 38795 37247
rect 44925 37213 44959 37247
rect 45201 37213 45235 37247
rect 64153 37213 64187 37247
rect 79701 37213 79735 37247
rect 85773 37213 85807 37247
rect 86509 37213 86543 37247
rect 20545 37145 20579 37179
rect 34529 37145 34563 37179
rect 65901 37145 65935 37179
rect 79609 37145 79643 37179
rect 15577 37077 15611 37111
rect 31953 37077 31987 37111
rect 34161 37077 34195 37111
rect 41061 37077 41095 37111
rect 44649 37077 44683 37111
rect 46765 37077 46799 37111
rect 63509 37077 63543 37111
rect 65257 37077 65291 37111
rect 79977 37077 80011 37111
rect 81173 37077 81207 37111
rect 88533 37077 88567 37111
rect 5457 36873 5491 36907
rect 9781 36873 9815 36907
rect 9965 36873 9999 36907
rect 33149 36873 33183 36907
rect 38669 36873 38703 36907
rect 43545 36873 43579 36907
rect 50721 36873 50755 36907
rect 64245 36873 64279 36907
rect 65533 36873 65567 36907
rect 78781 36873 78815 36907
rect 80069 36873 80103 36907
rect 83914 36873 83948 36907
rect 84761 36873 84795 36907
rect 85773 36873 85807 36907
rect 85957 36873 85991 36907
rect 86233 36873 86267 36907
rect 4997 36805 5031 36839
rect 16681 36805 16715 36839
rect 22293 36805 22327 36839
rect 26341 36805 26375 36839
rect 48237 36805 48271 36839
rect 51457 36805 51491 36839
rect 65349 36805 65383 36839
rect 66085 36805 66119 36839
rect 78965 36805 78999 36839
rect 81541 36805 81575 36839
rect 84025 36805 84059 36839
rect 8309 36737 8343 36771
rect 9137 36737 9171 36771
rect 20821 36737 20855 36771
rect 21557 36737 21591 36771
rect 22201 36737 22235 36771
rect 26433 36737 26467 36771
rect 37197 36737 37231 36771
rect 43269 36737 43303 36771
rect 46949 36737 46983 36771
rect 52009 36737 52043 36771
rect 64889 36737 64923 36771
rect 66453 36737 66487 36771
rect 71145 36737 71179 36771
rect 86693 36737 86727 36771
rect 87245 36737 87279 36771
rect 3893 36669 3927 36703
rect 4077 36669 4111 36703
rect 4629 36669 4663 36703
rect 4813 36669 4847 36703
rect 9045 36669 9079 36703
rect 9413 36669 9447 36703
rect 9597 36669 9631 36703
rect 13553 36669 13587 36703
rect 14289 36669 14323 36703
rect 14565 36669 14599 36703
rect 15945 36669 15979 36703
rect 16497 36669 16531 36703
rect 21465 36669 21499 36703
rect 21833 36669 21867 36703
rect 22017 36669 22051 36703
rect 26212 36669 26246 36703
rect 31953 36669 31987 36703
rect 32137 36669 32171 36703
rect 32689 36669 32723 36703
rect 32873 36669 32907 36703
rect 37473 36669 37507 36703
rect 37657 36669 37691 36703
rect 38255 36669 38289 36703
rect 38393 36669 38427 36703
rect 41797 36669 41831 36703
rect 41981 36669 42015 36703
rect 42165 36669 42199 36703
rect 42717 36669 42751 36703
rect 42901 36669 42935 36703
rect 46673 36669 46707 36703
rect 50629 36669 50663 36703
rect 51733 36669 51767 36703
rect 58173 36669 58207 36703
rect 58449 36669 58483 36703
rect 64429 36669 64463 36703
rect 64613 36669 64647 36703
rect 64981 36669 65015 36703
rect 65993 36669 66027 36703
rect 66269 36669 66303 36703
rect 70869 36669 70903 36703
rect 75929 36669 75963 36703
rect 78689 36669 78723 36703
rect 79793 36669 79827 36703
rect 79977 36669 80011 36703
rect 80437 36669 80471 36703
rect 81449 36669 81483 36703
rect 81725 36669 81759 36703
rect 84088 36669 84122 36703
rect 86785 36669 86819 36703
rect 87153 36669 87187 36703
rect 88165 36669 88199 36703
rect 88441 36669 88475 36703
rect 8401 36601 8435 36635
rect 15761 36601 15795 36635
rect 22477 36601 22511 36635
rect 26065 36601 26099 36635
rect 31861 36601 31895 36635
rect 59829 36601 59863 36635
rect 83749 36601 83783 36635
rect 84485 36601 84519 36635
rect 88349 36601 88383 36635
rect 88901 36601 88935 36635
rect 3709 36533 3743 36567
rect 5549 36533 5583 36567
rect 5733 36533 5767 36567
rect 13645 36533 13679 36567
rect 16037 36533 16071 36567
rect 25697 36533 25731 36567
rect 25881 36533 25915 36567
rect 26709 36533 26743 36567
rect 37381 36533 37415 36567
rect 48513 36533 48547 36567
rect 53113 36533 53147 36567
rect 59921 36533 59955 36567
rect 72433 36533 72467 36567
rect 72709 36533 72743 36567
rect 76113 36533 76147 36567
rect 81909 36533 81943 36567
rect 84577 36533 84611 36567
rect 85037 36533 85071 36567
rect 87981 36533 88015 36567
rect 5365 36329 5399 36363
rect 16497 36329 16531 36363
rect 17141 36329 17175 36363
rect 37473 36329 37507 36363
rect 56333 36329 56367 36363
rect 56517 36329 56551 36363
rect 68569 36329 68603 36363
rect 74549 36329 74583 36363
rect 74641 36329 74675 36363
rect 86601 36329 86635 36363
rect 33885 36261 33919 36295
rect 39037 36261 39071 36295
rect 47869 36261 47903 36295
rect 48145 36261 48179 36295
rect 52469 36261 52503 36295
rect 63233 36261 63267 36295
rect 67005 36261 67039 36295
rect 86785 36261 86819 36295
rect 87337 36261 87371 36295
rect 5273 36193 5307 36227
rect 5825 36193 5859 36227
rect 15301 36193 15335 36227
rect 16129 36193 16163 36227
rect 16313 36193 16347 36227
rect 17325 36193 17359 36227
rect 19717 36193 19751 36227
rect 21557 36193 21591 36227
rect 21925 36193 21959 36227
rect 22201 36193 22235 36227
rect 22477 36193 22511 36227
rect 26525 36193 26559 36227
rect 26672 36193 26706 36227
rect 32781 36193 32815 36227
rect 32873 36193 32907 36227
rect 33241 36193 33275 36227
rect 33333 36193 33367 36227
rect 37749 36193 37783 36227
rect 37933 36193 37967 36227
rect 38485 36193 38519 36227
rect 38669 36193 38703 36227
rect 45477 36193 45511 36227
rect 47777 36193 47811 36227
rect 57069 36193 57103 36227
rect 57621 36193 57655 36227
rect 57805 36193 57839 36227
rect 63141 36193 63175 36227
rect 67649 36193 67683 36227
rect 68017 36193 68051 36227
rect 71513 36193 71547 36227
rect 74825 36193 74859 36227
rect 75285 36193 75319 36227
rect 75377 36193 75411 36227
rect 79977 36193 80011 36227
rect 80069 36193 80103 36227
rect 85773 36193 85807 36227
rect 86049 36193 86083 36227
rect 86969 36193 87003 36227
rect 88717 36193 88751 36227
rect 15853 36125 15887 36159
rect 20913 36125 20947 36159
rect 21649 36125 21683 36159
rect 21833 36125 21867 36159
rect 26893 36125 26927 36159
rect 45201 36125 45235 36159
rect 50813 36125 50847 36159
rect 51089 36125 51123 36159
rect 56793 36125 56827 36159
rect 56885 36125 56919 36159
rect 67741 36125 67775 36159
rect 67925 36125 67959 36159
rect 71789 36125 71823 36159
rect 75837 36125 75871 36159
rect 88441 36125 88475 36159
rect 19901 36057 19935 36091
rect 27169 36057 27203 36091
rect 39221 36057 39255 36091
rect 68293 36057 68327 36091
rect 75101 36057 75135 36091
rect 85865 36057 85899 36091
rect 15117 35989 15151 36023
rect 17509 35989 17543 36023
rect 26249 35989 26283 36023
rect 26801 35989 26835 36023
rect 34161 35989 34195 36023
rect 34253 35989 34287 36023
rect 46765 35989 46799 36023
rect 46949 35989 46983 36023
rect 50629 35989 50663 36023
rect 58081 35989 58115 36023
rect 68753 35989 68787 36023
rect 72893 35989 72927 36023
rect 73353 35989 73387 36023
rect 79609 35989 79643 36023
rect 79793 35989 79827 36023
rect 80253 35989 80287 36023
rect 88257 35989 88291 36023
rect 89821 35989 89855 36023
rect 21649 35785 21683 35819
rect 26157 35785 26191 35819
rect 66085 35785 66119 35819
rect 67373 35785 67407 35819
rect 72249 35785 72283 35819
rect 76941 35785 76975 35819
rect 81357 35785 81391 35819
rect 6009 35717 6043 35751
rect 29469 35717 29503 35751
rect 47041 35717 47075 35751
rect 52009 35717 52043 35751
rect 85497 35717 85531 35751
rect 2605 35649 2639 35683
rect 2881 35649 2915 35683
rect 8677 35649 8711 35683
rect 16589 35649 16623 35683
rect 33333 35649 33367 35683
rect 44281 35649 44315 35683
rect 46857 35649 46891 35683
rect 58725 35649 58759 35683
rect 60105 35649 60139 35683
rect 67189 35649 67223 35683
rect 71421 35649 71455 35683
rect 71973 35649 72007 35683
rect 74733 35649 74767 35683
rect 75837 35649 75871 35683
rect 80069 35649 80103 35683
rect 85865 35649 85899 35683
rect 88349 35649 88383 35683
rect 4353 35581 4387 35615
rect 5365 35581 5399 35615
rect 5641 35581 5675 35615
rect 8401 35581 8435 35615
rect 10149 35581 10183 35615
rect 13369 35581 13403 35615
rect 14105 35581 14139 35615
rect 14381 35581 14415 35615
rect 15301 35581 15335 35615
rect 15853 35581 15887 35615
rect 16129 35581 16163 35615
rect 16313 35581 16347 35615
rect 20361 35581 20395 35615
rect 21465 35581 21499 35615
rect 21925 35581 21959 35615
rect 26341 35581 26375 35615
rect 26525 35581 26559 35615
rect 26893 35581 26927 35615
rect 26985 35581 27019 35615
rect 29285 35581 29319 35615
rect 32045 35581 32079 35615
rect 32229 35581 32263 35615
rect 32689 35581 32723 35615
rect 32781 35581 32815 35615
rect 33977 35581 34011 35615
rect 34161 35581 34195 35615
rect 42809 35581 42843 35615
rect 42993 35581 43027 35615
rect 43177 35581 43211 35615
rect 43729 35581 43763 35615
rect 43913 35581 43947 35615
rect 46949 35581 46983 35615
rect 51917 35581 51951 35615
rect 58449 35581 58483 35615
rect 63141 35581 63175 35615
rect 66269 35581 66303 35615
rect 66453 35581 66487 35615
rect 66821 35581 66855 35615
rect 66913 35581 66947 35615
rect 71513 35581 71547 35615
rect 74365 35581 74399 35615
rect 74825 35581 74859 35615
rect 75561 35581 75595 35615
rect 79793 35581 79827 35615
rect 85405 35581 85439 35615
rect 85681 35581 85715 35615
rect 86233 35581 86267 35615
rect 87889 35581 87923 35615
rect 88073 35581 88107 35615
rect 88533 35581 88567 35615
rect 15209 35513 15243 35547
rect 29745 35513 29779 35547
rect 74178 35513 74212 35547
rect 4169 35445 4203 35479
rect 5181 35445 5215 35479
rect 9781 35445 9815 35479
rect 13461 35445 13495 35479
rect 16497 35445 16531 35479
rect 20545 35445 20579 35479
rect 27169 35445 27203 35479
rect 27445 35445 27479 35479
rect 33517 35445 33551 35479
rect 33701 35445 33735 35479
rect 44465 35445 44499 35479
rect 60197 35445 60231 35479
rect 63233 35445 63267 35479
rect 65625 35445 65659 35479
rect 72157 35445 72191 35479
rect 75009 35445 75043 35479
rect 77309 35445 77343 35479
rect 79517 35445 79551 35479
rect 4629 35241 4663 35275
rect 5457 35241 5491 35275
rect 6193 35241 6227 35275
rect 16957 35241 16991 35275
rect 17509 35241 17543 35275
rect 21097 35241 21131 35275
rect 21373 35241 21407 35275
rect 32689 35241 32723 35275
rect 32965 35241 32999 35275
rect 48789 35241 48823 35275
rect 26525 35173 26559 35207
rect 36369 35173 36403 35207
rect 38393 35173 38427 35207
rect 40141 35173 40175 35207
rect 44557 35173 44591 35207
rect 44833 35173 44867 35207
rect 4813 35105 4847 35139
rect 5089 35105 5123 35139
rect 6101 35105 6135 35139
rect 6653 35105 6687 35139
rect 14105 35105 14139 35139
rect 16957 35105 16991 35139
rect 17049 35105 17083 35139
rect 20913 35105 20947 35139
rect 27169 35105 27203 35139
rect 27537 35105 27571 35139
rect 32505 35105 32539 35139
rect 36553 35105 36587 35139
rect 43361 35105 43395 35139
rect 43729 35105 43763 35139
rect 44465 35105 44499 35139
rect 27261 35037 27295 35071
rect 27445 35037 27479 35071
rect 27905 35037 27939 35071
rect 38485 35037 38519 35071
rect 38761 35037 38795 35071
rect 43177 35037 43211 35071
rect 28089 34969 28123 35003
rect 36737 34969 36771 35003
rect 13921 34901 13955 34935
rect 14197 34901 14231 34935
rect 17233 34901 17267 34935
rect 43177 34901 43211 34935
rect 43545 34901 43579 34935
rect 48789 34901 48823 34935
rect 55321 35241 55355 35275
rect 57253 35241 57287 35275
rect 79517 35241 79551 35275
rect 88349 35241 88383 35275
rect 55505 35105 55539 35139
rect 55689 35105 55723 35139
rect 56241 35105 56275 35139
rect 56793 35105 56827 35139
rect 56977 35105 57011 35139
rect 57621 35105 57655 35139
rect 67925 35105 67959 35139
rect 72065 35105 72099 35139
rect 72341 35105 72375 35139
rect 75009 35105 75043 35139
rect 75193 35105 75227 35139
rect 77033 35105 77067 35139
rect 79333 35105 79367 35139
rect 88257 35105 88291 35139
rect 55321 35037 55355 35071
rect 55873 35037 55907 35071
rect 56057 35037 56091 35071
rect 75561 35037 75595 35071
rect 72157 34969 72191 35003
rect 55321 34901 55355 34935
rect 68017 34901 68051 34935
rect 75745 34901 75779 34935
rect 77125 34901 77159 34935
rect 5549 34697 5583 34731
rect 21833 34697 21867 34731
rect 22109 34697 22143 34731
rect 27353 34697 27387 34731
rect 37013 34697 37047 34731
rect 39681 34697 39715 34731
rect 40325 34697 40359 34731
rect 51457 34697 51491 34731
rect 53297 34697 53331 34731
rect 62681 34697 62715 34731
rect 64429 34697 64463 34731
rect 67741 34697 67775 34731
rect 68109 34697 68143 34731
rect 76665 34697 76699 34731
rect 77125 34697 77159 34731
rect 7297 34629 7331 34663
rect 15117 34629 15151 34663
rect 21925 34629 21959 34663
rect 44281 34629 44315 34663
rect 44649 34629 44683 34663
rect 44833 34629 44867 34663
rect 60841 34629 60875 34663
rect 61209 34629 61243 34663
rect 64061 34629 64095 34663
rect 64705 34629 64739 34663
rect 20269 34561 20303 34595
rect 21005 34561 21039 34595
rect 21649 34561 21683 34595
rect 36645 34561 36679 34595
rect 40325 34561 40359 34595
rect 51917 34561 51951 34595
rect 52653 34561 52687 34595
rect 59461 34561 59495 34595
rect 59737 34561 59771 34595
rect 68293 34629 68327 34663
rect 85497 34629 85531 34663
rect 67925 34561 67959 34595
rect 68569 34561 68603 34595
rect 75653 34561 75687 34595
rect 89453 34561 89487 34595
rect 4905 34493 4939 34527
rect 5181 34493 5215 34527
rect 7113 34493 7147 34527
rect 8217 34493 8251 34527
rect 8769 34493 8803 34527
rect 13093 34493 13127 34527
rect 15761 34493 15795 34527
rect 16037 34493 16071 34527
rect 16221 34493 16255 34527
rect 20913 34493 20947 34527
rect 21281 34493 21315 34527
rect 21465 34493 21499 34527
rect 25789 34493 25823 34527
rect 26065 34493 26099 34527
rect 37197 34493 37231 34527
rect 37381 34493 37415 34527
rect 37749 34493 37783 34527
rect 37933 34493 37967 34527
rect 39313 34493 39347 34527
rect 42901 34493 42935 34527
rect 43085 34493 43119 34527
rect 43269 34493 43303 34527
rect 43729 34493 43763 34527
rect 43821 34493 43855 34527
rect 51733 34493 51767 34527
rect 52561 34493 52595 34527
rect 52929 34493 52963 34527
rect 53113 34493 53147 34527
rect 62957 34493 62991 34527
rect 63141 34493 63175 34527
rect 63601 34493 63635 34527
rect 63693 34493 63727 34527
rect 65625 34493 65659 34527
rect 67741 34493 67775 34527
rect 68753 34493 68787 34527
rect 69213 34493 69247 34527
rect 69305 34493 69339 34527
rect 75561 34493 75595 34527
rect 75837 34493 75871 34527
rect 77033 34493 77067 34527
rect 85405 34493 85439 34527
rect 88165 34493 88199 34527
rect 89361 34493 89395 34527
rect 5365 34425 5399 34459
rect 8953 34425 8987 34459
rect 15209 34425 15243 34459
rect 65717 34425 65751 34459
rect 76849 34425 76883 34459
rect 87981 34425 88015 34459
rect 88533 34425 88567 34459
rect 13185 34357 13219 34391
rect 27537 34357 27571 34391
rect 36461 34357 36495 34391
rect 39405 34357 39439 34391
rect 54401 34357 54435 34391
rect 62405 34357 62439 34391
rect 69765 34357 69799 34391
rect 70133 34357 70167 34391
rect 76113 34357 76147 34391
rect 4353 34153 4387 34187
rect 5733 34153 5767 34187
rect 9321 34153 9355 34187
rect 11529 34153 11563 34187
rect 16037 34153 16071 34187
rect 75193 34153 75227 34187
rect 87981 34153 88015 34187
rect 16681 34085 16715 34119
rect 37197 34085 37231 34119
rect 37381 34085 37415 34119
rect 39037 34085 39071 34119
rect 50629 34085 50663 34119
rect 56793 34085 56827 34119
rect 58265 34085 58299 34119
rect 64705 34085 64739 34119
rect 74549 34085 74583 34119
rect 85037 34085 85071 34119
rect 4537 34017 4571 34051
rect 4629 34017 4663 34051
rect 5549 34017 5583 34051
rect 9505 34017 9539 34051
rect 11989 34017 12023 34051
rect 15577 34017 15611 34051
rect 15669 34017 15703 34051
rect 15853 34017 15887 34051
rect 18429 34017 18463 34051
rect 18705 34017 18739 34051
rect 19073 34017 19107 34051
rect 21649 34017 21683 34051
rect 21741 34017 21775 34051
rect 25421 34017 25455 34051
rect 25513 34017 25547 34051
rect 26709 34017 26743 34051
rect 27261 34017 27295 34051
rect 27445 34017 27479 34051
rect 28089 34017 28123 34051
rect 28273 34017 28307 34051
rect 32137 34017 32171 34051
rect 37933 34017 37967 34051
rect 38485 34017 38519 34051
rect 38669 34017 38703 34051
rect 44649 34017 44683 34051
rect 49525 34017 49559 34051
rect 50077 34017 50111 34051
rect 50261 34017 50295 34051
rect 54769 34017 54803 34051
rect 55321 34017 55355 34051
rect 55505 34017 55539 34051
rect 56057 34017 56091 34051
rect 56977 34017 57011 34051
rect 57161 34017 57195 34051
rect 57713 34017 57747 34051
rect 57897 34017 57931 34051
rect 63325 34017 63359 34051
rect 67465 34017 67499 34051
rect 68937 34017 68971 34051
rect 73261 34017 73295 34051
rect 73997 34017 74031 34051
rect 75377 34017 75411 34051
rect 77217 34017 77251 34051
rect 77309 34017 77343 34051
rect 87153 34017 87187 34051
rect 88257 34017 88291 34051
rect 88441 34017 88475 34051
rect 88533 34017 88567 34051
rect 89821 34017 89855 34051
rect 11713 33949 11747 33983
rect 17877 33949 17911 33983
rect 18889 33949 18923 33983
rect 26249 33949 26283 33983
rect 26525 33949 26559 33983
rect 37565 33949 37599 33983
rect 37749 33949 37783 33983
rect 44373 33949 44407 33983
rect 45753 33949 45787 33983
rect 49341 33949 49375 33983
rect 54585 33949 54619 33983
rect 56701 33949 56735 33983
rect 62865 33949 62899 33983
rect 63049 33949 63083 33983
rect 67189 33949 67223 33983
rect 68569 33949 68603 33983
rect 74273 33949 74307 33983
rect 75745 33949 75779 33983
rect 76113 33949 76147 33983
rect 83381 33949 83415 33983
rect 83657 33949 83691 33983
rect 21925 33881 21959 33915
rect 48697 33881 48731 33915
rect 54033 33881 54067 33915
rect 54217 33881 54251 33915
rect 55781 33881 55815 33915
rect 73537 33881 73571 33915
rect 75653 33881 75687 33915
rect 77033 33881 77067 33915
rect 90005 33881 90039 33915
rect 13093 33813 13127 33847
rect 16497 33813 16531 33847
rect 21649 33813 21683 33847
rect 27721 33813 27755 33847
rect 32229 33813 32263 33847
rect 37013 33813 37047 33847
rect 37565 33813 37599 33847
rect 48973 33813 49007 33847
rect 49157 33813 49191 33847
rect 58541 33813 58575 33847
rect 58633 33813 58667 33847
rect 75542 33813 75576 33847
rect 76205 33813 76239 33847
rect 77493 33813 77527 33847
rect 83197 33813 83231 33847
rect 87245 33813 87279 33847
rect 88717 33813 88751 33847
rect 4445 33609 4479 33643
rect 49249 33609 49283 33643
rect 50629 33609 50663 33643
rect 53941 33609 53975 33643
rect 56885 33609 56919 33643
rect 59001 33609 59035 33643
rect 68734 33609 68768 33643
rect 85497 33609 85531 33643
rect 87061 33609 87095 33643
rect 89821 33609 89855 33643
rect 9689 33541 9723 33575
rect 15025 33541 15059 33575
rect 17325 33541 17359 33575
rect 18153 33541 18187 33575
rect 18981 33541 19015 33575
rect 24869 33541 24903 33575
rect 26341 33541 26375 33575
rect 32137 33541 32171 33575
rect 33149 33541 33183 33575
rect 60933 33541 60967 33575
rect 68845 33541 68879 33575
rect 2605 33473 2639 33507
rect 2881 33473 2915 33507
rect 37289 33473 37323 33507
rect 38025 33473 38059 33507
rect 49433 33473 49467 33507
rect 51365 33473 51399 33507
rect 52561 33473 52595 33507
rect 53297 33473 53331 33507
rect 55321 33473 55355 33507
rect 57345 33473 57379 33507
rect 61025 33473 61059 33507
rect 68937 33473 68971 33507
rect 76297 33473 76331 33507
rect 80805 33473 80839 33507
rect 80897 33473 80931 33507
rect 88533 33473 88567 33507
rect 7389 33405 7423 33439
rect 8769 33405 8803 33439
rect 9321 33405 9355 33439
rect 15209 33405 15243 33439
rect 15301 33405 15335 33439
rect 16589 33405 16623 33439
rect 16773 33405 16807 33439
rect 18061 33405 18095 33439
rect 18337 33405 18371 33439
rect 19901 33405 19935 33439
rect 24961 33405 24995 33439
rect 25237 33405 25271 33439
rect 27445 33405 27479 33439
rect 30573 33405 30607 33439
rect 30849 33405 30883 33439
rect 33057 33405 33091 33439
rect 35449 33405 35483 33439
rect 35633 33405 35667 33439
rect 37013 33405 37047 33439
rect 37933 33405 37967 33439
rect 38301 33405 38335 33439
rect 38485 33405 38519 33439
rect 49617 33405 49651 33439
rect 50169 33405 50203 33439
rect 50353 33405 50387 33439
rect 52469 33405 52503 33439
rect 52837 33405 52871 33439
rect 53021 33405 53055 33439
rect 54217 33405 54251 33439
rect 54309 33405 54343 33439
rect 54769 33405 54803 33439
rect 54953 33405 54987 33439
rect 57529 33405 57563 33439
rect 57989 33405 58023 33439
rect 58169 33405 58203 33439
rect 60804 33405 60838 33439
rect 61393 33405 61427 33439
rect 69305 33405 69339 33439
rect 76021 33405 76055 33439
rect 77769 33405 77803 33439
rect 81173 33405 81207 33439
rect 85405 33405 85439 33439
rect 86969 33405 87003 33439
rect 88257 33405 88291 33439
rect 51457 33337 51491 33371
rect 51825 33337 51859 33371
rect 53481 33337 53515 33371
rect 53665 33337 53699 33371
rect 57069 33337 57103 33371
rect 58633 33337 58667 33371
rect 60657 33337 60691 33371
rect 68569 33337 68603 33371
rect 86785 33337 86819 33371
rect 4169 33269 4203 33303
rect 7573 33269 7607 33303
rect 9045 33269 9079 33303
rect 16865 33269 16899 33303
rect 17877 33269 17911 33303
rect 18521 33269 18555 33303
rect 19993 33269 20027 33303
rect 27537 33269 27571 33303
rect 32321 33269 32355 33303
rect 33333 33269 33367 33303
rect 35817 33269 35851 33303
rect 37197 33269 37231 33303
rect 48881 33269 48915 33303
rect 49065 33269 49099 33303
rect 53205 33269 53239 33303
rect 55597 33269 55631 33303
rect 58909 33269 58943 33303
rect 77401 33269 77435 33303
rect 82277 33269 82311 33303
rect 86693 33269 86727 33303
rect 88073 33269 88107 33303
rect 8953 33065 8987 33099
rect 10609 33065 10643 33099
rect 49433 33065 49467 33099
rect 63693 33065 63727 33099
rect 68753 33065 68787 33099
rect 75561 33065 75595 33099
rect 77769 33065 77803 33099
rect 85313 33065 85347 33099
rect 88533 33065 88567 33099
rect 15025 32997 15059 33031
rect 17877 32997 17911 33031
rect 29285 32997 29319 33031
rect 29377 32997 29411 33031
rect 31033 32997 31067 33031
rect 49157 32997 49191 33031
rect 67005 32997 67039 33031
rect 68845 32997 68879 33031
rect 85681 32997 85715 33031
rect 88257 32997 88291 33031
rect 8033 32929 8067 32963
rect 8585 32929 8619 32963
rect 9689 32929 9723 32963
rect 10241 32929 10275 32963
rect 15301 32929 15335 32963
rect 17785 32929 17819 32963
rect 19625 32929 19659 32963
rect 20913 32929 20947 32963
rect 29929 32929 29963 32963
rect 30389 32929 30423 32963
rect 30481 32929 30515 32963
rect 31861 32929 31895 32963
rect 32321 32929 32355 32963
rect 32873 32929 32907 32963
rect 33057 32929 33091 32963
rect 38117 32929 38151 32963
rect 42165 32929 42199 32963
rect 45477 32929 45511 32963
rect 46305 32929 46339 32963
rect 49065 32929 49099 32963
rect 49985 32929 50019 32963
rect 50353 32929 50387 32963
rect 50537 32929 50571 32963
rect 61853 32929 61887 32963
rect 62037 32929 62071 32963
rect 62497 32929 62531 32963
rect 62589 32929 62623 32963
rect 63325 32929 63359 32963
rect 67373 32929 67407 32963
rect 67465 32929 67499 32963
rect 67925 32929 67959 32963
rect 68109 32929 68143 32963
rect 73997 32929 74031 32963
rect 74273 32929 74307 32963
rect 74457 32929 74491 32963
rect 75469 32929 75503 32963
rect 75745 32929 75779 32963
rect 77953 32929 77987 32963
rect 80437 32929 80471 32963
rect 80529 32929 80563 32963
rect 81449 32929 81483 32963
rect 82185 32929 82219 32963
rect 82645 32929 82679 32963
rect 83197 32929 83231 32963
rect 86325 32929 86359 32963
rect 86693 32929 86727 32963
rect 86785 32929 86819 32963
rect 88441 32929 88475 32963
rect 88901 32929 88935 32963
rect 8677 32861 8711 32895
rect 10425 32861 10459 32895
rect 15577 32861 15611 32895
rect 29745 32861 29779 32895
rect 31493 32861 31527 32895
rect 32137 32861 32171 32895
rect 43821 32861 43855 32895
rect 44097 32861 44131 32895
rect 50077 32861 50111 32895
rect 68477 32861 68511 32895
rect 73445 32861 73479 32895
rect 83473 32861 83507 32895
rect 86233 32861 86267 32895
rect 19809 32793 19843 32827
rect 21097 32793 21131 32827
rect 31217 32793 31251 32827
rect 33609 32793 33643 32827
rect 42349 32793 42383 32827
rect 61669 32793 61703 32827
rect 81633 32793 81667 32827
rect 82737 32793 82771 32827
rect 16681 32725 16715 32759
rect 17601 32725 17635 32759
rect 29561 32725 29595 32759
rect 31493 32725 31527 32759
rect 31585 32725 31619 32759
rect 33333 32725 33367 32759
rect 37933 32725 37967 32759
rect 38301 32725 38335 32759
rect 41981 32725 42015 32759
rect 46397 32725 46431 32759
rect 63049 32725 63083 32759
rect 63509 32725 63543 32759
rect 82369 32725 82403 32759
rect 85589 32725 85623 32759
rect 10425 32521 10459 32555
rect 35449 32521 35483 32555
rect 36185 32521 36219 32555
rect 37657 32521 37691 32555
rect 42165 32521 42199 32555
rect 54585 32521 54619 32555
rect 15853 32453 15887 32487
rect 16865 32453 16899 32487
rect 18705 32453 18739 32487
rect 21373 32453 21407 32487
rect 21557 32453 21591 32487
rect 27261 32453 27295 32487
rect 40785 32453 40819 32487
rect 42441 32453 42475 32487
rect 42993 32453 43027 32487
rect 54769 32453 54803 32487
rect 61669 32453 61703 32487
rect 69673 32453 69707 32487
rect 3157 32385 3191 32419
rect 8493 32385 8527 32419
rect 8861 32385 8895 32419
rect 10057 32385 10091 32419
rect 24777 32385 24811 32419
rect 24961 32385 24995 32419
rect 26065 32385 26099 32419
rect 26433 32385 26467 32419
rect 26617 32385 26651 32419
rect 31585 32385 31619 32419
rect 31861 32385 31895 32419
rect 37289 32385 37323 32419
rect 40969 32385 41003 32419
rect 53205 32385 53239 32419
rect 54309 32385 54343 32419
rect 81541 32385 81575 32419
rect 82093 32385 82127 32419
rect 82553 32385 82587 32419
rect 82645 32385 82679 32419
rect 2881 32317 2915 32351
rect 8033 32317 8067 32351
rect 8401 32317 8435 32351
rect 9689 32317 9723 32351
rect 9965 32317 9999 32351
rect 15669 32317 15703 32351
rect 16773 32317 16807 32351
rect 18613 32317 18647 32351
rect 19993 32317 20027 32351
rect 20085 32317 20119 32351
rect 20545 32317 20579 32351
rect 20729 32317 20763 32351
rect 25053 32317 25087 32351
rect 25605 32317 25639 32351
rect 25789 32317 25823 32351
rect 27077 32317 27111 32351
rect 33241 32317 33275 32351
rect 35265 32317 35299 32351
rect 36369 32317 36403 32351
rect 37473 32317 37507 32351
rect 41153 32317 41187 32351
rect 41613 32317 41647 32351
rect 41705 32317 41739 32351
rect 42625 32317 42659 32351
rect 43177 32317 43211 32351
rect 44373 32317 44407 32351
rect 48145 32317 48179 32351
rect 53297 32317 53331 32351
rect 53757 32317 53791 32351
rect 53849 32317 53883 32351
rect 60565 32317 60599 32351
rect 60749 32317 60783 32351
rect 61301 32317 61335 32351
rect 61485 32317 61519 32351
rect 62129 32317 62163 32351
rect 68569 32317 68603 32351
rect 68753 32317 68787 32351
rect 69213 32317 69247 32351
rect 69305 32317 69339 32351
rect 70041 32317 70075 32351
rect 74181 32317 74215 32351
rect 74457 32317 74491 32351
rect 82369 32317 82403 32351
rect 21741 32249 21775 32283
rect 40601 32249 40635 32283
rect 44465 32249 44499 32283
rect 62221 32249 62255 32283
rect 75929 32249 75963 32283
rect 4261 32181 4295 32215
rect 4721 32181 4755 32215
rect 21005 32181 21039 32215
rect 26893 32181 26927 32215
rect 33333 32181 33367 32215
rect 35081 32181 35115 32215
rect 36553 32181 36587 32215
rect 43361 32181 43395 32215
rect 47961 32181 47995 32215
rect 55045 32181 55079 32215
rect 60381 32181 60415 32215
rect 62405 32181 62439 32215
rect 68293 32181 68327 32215
rect 75561 32181 75595 32215
rect 10885 31977 10919 32011
rect 34897 31977 34931 32011
rect 40969 31977 41003 32011
rect 42625 31977 42659 32011
rect 42809 31977 42843 32011
rect 44741 31977 44775 32011
rect 53389 31977 53423 32011
rect 54401 31977 54435 32011
rect 54861 31977 54895 32011
rect 68753 31977 68787 32011
rect 74457 31977 74491 32011
rect 76021 31977 76055 32011
rect 76297 31977 76331 32011
rect 81173 31977 81207 32011
rect 88441 31977 88475 32011
rect 42349 31909 42383 31943
rect 87429 31909 87463 31943
rect 10977 31841 11011 31875
rect 16497 31841 16531 31875
rect 17049 31841 17083 31875
rect 17233 31841 17267 31875
rect 17417 31841 17451 31875
rect 17877 31841 17911 31875
rect 19533 31841 19567 31875
rect 34713 31841 34747 31875
rect 41245 31841 41279 31875
rect 41885 31841 41919 31875
rect 41981 31841 42015 31875
rect 43637 31841 43671 31875
rect 53297 31841 53331 31875
rect 54401 31841 54435 31875
rect 54585 31841 54619 31875
rect 67465 31841 67499 31875
rect 67925 31841 67959 31875
rect 68017 31841 68051 31875
rect 74365 31841 74399 31875
rect 74641 31841 74675 31875
rect 75837 31841 75871 31875
rect 80529 31841 80563 31875
rect 80676 31841 80710 31875
rect 81357 31841 81391 31875
rect 85405 31841 85439 31875
rect 86785 31841 86819 31875
rect 86969 31841 87003 31875
rect 87337 31841 87371 31875
rect 88257 31841 88291 31875
rect 11253 31773 11287 31807
rect 16221 31773 16255 31807
rect 16589 31773 16623 31807
rect 17969 31773 18003 31807
rect 19441 31773 19475 31807
rect 34529 31773 34563 31807
rect 41061 31773 41095 31807
rect 43361 31773 43395 31807
rect 66913 31773 66947 31807
rect 67281 31773 67315 31807
rect 80897 31773 80931 31807
rect 85497 31773 85531 31807
rect 18245 31705 18279 31739
rect 40785 31705 40819 31739
rect 12541 31637 12575 31671
rect 19717 31637 19751 31671
rect 53113 31637 53147 31671
rect 54677 31637 54711 31671
rect 67097 31637 67131 31671
rect 68477 31637 68511 31671
rect 69029 31637 69063 31671
rect 80805 31637 80839 31671
rect 12081 31433 12115 31467
rect 12173 31433 12207 31467
rect 3157 31297 3191 31331
rect 57161 31433 57195 31467
rect 62129 31433 62163 31467
rect 63233 31433 63267 31467
rect 63601 31433 63635 31467
rect 68707 31433 68741 31467
rect 68845 31433 68879 31467
rect 75745 31433 75779 31467
rect 75929 31433 75963 31467
rect 84209 31433 84243 31467
rect 85129 31433 85163 31467
rect 23765 31365 23799 31399
rect 35265 31365 35299 31399
rect 35541 31365 35575 31399
rect 41981 31365 42015 31399
rect 16129 31297 16163 31331
rect 69029 31365 69063 31399
rect 85497 31365 85531 31399
rect 24777 31297 24811 31331
rect 46581 31297 46615 31331
rect 46765 31297 46799 31331
rect 57161 31297 57195 31331
rect 61945 31297 61979 31331
rect 63104 31297 63138 31331
rect 63325 31297 63359 31331
rect 68937 31297 68971 31331
rect 74181 31297 74215 31331
rect 2881 31229 2915 31263
rect 11897 31229 11931 31263
rect 12173 31229 12207 31263
rect 15761 31229 15795 31263
rect 23765 31229 23799 31263
rect 23857 31229 23891 31263
rect 24685 31229 24719 31263
rect 25054 31229 25088 31263
rect 25145 31229 25179 31263
rect 29285 31229 29319 31263
rect 35357 31229 35391 31263
rect 36461 31229 36495 31263
rect 36737 31229 36771 31263
rect 42073 31229 42107 31263
rect 43177 31229 43211 31263
rect 47133 31229 47167 31263
rect 47317 31229 47351 31263
rect 47869 31229 47903 31263
rect 48053 31229 48087 31263
rect 53665 31229 53699 31263
rect 53757 31229 53791 31263
rect 54125 31229 54159 31263
rect 54217 31229 54251 31263
rect 55137 31229 55171 31263
rect 59001 31229 59035 31263
rect 60657 31229 60691 31263
rect 60841 31229 60875 31263
rect 61301 31229 61335 31263
rect 61393 31229 61427 31263
rect 74365 31229 74399 31263
rect 74825 31229 74859 31263
rect 74917 31229 74951 31263
rect 79793 31229 79827 31263
rect 79977 31229 80011 31263
rect 80437 31229 80471 31263
rect 82369 31229 82403 31263
rect 82737 31229 82771 31263
rect 83657 31229 83691 31263
rect 83749 31229 83783 31263
rect 83933 31229 83967 31263
rect 84025 31229 84059 31263
rect 85681 31229 85715 31263
rect 85957 31229 85991 31263
rect 87429 31229 87463 31263
rect 87705 31229 87739 31263
rect 15577 31161 15611 31195
rect 24041 31161 24075 31195
rect 38117 31161 38151 31195
rect 48421 31161 48455 31195
rect 54953 31161 54987 31195
rect 60289 31161 60323 31195
rect 62957 31161 62991 31195
rect 68569 31161 68603 31195
rect 80345 31161 80379 31195
rect 82185 31161 82219 31195
rect 87613 31161 87647 31195
rect 88165 31161 88199 31195
rect 4261 31093 4295 31127
rect 4721 31093 4755 31127
rect 11713 31093 11747 31127
rect 29377 31093 29411 31127
rect 29653 31093 29687 31127
rect 42257 31093 42291 31127
rect 43269 31093 43303 31127
rect 43545 31093 43579 31127
rect 46949 31093 46983 31127
rect 54677 31093 54711 31127
rect 59093 31093 59127 31127
rect 60473 31093 60507 31127
rect 62313 31093 62347 31127
rect 73721 31093 73755 31127
rect 73905 31093 73939 31127
rect 75377 31093 75411 31127
rect 87245 31093 87279 31127
rect 13001 30889 13035 30923
rect 18245 30889 18279 30923
rect 25237 30889 25271 30923
rect 30941 30889 30975 30923
rect 36921 30889 36955 30923
rect 66085 30889 66119 30923
rect 67465 30889 67499 30923
rect 68293 30889 68327 30923
rect 69673 30889 69707 30923
rect 86233 30889 86267 30923
rect 87981 30889 88015 30923
rect 89729 30889 89763 30923
rect 11161 30821 11195 30855
rect 35265 30821 35299 30855
rect 36737 30821 36771 30855
rect 5181 30753 5215 30787
rect 11069 30753 11103 30787
rect 11713 30753 11747 30787
rect 11805 30753 11839 30787
rect 12081 30753 12115 30787
rect 12633 30753 12667 30787
rect 16957 30753 16991 30787
rect 19441 30753 19475 30787
rect 24041 30753 24075 30787
rect 25053 30753 25087 30787
rect 35449 30753 35483 30787
rect 35633 30753 35667 30787
rect 36185 30753 36219 30787
rect 36369 30753 36403 30787
rect 4905 30685 4939 30719
rect 12449 30685 12483 30719
rect 16497 30685 16531 30719
rect 16681 30685 16715 30719
rect 29101 30685 29135 30719
rect 29377 30685 29411 30719
rect 62405 30821 62439 30855
rect 68109 30821 68143 30855
rect 74825 30821 74859 30855
rect 75101 30821 75135 30855
rect 75193 30821 75227 30855
rect 83749 30821 83783 30855
rect 86417 30821 86451 30855
rect 37105 30753 37139 30787
rect 37289 30753 37323 30787
rect 37933 30753 37967 30787
rect 38393 30753 38427 30787
rect 38485 30753 38519 30787
rect 40969 30753 41003 30787
rect 41153 30753 41187 30787
rect 41705 30753 41739 30787
rect 41889 30753 41923 30787
rect 42441 30753 42475 30787
rect 43361 30753 43395 30787
rect 46397 30753 46431 30787
rect 46949 30753 46983 30787
rect 47133 30753 47167 30787
rect 49249 30753 49283 30787
rect 54585 30753 54619 30787
rect 56241 30753 56275 30787
rect 56425 30753 56459 30787
rect 56885 30753 56919 30787
rect 57437 30753 57471 30787
rect 57621 30753 57655 30787
rect 58909 30753 58943 30787
rect 61301 30753 61335 30787
rect 61767 30753 61801 30787
rect 61941 30753 61975 30787
rect 62773 30753 62807 30787
rect 66453 30753 66487 30787
rect 66913 30753 66947 30787
rect 67005 30753 67039 30787
rect 68477 30753 68511 30787
rect 68661 30753 68695 30787
rect 69121 30753 69155 30787
rect 69213 30753 69247 30787
rect 70133 30753 70167 30787
rect 73721 30753 73755 30787
rect 74181 30753 74215 30787
rect 74273 30753 74307 30787
rect 79517 30753 79551 30787
rect 79609 30753 79643 30787
rect 79885 30753 79919 30787
rect 80897 30753 80931 30787
rect 84209 30753 84243 30787
rect 86601 30753 86635 30787
rect 88349 30753 88383 30787
rect 88625 30753 88659 30787
rect 37749 30685 37783 30719
rect 40785 30685 40819 30719
rect 42257 30685 42291 30719
rect 46213 30685 46247 30719
rect 48973 30685 49007 30719
rect 56609 30685 56643 30719
rect 56701 30685 56735 30719
rect 61025 30685 61059 30719
rect 61117 30685 61151 30719
rect 66269 30685 66303 30719
rect 73537 30685 73571 30719
rect 78781 30685 78815 30719
rect 79977 30685 80011 30719
rect 80713 30685 80747 30719
rect 83933 30685 83967 30719
rect 12817 30617 12851 30651
rect 30665 30617 30699 30651
rect 36921 30617 36955 30651
rect 38853 30617 38887 30651
rect 40509 30617 40543 30651
rect 40693 30617 40727 30651
rect 46029 30617 46063 30651
rect 57805 30617 57839 30651
rect 59001 30617 59035 30651
rect 80161 30617 80195 30651
rect 81081 30617 81115 30651
rect 6285 30549 6319 30583
rect 6653 30549 6687 30583
rect 19625 30549 19659 30583
rect 24133 30549 24167 30583
rect 37473 30549 37507 30583
rect 43453 30549 43487 30583
rect 43729 30549 43763 30583
rect 47409 30549 47443 30583
rect 48789 30549 48823 30583
rect 50353 30549 50387 30583
rect 54677 30549 54711 30583
rect 59185 30549 59219 30583
rect 60749 30549 60783 30583
rect 62681 30549 62715 30583
rect 67741 30549 67775 30583
rect 68017 30549 68051 30583
rect 70041 30549 70075 30583
rect 73169 30549 73203 30583
rect 73353 30549 73387 30583
rect 78965 30549 78999 30583
rect 85313 30549 85347 30583
rect 86693 30549 86727 30583
rect 31033 30345 31067 30379
rect 38209 30345 38243 30379
rect 54125 30345 54159 30379
rect 60197 30345 60231 30379
rect 84669 30345 84703 30379
rect 28181 30277 28215 30311
rect 37565 30277 37599 30311
rect 43177 30277 43211 30311
rect 48789 30277 48823 30311
rect 52561 30277 52595 30311
rect 61485 30277 61519 30311
rect 61945 30277 61979 30311
rect 65717 30277 65751 30311
rect 65901 30277 65935 30311
rect 71421 30277 71455 30311
rect 84393 30277 84427 30311
rect 2605 30209 2639 30243
rect 4629 30209 4663 30243
rect 9965 30209 9999 30243
rect 25053 30209 25087 30243
rect 52745 30209 52779 30243
rect 58817 30209 58851 30243
rect 66269 30209 66303 30243
rect 68661 30209 68695 30243
rect 87705 30209 87739 30243
rect 2881 30141 2915 30175
rect 7941 30141 7975 30175
rect 10609 30141 10643 30175
rect 10793 30141 10827 30175
rect 10977 30141 11011 30175
rect 11345 30141 11379 30175
rect 11529 30141 11563 30175
rect 15485 30141 15519 30175
rect 19809 30141 19843 30175
rect 21833 30141 21867 30175
rect 22017 30141 22051 30175
rect 24777 30141 24811 30175
rect 24961 30141 24995 30175
rect 25421 30141 25455 30175
rect 26985 30141 27019 30175
rect 27169 30141 27203 30175
rect 27629 30141 27663 30175
rect 27809 30141 27843 30175
rect 29285 30141 29319 30175
rect 29561 30141 29595 30175
rect 35633 30141 35667 30175
rect 35909 30141 35943 30175
rect 37473 30141 37507 30175
rect 38117 30141 38151 30175
rect 41613 30141 41647 30175
rect 41889 30141 41923 30175
rect 43361 30141 43395 30175
rect 43637 30141 43671 30175
rect 46949 30141 46983 30175
rect 47225 30141 47259 30175
rect 53021 30141 53055 30175
rect 57437 30141 57471 30175
rect 57713 30141 57747 30175
rect 59737 30141 59771 30175
rect 60381 30141 60415 30175
rect 60565 30141 60599 30175
rect 61025 30141 61059 30175
rect 61205 30141 61239 30175
rect 62037 30141 62071 30175
rect 66453 30141 66487 30175
rect 67005 30141 67039 30175
rect 67189 30141 67223 30175
rect 68569 30141 68603 30175
rect 74365 30141 74399 30175
rect 79793 30141 79827 30175
rect 80069 30141 80103 30175
rect 84301 30141 84335 30175
rect 86141 30141 86175 30175
rect 86325 30141 86359 30175
rect 86693 30141 86727 30175
rect 87613 30141 87647 30175
rect 10057 30073 10091 30107
rect 22293 30073 22327 30107
rect 45017 30073 45051 30107
rect 79517 30073 79551 30107
rect 86969 30073 87003 30107
rect 3985 30005 4019 30039
rect 4445 30005 4479 30039
rect 7757 30005 7791 30039
rect 11621 30005 11655 30039
rect 11897 30005 11931 30039
rect 15577 30005 15611 30039
rect 19993 30005 20027 30039
rect 22477 30005 22511 30039
rect 26801 30005 26835 30039
rect 28457 30005 28491 30039
rect 28733 30005 28767 30039
rect 28917 30005 28951 30039
rect 30849 30005 30883 30039
rect 37013 30005 37047 30039
rect 37933 30005 37967 30039
rect 48329 30005 48363 30039
rect 59185 30005 59219 30039
rect 59553 30005 59587 30039
rect 60013 30005 60047 30039
rect 66085 30005 66119 30039
rect 67465 30005 67499 30039
rect 68845 30005 68879 30039
rect 74457 30005 74491 30039
rect 81173 30005 81207 30039
rect 87061 30005 87095 30039
rect 15485 29801 15519 29835
rect 17969 29801 18003 29835
rect 19349 29801 19383 29835
rect 28181 29801 28215 29835
rect 36737 29801 36771 29835
rect 40969 29801 41003 29835
rect 42257 29801 42291 29835
rect 42625 29801 42659 29835
rect 53113 29801 53147 29835
rect 69397 29801 69431 29835
rect 73169 29801 73203 29835
rect 75193 29801 75227 29835
rect 79333 29801 79367 29835
rect 80621 29801 80655 29835
rect 6561 29733 6595 29767
rect 26801 29733 26835 29767
rect 28457 29733 28491 29767
rect 29285 29733 29319 29767
rect 29561 29733 29595 29767
rect 35449 29733 35483 29767
rect 45477 29733 45511 29767
rect 56425 29733 56459 29767
rect 56609 29733 56643 29767
rect 58265 29733 58299 29767
rect 61945 29733 61979 29767
rect 72893 29733 72927 29767
rect 4721 29665 4755 29699
rect 4997 29665 5031 29699
rect 9689 29665 9723 29699
rect 9965 29665 9999 29699
rect 11345 29665 11379 29699
rect 15301 29665 15335 29699
rect 18061 29665 18095 29699
rect 18153 29665 18187 29699
rect 19533 29665 19567 29699
rect 23857 29665 23891 29699
rect 26985 29665 27019 29699
rect 27169 29665 27203 29699
rect 27629 29665 27663 29699
rect 27721 29665 27755 29699
rect 28733 29665 28767 29699
rect 28825 29665 28859 29699
rect 29193 29665 29227 29699
rect 35265 29665 35299 29699
rect 36645 29665 36679 29699
rect 36921 29665 36955 29699
rect 41061 29665 41095 29699
rect 41245 29665 41279 29699
rect 41797 29665 41831 29699
rect 41981 29665 42015 29699
rect 44281 29665 44315 29699
rect 47041 29665 47075 29699
rect 48237 29665 48271 29699
rect 51273 29665 51307 29699
rect 51457 29665 51491 29699
rect 51641 29665 51675 29699
rect 52101 29665 52135 29699
rect 52653 29665 52687 29699
rect 52837 29665 52871 29699
rect 55137 29665 55171 29699
rect 55505 29665 55539 29699
rect 56793 29665 56827 29699
rect 56977 29665 57011 29699
rect 57161 29665 57195 29699
rect 57713 29665 57747 29699
rect 57897 29665 57931 29699
rect 58449 29665 58483 29699
rect 60473 29665 60507 29699
rect 67925 29665 67959 29699
rect 71237 29665 71271 29699
rect 71789 29665 71823 29699
rect 72341 29665 72375 29699
rect 72525 29665 72559 29699
rect 74089 29665 74123 29699
rect 79241 29665 79275 29699
rect 80529 29665 80563 29699
rect 19441 29597 19475 29631
rect 23489 29597 23523 29631
rect 23581 29597 23615 29631
rect 42717 29597 42751 29631
rect 47869 29597 47903 29631
rect 48053 29529 48087 29563
rect 51825 29597 51859 29631
rect 52009 29597 52043 29631
rect 53389 29597 53423 29631
rect 59461 29597 59495 29631
rect 60197 29597 60231 29631
rect 67649 29597 67683 29631
rect 71053 29597 71087 29631
rect 71421 29597 71455 29631
rect 71605 29597 71639 29631
rect 73813 29597 73847 29631
rect 75561 29597 75595 29631
rect 55321 29529 55355 29563
rect 59093 29529 59127 29563
rect 59553 29529 59587 29563
rect 71237 29529 71271 29563
rect 86877 29529 86911 29563
rect 87153 29529 87187 29563
rect 6101 29461 6135 29495
rect 9505 29461 9539 29495
rect 18337 29461 18371 29495
rect 19717 29461 19751 29495
rect 25145 29461 25179 29495
rect 35081 29461 35115 29495
rect 44097 29461 44131 29495
rect 45385 29461 45419 29495
rect 51273 29461 51307 29495
rect 58909 29461 58943 29495
rect 59185 29461 59219 29495
rect 59737 29461 59771 29495
rect 59921 29461 59955 29495
rect 61577 29461 61611 29495
rect 69029 29461 69063 29495
rect 86325 29461 86359 29495
rect 86509 29461 86543 29495
rect 86693 29461 86727 29495
rect 87245 29461 87279 29495
rect 87429 29461 87463 29495
rect 87613 29461 87647 29495
rect 4629 29257 4663 29291
rect 13185 29257 13219 29291
rect 21373 29189 21407 29223
rect 2789 29121 2823 29155
rect 3065 29121 3099 29155
rect 4169 29121 4203 29155
rect 12449 29121 12483 29155
rect 15393 29121 15427 29155
rect 20453 29121 20487 29155
rect 21189 29121 21223 29155
rect 12541 29053 12575 29087
rect 14565 29053 14599 29087
rect 20361 29053 20395 29087
rect 20565 29053 20599 29087
rect 23673 29053 23707 29087
rect 13001 28985 13035 29019
rect 14657 28985 14691 29019
rect 15025 28985 15059 29019
rect 21005 28985 21039 29019
rect 14841 28917 14875 28951
rect 14933 28917 14967 28951
rect 20177 28917 20211 28951
rect 23857 28917 23891 28951
rect 4537 28713 4571 28747
rect 13553 28713 13587 28747
rect 15393 28713 15427 28747
rect 4077 28577 4111 28611
rect 8217 28577 8251 28611
rect 9689 28577 9723 28611
rect 11253 28577 11287 28611
rect 8125 28441 8159 28475
rect 14013 28645 14047 28679
rect 15301 28645 15335 28679
rect 15853 28645 15887 28679
rect 15945 28645 15979 28679
rect 13829 28577 13863 28611
rect 13921 28577 13955 28611
rect 13645 28509 13679 28543
rect 14381 28509 14415 28543
rect 14565 28441 14599 28475
rect 15761 28577 15795 28611
rect 15577 28509 15611 28543
rect 16313 28509 16347 28543
rect 4261 28373 4295 28407
rect 8309 28373 8343 28407
rect 9873 28373 9907 28407
rect 11437 28373 11471 28407
rect 13553 28373 13587 28407
rect 15025 28373 15059 28407
rect 15301 28373 15335 28407
rect 9781 28169 9815 28203
rect 18429 28169 18463 28203
rect 20269 28169 20303 28203
rect 21189 28169 21223 28203
rect 24501 28169 24535 28203
rect 10057 28101 10091 28135
rect 15117 28101 15151 28135
rect 2605 28033 2639 28067
rect 2881 28033 2915 28067
rect 10701 28033 10735 28067
rect 15761 28033 15795 28067
rect 19901 28033 19935 28067
rect 20913 28033 20947 28067
rect 24777 28033 24811 28067
rect 25329 28033 25363 28067
rect 8125 27965 8159 27999
rect 9965 27965 9999 27999
rect 10241 27965 10275 27999
rect 14933 27965 14967 27999
rect 19165 27965 19199 27999
rect 19349 27965 19383 27999
rect 19441 27965 19475 27999
rect 19993 27965 20027 27999
rect 21005 27965 21039 27999
rect 25191 27965 25225 27999
rect 25605 27965 25639 27999
rect 25789 27965 25823 27999
rect 14197 27897 14231 27931
rect 14473 27897 14507 27931
rect 14565 27897 14599 27931
rect 15945 27897 15979 27931
rect 16129 27897 16163 27931
rect 16497 27897 16531 27931
rect 18613 27897 18647 27931
rect 20361 27897 20395 27931
rect 21649 27897 21683 27931
rect 3985 27829 4019 27863
rect 4445 27829 4479 27863
rect 8033 27829 8067 27863
rect 8309 27829 8343 27863
rect 14381 27829 14415 27863
rect 16037 27829 16071 27863
rect 13829 27625 13863 27659
rect 18245 27625 18279 27659
rect 22753 27625 22787 27659
rect 8769 27557 8803 27591
rect 14013 27557 14047 27591
rect 25697 27557 25731 27591
rect 6929 27489 6963 27523
rect 8033 27489 8067 27523
rect 8309 27489 8343 27523
rect 9689 27489 9723 27523
rect 9965 27489 9999 27523
rect 11253 27489 11287 27523
rect 12541 27489 12575 27523
rect 13645 27489 13679 27523
rect 13921 27489 13955 27523
rect 15393 27489 15427 27523
rect 18981 27489 19015 27523
rect 19165 27489 19199 27523
rect 19257 27489 19291 27523
rect 19901 27489 19935 27523
rect 22575 27489 22609 27523
rect 24225 27489 24259 27523
rect 24961 27489 24995 27523
rect 25329 27489 25363 27523
rect 25513 27489 25547 27523
rect 26709 27489 26743 27523
rect 27261 27489 27295 27523
rect 27445 27489 27479 27523
rect 10425 27421 10459 27455
rect 14381 27421 14415 27455
rect 15301 27421 15335 27455
rect 15853 27421 15887 27455
rect 18429 27421 18463 27455
rect 19717 27421 19751 27455
rect 24317 27421 24351 27455
rect 25053 27421 25087 27455
rect 26525 27421 26559 27455
rect 7941 27353 7975 27387
rect 8125 27353 8159 27387
rect 9781 27353 9815 27387
rect 20085 27353 20119 27387
rect 7113 27285 7147 27319
rect 11437 27285 11471 27319
rect 12725 27285 12759 27319
rect 20177 27285 20211 27319
rect 25881 27285 25915 27319
rect 26249 27285 26283 27319
rect 27721 27285 27755 27319
rect 4721 27081 4755 27115
rect 7297 27081 7331 27115
rect 23857 27081 23891 27115
rect 8309 27013 8343 27047
rect 9965 27013 9999 27047
rect 14105 27013 14139 27047
rect 26341 27013 26375 27047
rect 8953 26945 8987 26979
rect 3985 26877 4019 26911
rect 7113 26877 7147 26911
rect 7205 26877 7239 26911
rect 8217 26877 8251 26911
rect 8493 26877 8527 26911
rect 9873 26877 9907 26911
rect 10149 26877 10183 26911
rect 15301 26945 15335 26979
rect 26525 26945 26559 26979
rect 26801 26945 26835 26979
rect 14749 26877 14783 26911
rect 14841 26877 14875 26911
rect 15025 26877 15059 26911
rect 15669 26877 15703 26911
rect 23673 26877 23707 26911
rect 24777 26877 24811 26911
rect 3801 26809 3835 26843
rect 4353 26809 4387 26843
rect 10609 26809 10643 26843
rect 14105 26809 14139 26843
rect 14197 26809 14231 26843
rect 4537 26741 4571 26775
rect 7941 26741 7975 26775
rect 8033 26741 8067 26775
rect 24961 26741 24995 26775
rect 28089 26741 28123 26775
rect 6561 26537 6595 26571
rect 8401 26537 8435 26571
rect 9781 26537 9815 26571
rect 24225 26537 24259 26571
rect 28089 26537 28123 26571
rect 4261 26469 4295 26503
rect 5641 26469 5675 26503
rect 6377 26469 6411 26503
rect 24133 26469 24167 26503
rect 4169 26401 4203 26435
rect 4353 26401 4387 26435
rect 5825 26401 5859 26435
rect 8217 26401 8251 26435
rect 9689 26401 9723 26435
rect 9965 26401 9999 26435
rect 10701 26401 10735 26435
rect 17325 26401 17359 26435
rect 18613 26401 18647 26435
rect 22661 26401 22695 26435
rect 23397 26401 23431 26435
rect 23765 26401 23799 26435
rect 23949 26401 23983 26435
rect 24777 26401 24811 26435
rect 27997 26401 28031 26435
rect 4813 26333 4847 26367
rect 6101 26333 6135 26367
rect 17141 26333 17175 26367
rect 17233 26333 17267 26367
rect 18760 26333 18794 26367
rect 18981 26333 19015 26367
rect 22753 26333 22787 26367
rect 23489 26333 23523 26367
rect 24501 26333 24535 26367
rect 4997 26265 5031 26299
rect 10885 26265 10919 26299
rect 18889 26265 18923 26299
rect 24869 26265 24903 26299
rect 28365 26265 28399 26299
rect 5181 26197 5215 26231
rect 8033 26197 8067 26231
rect 17509 26197 17543 26231
rect 19073 26197 19107 26231
rect 8309 25993 8343 26027
rect 15945 25993 15979 26027
rect 18429 25993 18463 26027
rect 18797 25993 18831 26027
rect 14933 25925 14967 25959
rect 2881 25857 2915 25891
rect 18521 25857 18555 25891
rect 2605 25789 2639 25823
rect 8125 25789 8159 25823
rect 15117 25789 15151 25823
rect 16129 25789 16163 25823
rect 18613 25789 18647 25823
rect 3985 25653 4019 25687
rect 4445 25653 4479 25687
rect 7941 25653 7975 25687
rect 15209 25653 15243 25687
rect 16221 25653 16255 25687
rect 13093 25449 13127 25483
rect 21649 25449 21683 25483
rect 23121 25449 23155 25483
rect 24133 25449 24167 25483
rect 15301 25381 15335 25415
rect 25697 25381 25731 25415
rect 5641 25313 5675 25347
rect 7389 25313 7423 25347
rect 11161 25313 11195 25347
rect 11713 25313 11747 25347
rect 11897 25313 11931 25347
rect 13185 25313 13219 25347
rect 15945 25313 15979 25347
rect 16313 25313 16347 25347
rect 16497 25313 16531 25347
rect 18981 25313 19015 25347
rect 19211 25313 19245 25347
rect 22385 25313 22419 25347
rect 22753 25313 22787 25347
rect 22937 25313 22971 25347
rect 24409 25313 24443 25347
rect 24961 25313 24995 25347
rect 25145 25313 25179 25347
rect 26525 25313 26559 25347
rect 5917 25245 5951 25279
rect 10885 25245 10919 25279
rect 11069 25245 11103 25279
rect 15853 25245 15887 25279
rect 19349 25245 19383 25279
rect 21741 25245 21775 25279
rect 22477 25245 22511 25279
rect 23213 25245 23247 25279
rect 24317 25245 24351 25279
rect 12081 25177 12115 25211
rect 19146 25177 19180 25211
rect 7205 25109 7239 25143
rect 12541 25109 12575 25143
rect 12725 25109 12759 25143
rect 13369 25109 13403 25143
rect 19625 25109 19659 25143
rect 25421 25109 25455 25143
rect 26709 25109 26743 25143
rect 24317 24905 24351 24939
rect 7205 24837 7239 24871
rect 19073 24837 19107 24871
rect 6101 24769 6135 24803
rect 25513 24769 25547 24803
rect 5181 24701 5215 24735
rect 5365 24701 5399 24735
rect 5457 24701 5491 24735
rect 6837 24701 6871 24735
rect 12633 24701 12667 24735
rect 12817 24701 12851 24735
rect 13369 24701 13403 24735
rect 13645 24701 13679 24735
rect 18061 24701 18095 24735
rect 18429 24701 18463 24735
rect 18797 24701 18831 24735
rect 19073 24701 19107 24735
rect 20269 24701 20303 24735
rect 24133 24701 24167 24735
rect 25145 24701 25179 24735
rect 25237 24701 25271 24735
rect 5917 24633 5951 24667
rect 13921 24633 13955 24667
rect 26893 24633 26927 24667
rect 5089 24565 5123 24599
rect 6929 24565 6963 24599
rect 20361 24565 20395 24599
rect 6193 24361 6227 24395
rect 26617 24361 26651 24395
rect 18705 24293 18739 24327
rect 24685 24293 24719 24327
rect 5181 24225 5215 24259
rect 5733 24225 5767 24259
rect 5917 24225 5951 24259
rect 11529 24225 11563 24259
rect 18245 24225 18279 24259
rect 23121 24225 23155 24259
rect 23213 24225 23247 24259
rect 23397 24225 23431 24259
rect 23857 24225 23891 24259
rect 23949 24225 23983 24259
rect 24869 24225 24903 24259
rect 26525 24225 26559 24259
rect 4997 24157 5031 24191
rect 11253 24157 11287 24191
rect 18153 24157 18187 24191
rect 24317 24089 24351 24123
rect 4813 24021 4847 24055
rect 11161 24021 11195 24055
rect 12817 24021 12851 24055
rect 26893 24021 26927 24055
rect 28917 24021 28951 24055
rect 12909 23749 12943 23783
rect 4261 23681 4295 23715
rect 6009 23681 6043 23715
rect 15209 23681 15243 23715
rect 19441 23681 19475 23715
rect 25789 23681 25823 23715
rect 4537 23613 4571 23647
rect 5917 23613 5951 23647
rect 6837 23613 6871 23647
rect 12817 23613 12851 23647
rect 13921 23613 13955 23647
rect 14289 23613 14323 23647
rect 14473 23613 14507 23647
rect 14749 23613 14783 23647
rect 14933 23613 14967 23647
rect 18889 23613 18923 23647
rect 18981 23613 19015 23647
rect 24133 23613 24167 23647
rect 24409 23613 24443 23647
rect 7205 23545 7239 23579
rect 13829 23545 13863 23579
rect 6929 23477 6963 23511
rect 12725 23477 12759 23511
rect 18705 23477 18739 23511
rect 24041 23477 24075 23511
rect 12817 23273 12851 23307
rect 22661 23273 22695 23307
rect 24777 23273 24811 23307
rect 9505 23205 9539 23239
rect 26617 23205 26651 23239
rect 4522 23137 4556 23171
rect 5089 23137 5123 23171
rect 5273 23137 5307 23171
rect 4353 23069 4387 23103
rect 5549 23069 5583 23103
rect 13553 23137 13587 23171
rect 13829 23137 13863 23171
rect 14105 23137 14139 23171
rect 17693 23137 17727 23171
rect 22569 23137 22603 23171
rect 22937 23137 22971 23171
rect 23765 23137 23799 23171
rect 24317 23137 24351 23171
rect 24501 23137 24535 23171
rect 26525 23137 26559 23171
rect 13185 23069 13219 23103
rect 23397 23069 23431 23103
rect 23581 23069 23615 23103
rect 4261 22933 4295 22967
rect 9505 22933 9539 22967
rect 17877 22933 17911 22967
rect 8861 22729 8895 22763
rect 17877 22729 17911 22763
rect 20637 22729 20671 22763
rect 15117 22661 15151 22695
rect 2605 22593 2639 22627
rect 2789 22593 2823 22627
rect 13645 22593 13679 22627
rect 18245 22593 18279 22627
rect 23397 22593 23431 22627
rect 2881 22525 2915 22559
rect 3433 22525 3467 22559
rect 3617 22525 3651 22559
rect 8493 22525 8527 22559
rect 13737 22525 13771 22559
rect 14105 22525 14139 22559
rect 14289 22525 14323 22559
rect 14565 22525 14599 22559
rect 14749 22525 14783 22559
rect 18613 22525 18647 22559
rect 18797 22525 18831 22559
rect 18981 22525 19015 22559
rect 19165 22525 19199 22559
rect 20545 22525 20579 22559
rect 23949 22525 23983 22559
rect 24041 22525 24075 22559
rect 24501 22525 24535 22559
rect 24685 22525 24719 22559
rect 25973 22525 26007 22559
rect 19717 22457 19751 22491
rect 26065 22457 26099 22491
rect 3893 22389 3927 22423
rect 8585 22389 8619 22423
rect 18153 22389 18187 22423
rect 24961 22389 24995 22423
rect 8033 22185 8067 22219
rect 13093 22185 13127 22219
rect 12909 22117 12943 22151
rect 13737 22117 13771 22151
rect 4077 22049 4111 22083
rect 4169 22049 4203 22083
rect 7021 22049 7055 22083
rect 7573 22049 7607 22083
rect 7757 22049 7791 22083
rect 11621 22049 11655 22083
rect 12173 22049 12207 22083
rect 12357 22049 12391 22083
rect 13645 22049 13679 22083
rect 15577 22049 15611 22083
rect 18337 22049 18371 22083
rect 18705 22049 18739 22083
rect 18889 22049 18923 22083
rect 19165 22049 19199 22083
rect 19257 22049 19291 22083
rect 24133 22049 24167 22083
rect 6837 21981 6871 22015
rect 11437 21981 11471 22015
rect 23857 21981 23891 22015
rect 18061 21913 18095 21947
rect 4445 21845 4479 21879
rect 6653 21845 6687 21879
rect 11253 21845 11287 21879
rect 12633 21845 12667 21879
rect 14013 21845 14047 21879
rect 15761 21845 15795 21879
rect 18153 21845 18187 21879
rect 19717 21845 19751 21879
rect 23765 21845 23799 21879
rect 25421 21845 25455 21879
rect 5825 21641 5859 21675
rect 9321 21641 9355 21675
rect 25973 21641 26007 21675
rect 4353 21573 4387 21607
rect 3065 21505 3099 21539
rect 7757 21505 7791 21539
rect 8033 21505 8067 21539
rect 12725 21505 12759 21539
rect 24685 21505 24719 21539
rect 2789 21437 2823 21471
rect 5641 21437 5675 21471
rect 9505 21437 9539 21471
rect 12173 21437 12207 21471
rect 12449 21437 12483 21471
rect 15669 21437 15703 21471
rect 24409 21437 24443 21471
rect 14105 21369 14139 21403
rect 4629 21301 4663 21335
rect 15761 21301 15795 21335
rect 24225 21301 24259 21335
rect 23673 21029 23707 21063
rect 22017 20893 22051 20927
rect 22293 20893 22327 20927
rect 23857 20757 23891 20791
rect 4445 20553 4479 20587
rect 16313 20553 16347 20587
rect 16589 20553 16623 20587
rect 23857 20553 23891 20587
rect 3985 20485 4019 20519
rect 2881 20417 2915 20451
rect 14749 20417 14783 20451
rect 18429 20417 18463 20451
rect 2605 20349 2639 20383
rect 6837 20349 6871 20383
rect 8125 20349 8159 20383
rect 10609 20349 10643 20383
rect 15117 20349 15151 20383
rect 15301 20349 15335 20383
rect 15577 20349 15611 20383
rect 15669 20349 15703 20383
rect 18061 20349 18095 20383
rect 22569 20349 22603 20383
rect 23679 20349 23713 20383
rect 26341 20349 26375 20383
rect 4629 20213 4663 20247
rect 7021 20213 7055 20247
rect 8309 20213 8343 20247
rect 10793 20213 10827 20247
rect 14657 20213 14691 20247
rect 16129 20213 16163 20247
rect 18153 20213 18187 20247
rect 22661 20213 22695 20247
rect 24041 20213 24075 20247
rect 26433 20213 26467 20247
rect 17969 20009 18003 20043
rect 20453 20009 20487 20043
rect 21373 20009 21407 20043
rect 22661 20009 22695 20043
rect 5365 19873 5399 19907
rect 5917 19873 5951 19907
rect 6101 19873 6135 19907
rect 11437 19873 11471 19907
rect 11989 19873 12023 19907
rect 12173 19873 12207 19907
rect 20361 19873 20395 19907
rect 21465 19873 21499 19907
rect 21649 19873 21683 19907
rect 22201 19873 22235 19907
rect 22385 19873 22419 19907
rect 24869 19873 24903 19907
rect 26525 19873 26559 19907
rect 5181 19805 5215 19839
rect 11253 19805 11287 19839
rect 16589 19805 16623 19839
rect 16865 19805 16899 19839
rect 6285 19737 6319 19771
rect 16405 19737 16439 19771
rect 4997 19669 5031 19703
rect 11161 19669 11195 19703
rect 12449 19669 12483 19703
rect 20177 19669 20211 19703
rect 25053 19669 25087 19703
rect 26617 19669 26651 19703
rect 26985 19465 27019 19499
rect 13001 19397 13035 19431
rect 9413 19329 9447 19363
rect 6837 19261 6871 19295
rect 6929 19261 6963 19295
rect 8125 19261 8159 19295
rect 8309 19261 8343 19295
rect 8861 19261 8895 19295
rect 9045 19261 9079 19295
rect 10333 19261 10367 19295
rect 12817 19261 12851 19295
rect 12909 19261 12943 19295
rect 16773 19261 16807 19295
rect 16865 19261 16899 19295
rect 25421 19261 25455 19295
rect 25605 19261 25639 19295
rect 25881 19261 25915 19295
rect 10425 19193 10459 19227
rect 7205 19125 7239 19159
rect 7941 19125 7975 19159
rect 10701 19125 10735 19159
rect 12817 19125 12851 19159
rect 13277 19125 13311 19159
rect 17049 19125 17083 19159
rect 6285 18921 6319 18955
rect 16221 18921 16255 18955
rect 17509 18921 17543 18955
rect 20361 18921 20395 18955
rect 23949 18921 23983 18955
rect 24041 18921 24075 18955
rect 26249 18921 26283 18955
rect 27721 18921 27755 18955
rect 4997 18785 5031 18819
rect 9965 18785 9999 18819
rect 12449 18785 12483 18819
rect 16313 18785 16347 18819
rect 16497 18785 16531 18819
rect 17049 18785 17083 18819
rect 17233 18785 17267 18819
rect 19441 18785 19475 18819
rect 19809 18785 19843 18819
rect 19993 18785 20027 18819
rect 23949 18785 23983 18819
rect 24225 18785 24259 18819
rect 24409 18785 24443 18819
rect 24961 18785 24995 18819
rect 25145 18785 25179 18819
rect 26709 18785 26743 18819
rect 26801 18785 26835 18819
rect 27169 18785 27203 18819
rect 27261 18785 27295 18819
rect 4721 18717 4755 18751
rect 6469 18717 6503 18751
rect 9689 18717 9723 18751
rect 11437 18717 11471 18751
rect 11989 18717 12023 18751
rect 12173 18717 12207 18751
rect 18797 18717 18831 18751
rect 19349 18717 19383 18751
rect 20177 18717 20211 18751
rect 25329 18649 25363 18683
rect 11253 18581 11287 18615
rect 13737 18581 13771 18615
rect 4445 18377 4479 18411
rect 20269 18377 20303 18411
rect 26249 18377 26283 18411
rect 2605 18241 2639 18275
rect 2881 18241 2915 18275
rect 25145 18241 25179 18275
rect 9873 18173 9907 18207
rect 14197 18173 14231 18207
rect 19165 18173 19199 18207
rect 19349 18173 19383 18207
rect 19717 18173 19751 18207
rect 19901 18173 19935 18207
rect 24869 18173 24903 18207
rect 18705 18105 18739 18139
rect 20085 18105 20119 18139
rect 4169 18037 4203 18071
rect 4629 18037 4663 18071
rect 9689 18037 9723 18071
rect 14289 18037 14323 18071
rect 24777 18037 24811 18071
rect 20085 17833 20119 17867
rect 20269 17833 20303 17867
rect 21005 17765 21039 17799
rect 7849 17697 7883 17731
rect 14105 17697 14139 17731
rect 18429 17697 18463 17731
rect 18705 17697 18739 17731
rect 19257 17697 19291 17731
rect 19441 17697 19475 17731
rect 20913 17697 20947 17731
rect 27997 17697 28031 17731
rect 13553 17629 13587 17663
rect 18613 17629 18647 17663
rect 14197 17561 14231 17595
rect 19625 17561 19659 17595
rect 7941 17493 7975 17527
rect 8217 17493 8251 17527
rect 21189 17493 21223 17527
rect 28089 17493 28123 17527
rect 4445 17289 4479 17323
rect 13185 17289 13219 17323
rect 15301 17289 15335 17323
rect 2605 17153 2639 17187
rect 2881 17153 2915 17187
rect 13461 17153 13495 17187
rect 19441 17153 19475 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 7573 17085 7607 17119
rect 7757 17085 7791 17119
rect 13369 17085 13403 17119
rect 13737 17085 13771 17119
rect 14013 17085 14047 17119
rect 14197 17085 14231 17119
rect 14381 17085 14415 17119
rect 15117 17085 15151 17119
rect 19165 17085 19199 17119
rect 26617 17085 26651 17119
rect 27169 17085 27203 17119
rect 27353 17085 27387 17119
rect 6561 17017 6595 17051
rect 13093 17017 13127 17051
rect 20821 17017 20855 17051
rect 4169 16949 4203 16983
rect 4629 16949 4663 16983
rect 8033 16949 8067 16983
rect 14841 16949 14875 16983
rect 21005 16949 21039 16983
rect 27629 16949 27663 16983
rect 8585 16745 8619 16779
rect 20177 16745 20211 16779
rect 20269 16745 20303 16779
rect 23673 16745 23707 16779
rect 26249 16745 26283 16779
rect 28089 16745 28123 16779
rect 12357 16677 12391 16711
rect 7021 16609 7055 16643
rect 7297 16609 7331 16643
rect 12449 16609 12483 16643
rect 13093 16609 13127 16643
rect 13185 16609 13219 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 18429 16609 18463 16643
rect 18613 16609 18647 16643
rect 18797 16609 18831 16643
rect 19349 16609 19383 16643
rect 19533 16609 19567 16643
rect 23857 16609 23891 16643
rect 26525 16609 26559 16643
rect 26801 16609 26835 16643
rect 8769 16541 8803 16575
rect 19809 16405 19843 16439
rect 4445 16201 4479 16235
rect 8953 16201 8987 16235
rect 9597 16201 9631 16235
rect 14841 16201 14875 16235
rect 23673 16201 23707 16235
rect 24869 16201 24903 16235
rect 26525 16201 26559 16235
rect 2881 16065 2915 16099
rect 7205 16065 7239 16099
rect 8861 16065 8895 16099
rect 13277 16065 13311 16099
rect 19901 16065 19935 16099
rect 24961 16065 24995 16099
rect 2605 15997 2639 16031
rect 4537 15997 4571 16031
rect 7481 15997 7515 16031
rect 9689 15997 9723 16031
rect 13001 15997 13035 16031
rect 19625 15997 19659 16031
rect 23857 15997 23891 16031
rect 25237 15997 25271 16031
rect 21281 15929 21315 15963
rect 4169 15861 4203 15895
rect 9781 15861 9815 15895
rect 12817 15861 12851 15895
rect 14381 15861 14415 15895
rect 21465 15861 21499 15895
rect 24041 15861 24075 15895
rect 7665 15657 7699 15691
rect 21005 15657 21039 15691
rect 21281 15657 21315 15691
rect 25421 15657 25455 15691
rect 26617 15589 26651 15623
rect 6653 15521 6687 15555
rect 7205 15521 7239 15555
rect 7389 15521 7423 15555
rect 20913 15521 20947 15555
rect 24409 15521 24443 15555
rect 24961 15521 24995 15555
rect 25145 15521 25179 15555
rect 26525 15521 26559 15555
rect 6561 15453 6595 15487
rect 24041 15453 24075 15487
rect 24225 15453 24259 15487
rect 6377 15385 6411 15419
rect 4537 15113 4571 15147
rect 2973 14977 3007 15011
rect 13829 14977 13863 15011
rect 2697 14909 2731 14943
rect 13553 14909 13587 14943
rect 4077 14773 4111 14807
rect 4629 14773 4663 14807
rect 13369 14773 13403 14807
rect 15117 14773 15151 14807
rect 21741 14569 21775 14603
rect 14381 14501 14415 14535
rect 18061 14501 18095 14535
rect 8309 14433 8343 14467
rect 16405 14433 16439 14467
rect 18153 14433 18187 14467
rect 20913 14433 20947 14467
rect 8217 14365 8251 14399
rect 12725 14365 12759 14399
rect 13001 14365 13035 14399
rect 16681 14365 16715 14399
rect 8493 14229 8527 14263
rect 12633 14229 12667 14263
rect 21557 14229 21591 14263
rect 4629 14025 4663 14059
rect 7205 14025 7239 14059
rect 8953 14025 8987 14059
rect 10609 14025 10643 14059
rect 20729 14025 20763 14059
rect 25421 14025 25455 14059
rect 2605 13889 2639 13923
rect 2881 13889 2915 13923
rect 4445 13889 4479 13923
rect 12725 13889 12759 13923
rect 14013 13889 14047 13923
rect 14565 13889 14599 13923
rect 20913 13889 20947 13923
rect 25605 13889 25639 13923
rect 27905 13889 27939 13923
rect 7389 13821 7423 13855
rect 8309 13821 8343 13855
rect 8493 13821 8527 13855
rect 8769 13821 8803 13855
rect 9321 13821 9355 13855
rect 10793 13821 10827 13855
rect 12449 13821 12483 13855
rect 12541 13821 12575 13855
rect 14657 13821 14691 13855
rect 15025 13821 15059 13855
rect 15209 13821 15243 13855
rect 21189 13821 21223 13855
rect 25789 13821 25823 13855
rect 26341 13821 26375 13855
rect 26525 13821 26559 13855
rect 27813 13821 27847 13855
rect 8677 13753 8711 13787
rect 3985 13685 4019 13719
rect 7573 13685 7607 13719
rect 15393 13685 15427 13719
rect 22293 13685 22327 13719
rect 26801 13685 26835 13719
rect 6469 13481 6503 13515
rect 7573 13481 7607 13515
rect 10517 13481 10551 13515
rect 23489 13481 23523 13515
rect 26249 13481 26283 13515
rect 6837 13413 6871 13447
rect 17049 13413 17083 13447
rect 6653 13345 6687 13379
rect 6929 13345 6963 13379
rect 8309 13345 8343 13379
rect 8861 13345 8895 13379
rect 9873 13345 9907 13379
rect 17693 13345 17727 13379
rect 18061 13345 18095 13379
rect 21925 13345 21959 13379
rect 26525 13345 26559 13379
rect 26801 13345 26835 13379
rect 8217 13277 8251 13311
rect 9781 13277 9815 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 21649 13277 21683 13311
rect 23029 13277 23063 13311
rect 7113 13141 7147 13175
rect 8493 13141 8527 13175
rect 10057 13141 10091 13175
rect 18429 13141 18463 13175
rect 28089 13141 28123 13175
rect 4445 12937 4479 12971
rect 8677 12937 8711 12971
rect 9137 12937 9171 12971
rect 10425 12937 10459 12971
rect 15485 12937 15519 12971
rect 15761 12937 15795 12971
rect 24317 12937 24351 12971
rect 8217 12869 8251 12903
rect 2605 12801 2639 12835
rect 2881 12801 2915 12835
rect 24501 12801 24535 12835
rect 8493 12733 8527 12767
rect 10701 12733 10735 12767
rect 15393 12733 15427 12767
rect 24777 12733 24811 12767
rect 8401 12665 8435 12699
rect 10609 12665 10643 12699
rect 11161 12665 11195 12699
rect 4169 12597 4203 12631
rect 25881 12597 25915 12631
rect 7297 12393 7331 12427
rect 10609 12393 10643 12427
rect 11989 12393 12023 12427
rect 22661 12393 22695 12427
rect 22845 12393 22879 12427
rect 10333 12325 10367 12359
rect 11713 12325 11747 12359
rect 7021 12257 7055 12291
rect 7205 12257 7239 12291
rect 10517 12257 10551 12291
rect 11897 12257 11931 12291
rect 18981 12257 19015 12291
rect 23029 12257 23063 12291
rect 17233 12189 17267 12223
rect 17509 12189 17543 12223
rect 18889 12189 18923 12223
rect 8493 11849 8527 11883
rect 13829 11849 13863 11883
rect 19441 11849 19475 11883
rect 25053 11849 25087 11883
rect 2605 11713 2639 11747
rect 2881 11713 2915 11747
rect 12449 11713 12483 11747
rect 14197 11713 14231 11747
rect 18061 11713 18095 11747
rect 21005 11713 21039 11747
rect 25237 11713 25271 11747
rect 25513 11713 25547 11747
rect 8217 11645 8251 11679
rect 8401 11645 8435 11679
rect 12725 11645 12759 11679
rect 16865 11645 16899 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 19027 11645 19061 11679
rect 19165 11645 19199 11679
rect 4169 11509 4203 11543
rect 4445 11509 4479 11543
rect 17049 11509 17083 11543
rect 21649 11509 21683 11543
rect 26617 11509 26651 11543
rect 13185 11237 13219 11271
rect 5641 11169 5675 11203
rect 13829 11169 13863 11203
rect 14197 11169 14231 11203
rect 14289 11169 14323 11203
rect 14565 11169 14599 11203
rect 15945 11169 15979 11203
rect 16313 11169 16347 11203
rect 5917 11101 5951 11135
rect 7297 11101 7331 11135
rect 13921 11101 13955 11135
rect 7389 11033 7423 11067
rect 16129 11033 16163 11067
rect 8769 10761 8803 10795
rect 9229 10761 9263 10795
rect 22017 10761 22051 10795
rect 4445 10693 4479 10727
rect 2605 10625 2639 10659
rect 2881 10625 2915 10659
rect 14289 10625 14323 10659
rect 26065 10625 26099 10659
rect 7389 10557 7423 10591
rect 7665 10557 7699 10591
rect 14197 10557 14231 10591
rect 14565 10557 14599 10591
rect 14749 10557 14783 10591
rect 20637 10557 20671 10591
rect 20913 10557 20947 10591
rect 25789 10557 25823 10591
rect 13553 10489 13587 10523
rect 4169 10421 4203 10455
rect 20453 10421 20487 10455
rect 25605 10421 25639 10455
rect 27169 10421 27203 10455
rect 7665 10217 7699 10251
rect 12633 10217 12667 10251
rect 14105 10217 14139 10251
rect 22293 10217 22327 10251
rect 27905 10217 27939 10251
rect 8217 10081 8251 10115
rect 8585 10081 8619 10115
rect 12725 10081 12759 10115
rect 13001 10081 13035 10115
rect 19901 10081 19935 10115
rect 21189 10081 21223 10115
rect 26801 10081 26835 10115
rect 8125 10013 8159 10047
rect 8493 10013 8527 10047
rect 20913 10013 20947 10047
rect 26341 10013 26375 10047
rect 26525 10013 26559 10047
rect 19717 9877 19751 9911
rect 20637 9877 20671 9911
rect 15301 9673 15335 9707
rect 19441 9605 19475 9639
rect 6929 9537 6963 9571
rect 7573 9537 7607 9571
rect 13737 9537 13771 9571
rect 15485 9537 15519 9571
rect 18521 9537 18555 9571
rect 21281 9537 21315 9571
rect 7481 9469 7515 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 14013 9469 14047 9503
rect 18705 9469 18739 9503
rect 19073 9469 19107 9503
rect 19165 9469 19199 9503
rect 18061 9401 18095 9435
rect 21925 9333 21959 9367
rect 6561 9129 6595 9163
rect 6837 9061 6871 9095
rect 19441 9061 19475 9095
rect 4997 8993 5031 9027
rect 17785 8993 17819 9027
rect 18061 8993 18095 9027
rect 5273 8925 5307 8959
rect 19533 8925 19567 8959
rect 21741 8925 21775 8959
rect 21925 8925 21959 8959
rect 22201 8925 22235 8959
rect 23489 8789 23523 8823
rect 4445 8585 4479 8619
rect 9873 8585 9907 8619
rect 12633 8585 12667 8619
rect 14197 8585 14231 8619
rect 25053 8585 25087 8619
rect 2605 8449 2639 8483
rect 2881 8449 2915 8483
rect 8493 8449 8527 8483
rect 10241 8449 10275 8483
rect 13093 8449 13127 8483
rect 21465 8449 21499 8483
rect 23949 8449 23983 8483
rect 8769 8381 8803 8415
rect 12817 8381 12851 8415
rect 20821 8381 20855 8415
rect 23489 8381 23523 8415
rect 23673 8381 23707 8415
rect 3985 8245 4019 8279
rect 5641 8041 5675 8075
rect 5917 8041 5951 8075
rect 4077 7905 4111 7939
rect 8033 7905 8067 7939
rect 4353 7837 4387 7871
rect 8677 7837 8711 7871
rect 4353 7497 4387 7531
rect 9229 7497 9263 7531
rect 9689 7497 9723 7531
rect 15209 7497 15243 7531
rect 2605 7361 2639 7395
rect 2881 7361 2915 7395
rect 7849 7361 7883 7395
rect 8125 7293 8159 7327
rect 10793 7293 10827 7327
rect 13645 7293 13679 7327
rect 13921 7293 13955 7327
rect 13461 7225 13495 7259
rect 4169 7157 4203 7191
rect 11437 7157 11471 7191
rect 13921 6885 13955 6919
rect 8033 6817 8067 6851
rect 8677 6817 8711 6851
rect 12081 6817 12115 6851
rect 12265 6817 12299 6851
rect 12541 6817 12575 6851
rect 4905 6409 4939 6443
rect 3157 6273 3191 6307
rect 3433 6273 3467 6307
rect 4537 6069 4571 6103
rect 26341 5321 26375 5355
rect 26065 5253 26099 5287
rect 26709 5185 26743 5219
rect 26433 5117 26467 5151
rect 28089 5049 28123 5083
rect 11529 4777 11563 4811
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 11069 4437 11103 4471
rect 3893 4097 3927 4131
rect 5457 4097 5491 4131
rect 3617 4029 3651 4063
rect 5549 4029 5583 4063
rect 4997 3893 5031 3927
rect 4721 3145 4755 3179
rect 3249 3009 3283 3043
rect 2973 2941 3007 2975
rect 4905 2941 4939 2975
rect 4353 2805 4387 2839
<< metal1 >>
rect 4062 48356 4068 48408
rect 4120 48396 4126 48408
rect 14918 48396 14924 48408
rect 4120 48368 14924 48396
rect 4120 48356 4126 48368
rect 14918 48356 14924 48368
rect 14976 48356 14982 48408
rect 3970 48288 3976 48340
rect 4028 48328 4034 48340
rect 73062 48328 73068 48340
rect 4028 48300 73068 48328
rect 4028 48288 4034 48300
rect 73062 48288 73068 48300
rect 73120 48288 73126 48340
rect 1104 47898 108008 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 65686 47898
rect 65738 47846 65750 47898
rect 65802 47846 65814 47898
rect 65866 47846 65878 47898
rect 65930 47846 96406 47898
rect 96458 47846 96470 47898
rect 96522 47846 96534 47898
rect 96586 47846 96598 47898
rect 96650 47846 108008 47898
rect 1104 47824 108008 47846
rect 8386 47648 8392 47660
rect 8347 47620 8392 47648
rect 8386 47608 8392 47620
rect 8444 47608 8450 47660
rect 7926 47580 7932 47592
rect 7887 47552 7932 47580
rect 7926 47540 7932 47552
rect 7984 47540 7990 47592
rect 8481 47583 8539 47589
rect 8481 47549 8493 47583
rect 8527 47580 8539 47583
rect 13722 47580 13728 47592
rect 8527 47552 13728 47580
rect 8527 47549 8539 47552
rect 8481 47543 8539 47549
rect 13722 47540 13728 47552
rect 13780 47540 13786 47592
rect 12066 47404 12072 47456
rect 12124 47444 12130 47456
rect 22462 47444 22468 47456
rect 12124 47416 22468 47444
rect 12124 47404 12130 47416
rect 22462 47404 22468 47416
rect 22520 47404 22526 47456
rect 1104 47354 108008 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 50326 47354
rect 50378 47302 50390 47354
rect 50442 47302 50454 47354
rect 50506 47302 50518 47354
rect 50570 47302 81046 47354
rect 81098 47302 81110 47354
rect 81162 47302 81174 47354
rect 81226 47302 81238 47354
rect 81290 47302 108008 47354
rect 1104 47280 108008 47302
rect 7745 47243 7803 47249
rect 7745 47240 7757 47243
rect 5184 47212 7757 47240
rect 3418 47064 3424 47116
rect 3476 47104 3482 47116
rect 4525 47107 4583 47113
rect 3476 47076 4384 47104
rect 3476 47064 3482 47076
rect 4249 47039 4307 47045
rect 4249 47005 4261 47039
rect 4295 47005 4307 47039
rect 4356 47036 4384 47076
rect 4525 47073 4537 47107
rect 4571 47104 4583 47107
rect 5184 47104 5212 47212
rect 7745 47209 7757 47212
rect 7791 47209 7803 47243
rect 22278 47240 22284 47252
rect 7745 47203 7803 47209
rect 12084 47212 22284 47240
rect 7926 47104 7932 47116
rect 4571 47076 5212 47104
rect 7887 47076 7932 47104
rect 4571 47073 4583 47076
rect 4525 47067 4583 47073
rect 7926 47064 7932 47076
rect 7984 47064 7990 47116
rect 8205 47107 8263 47113
rect 8205 47073 8217 47107
rect 8251 47104 8263 47107
rect 8573 47107 8631 47113
rect 8573 47104 8585 47107
rect 8251 47076 8585 47104
rect 8251 47073 8263 47076
rect 8205 47067 8263 47073
rect 8573 47073 8585 47076
rect 8619 47104 8631 47107
rect 12084 47104 12112 47212
rect 22278 47200 22284 47212
rect 22336 47200 22342 47252
rect 22462 47240 22468 47252
rect 22423 47212 22468 47240
rect 22462 47200 22468 47212
rect 22520 47200 22526 47252
rect 13004 47144 13952 47172
rect 13004 47113 13032 47144
rect 8619 47076 12112 47104
rect 12437 47107 12495 47113
rect 8619 47073 8631 47076
rect 8573 47067 8631 47073
rect 12437 47073 12449 47107
rect 12483 47104 12495 47107
rect 12989 47107 13047 47113
rect 12989 47104 13001 47107
rect 12483 47076 13001 47104
rect 12483 47073 12495 47076
rect 12437 47067 12495 47073
rect 12989 47073 13001 47076
rect 13035 47073 13047 47107
rect 12989 47067 13047 47073
rect 13173 47107 13231 47113
rect 13173 47073 13185 47107
rect 13219 47104 13231 47107
rect 13219 47076 13860 47104
rect 13219 47073 13231 47076
rect 13173 47067 13231 47073
rect 5629 47039 5687 47045
rect 5629 47036 5641 47039
rect 4356 47008 5641 47036
rect 4249 46999 4307 47005
rect 5629 47005 5641 47008
rect 5675 47005 5687 47039
rect 5629 46999 5687 47005
rect 12253 47039 12311 47045
rect 12253 47005 12265 47039
rect 12299 47005 12311 47039
rect 12253 46999 12311 47005
rect 4264 46900 4292 46999
rect 6089 46971 6147 46977
rect 6089 46937 6101 46971
rect 6135 46968 6147 46971
rect 12066 46968 12072 46980
rect 6135 46940 6868 46968
rect 12027 46940 12072 46968
rect 6135 46937 6147 46940
rect 6089 46931 6147 46937
rect 4706 46900 4712 46912
rect 4264 46872 4712 46900
rect 4706 46860 4712 46872
rect 4764 46860 4770 46912
rect 6840 46900 6868 46940
rect 12066 46928 12072 46940
rect 12124 46968 12130 46980
rect 12268 46968 12296 46999
rect 13354 46968 13360 46980
rect 12124 46940 12296 46968
rect 13315 46940 13360 46968
rect 12124 46928 12130 46940
rect 13354 46928 13360 46940
rect 13412 46928 13418 46980
rect 13832 46977 13860 47076
rect 13924 47045 13952 47144
rect 22480 47104 22508 47200
rect 23290 47132 23296 47184
rect 23348 47172 23354 47184
rect 23348 47144 23612 47172
rect 23348 47132 23354 47144
rect 22649 47107 22707 47113
rect 22649 47104 22661 47107
rect 22480 47076 22661 47104
rect 22649 47073 22661 47076
rect 22695 47073 22707 47107
rect 22649 47067 22707 47073
rect 22833 47107 22891 47113
rect 22833 47073 22845 47107
rect 22879 47104 22891 47107
rect 23382 47104 23388 47116
rect 22879 47076 23388 47104
rect 22879 47073 22891 47076
rect 22833 47067 22891 47073
rect 23382 47064 23388 47076
rect 23440 47064 23446 47116
rect 23584 47113 23612 47144
rect 46676 47144 47164 47172
rect 46676 47116 46704 47144
rect 23569 47107 23627 47113
rect 23569 47073 23581 47107
rect 23615 47104 23627 47107
rect 25406 47104 25412 47116
rect 23615 47076 24256 47104
rect 25367 47076 25412 47104
rect 23615 47073 23627 47076
rect 23569 47067 23627 47073
rect 13909 47039 13967 47045
rect 13909 47005 13921 47039
rect 13955 47036 13967 47039
rect 17129 47039 17187 47045
rect 17129 47036 17141 47039
rect 13955 47008 14228 47036
rect 13955 47005 13967 47008
rect 13909 46999 13967 47005
rect 14200 46980 14228 47008
rect 16960 47008 17141 47036
rect 13817 46971 13875 46977
rect 13817 46937 13829 46971
rect 13863 46968 13875 46971
rect 13998 46968 14004 46980
rect 13863 46940 14004 46968
rect 13863 46937 13875 46940
rect 13817 46931 13875 46937
rect 13998 46928 14004 46940
rect 14056 46928 14062 46980
rect 14182 46968 14188 46980
rect 14143 46940 14188 46968
rect 14182 46928 14188 46940
rect 14240 46928 14246 46980
rect 7190 46900 7196 46912
rect 6840 46872 7196 46900
rect 7190 46860 7196 46872
rect 7248 46860 7254 46912
rect 15470 46860 15476 46912
rect 15528 46900 15534 46912
rect 16960 46909 16988 47008
rect 17129 47005 17141 47008
rect 17175 47005 17187 47039
rect 17129 46999 17187 47005
rect 17405 47039 17463 47045
rect 17405 47005 17417 47039
rect 17451 47036 17463 47039
rect 18046 47036 18052 47048
rect 17451 47008 18052 47036
rect 17451 47005 17463 47008
rect 17405 46999 17463 47005
rect 18046 46996 18052 47008
rect 18104 46996 18110 47048
rect 23382 46928 23388 46980
rect 23440 46968 23446 46980
rect 23934 46968 23940 46980
rect 23440 46940 23940 46968
rect 23440 46928 23446 46940
rect 23934 46928 23940 46940
rect 23992 46928 23998 46980
rect 24228 46977 24256 47076
rect 25406 47064 25412 47076
rect 25464 47064 25470 47116
rect 34333 47107 34391 47113
rect 34333 47104 34345 47107
rect 32600 47076 34345 47104
rect 32600 47048 32628 47076
rect 34333 47073 34345 47076
rect 34379 47073 34391 47107
rect 34333 47067 34391 47073
rect 43349 47107 43407 47113
rect 43349 47073 43361 47107
rect 43395 47104 43407 47107
rect 44358 47104 44364 47116
rect 43395 47076 44364 47104
rect 43395 47073 43407 47076
rect 43349 47067 43407 47073
rect 44358 47064 44364 47076
rect 44416 47064 44422 47116
rect 45557 47107 45615 47113
rect 45557 47073 45569 47107
rect 45603 47073 45615 47107
rect 45557 47067 45615 47073
rect 45925 47107 45983 47113
rect 45925 47073 45937 47107
rect 45971 47104 45983 47107
rect 46658 47104 46664 47116
rect 45971 47076 46664 47104
rect 45971 47073 45983 47076
rect 45925 47067 45983 47073
rect 32582 47036 32588 47048
rect 32543 47008 32588 47036
rect 32582 46996 32588 47008
rect 32640 46996 32646 47048
rect 32858 47036 32864 47048
rect 32819 47008 32864 47036
rect 32858 46996 32864 47008
rect 32916 46996 32922 47048
rect 38933 47039 38991 47045
rect 38933 47005 38945 47039
rect 38979 47005 38991 47039
rect 38933 46999 38991 47005
rect 39209 47039 39267 47045
rect 39209 47005 39221 47039
rect 39255 47036 39267 47039
rect 40586 47036 40592 47048
rect 39255 47008 40592 47036
rect 39255 47005 39267 47008
rect 39209 46999 39267 47005
rect 24213 46971 24271 46977
rect 24213 46937 24225 46971
rect 24259 46968 24271 46971
rect 25501 46971 25559 46977
rect 25501 46968 25513 46971
rect 24259 46940 25513 46968
rect 24259 46937 24271 46940
rect 24213 46931 24271 46937
rect 25501 46937 25513 46940
rect 25547 46937 25559 46971
rect 38746 46968 38752 46980
rect 38707 46940 38752 46968
rect 25501 46931 25559 46937
rect 16945 46903 17003 46909
rect 16945 46900 16957 46903
rect 15528 46872 16957 46900
rect 15528 46860 15534 46872
rect 16945 46869 16957 46872
rect 16991 46869 17003 46903
rect 16945 46863 17003 46869
rect 18693 46903 18751 46909
rect 18693 46869 18705 46903
rect 18739 46900 18751 46903
rect 19058 46900 19064 46912
rect 18739 46872 19064 46900
rect 18739 46869 18751 46872
rect 18693 46863 18751 46869
rect 19058 46860 19064 46872
rect 19116 46860 19122 46912
rect 23845 46903 23903 46909
rect 23845 46869 23857 46903
rect 23891 46900 23903 46903
rect 24026 46900 24032 46912
rect 23891 46872 24032 46900
rect 23891 46869 23903 46872
rect 23845 46863 23903 46869
rect 24026 46860 24032 46872
rect 24084 46860 24090 46912
rect 25516 46900 25544 46931
rect 38746 46928 38752 46940
rect 38804 46968 38810 46980
rect 38948 46968 38976 46999
rect 40586 46996 40592 47008
rect 40644 46996 40650 47048
rect 40678 46996 40684 47048
rect 40736 47036 40742 47048
rect 44913 47039 44971 47045
rect 44913 47036 44925 47039
rect 40736 47008 44925 47036
rect 40736 46996 40742 47008
rect 44913 47005 44925 47008
rect 44959 47005 44971 47039
rect 44913 46999 44971 47005
rect 45465 47039 45523 47045
rect 45465 47005 45477 47039
rect 45511 47005 45523 47039
rect 45465 46999 45523 47005
rect 38804 46940 38976 46968
rect 38804 46928 38810 46940
rect 31018 46900 31024 46912
rect 25516 46872 31024 46900
rect 31018 46860 31024 46872
rect 31076 46860 31082 46912
rect 33778 46860 33784 46912
rect 33836 46900 33842 46912
rect 33965 46903 34023 46909
rect 33965 46900 33977 46903
rect 33836 46872 33977 46900
rect 33836 46860 33842 46872
rect 33965 46869 33977 46872
rect 34011 46869 34023 46903
rect 33965 46863 34023 46869
rect 40034 46860 40040 46912
rect 40092 46900 40098 46912
rect 40313 46903 40371 46909
rect 40313 46900 40325 46903
rect 40092 46872 40325 46900
rect 40092 46860 40098 46872
rect 40313 46869 40325 46872
rect 40359 46869 40371 46903
rect 43438 46900 43444 46912
rect 43399 46872 43444 46900
rect 40313 46863 40371 46869
rect 43438 46860 43444 46872
rect 43496 46860 43502 46912
rect 45480 46900 45508 46999
rect 45572 46968 45600 47067
rect 46658 47064 46664 47076
rect 46716 47064 46722 47116
rect 47136 47113 47164 47144
rect 46937 47107 46995 47113
rect 46937 47073 46949 47107
rect 46983 47073 46995 47107
rect 46937 47067 46995 47073
rect 47121 47107 47179 47113
rect 47121 47073 47133 47107
rect 47167 47073 47179 47107
rect 47121 47067 47179 47073
rect 49421 47107 49479 47113
rect 49421 47073 49433 47107
rect 49467 47104 49479 47107
rect 50154 47104 50160 47116
rect 49467 47076 50160 47104
rect 49467 47073 49479 47076
rect 49421 47067 49479 47073
rect 46017 47039 46075 47045
rect 46017 47005 46029 47039
rect 46063 47036 46075 47039
rect 46293 47039 46351 47045
rect 46293 47036 46305 47039
rect 46063 47008 46305 47036
rect 46063 47005 46075 47008
rect 46017 46999 46075 47005
rect 46293 47005 46305 47008
rect 46339 47036 46351 47039
rect 46952 47036 46980 47067
rect 50154 47064 50160 47076
rect 50212 47064 50218 47116
rect 50522 47064 50528 47116
rect 50580 47104 50586 47116
rect 50801 47107 50859 47113
rect 50801 47104 50813 47107
rect 50580 47076 50813 47104
rect 50580 47064 50586 47076
rect 50801 47073 50813 47076
rect 50847 47073 50859 47107
rect 50801 47067 50859 47073
rect 50890 47064 50896 47116
rect 50948 47104 50954 47116
rect 50948 47076 50993 47104
rect 50948 47064 50954 47076
rect 51902 47064 51908 47116
rect 51960 47104 51966 47116
rect 52181 47107 52239 47113
rect 52181 47104 52193 47107
rect 51960 47076 52193 47104
rect 51960 47064 51966 47076
rect 52181 47073 52193 47076
rect 52227 47073 52239 47107
rect 56686 47104 56692 47116
rect 56647 47076 56692 47104
rect 52181 47067 52239 47073
rect 56686 47064 56692 47076
rect 56744 47064 56750 47116
rect 56778 47064 56784 47116
rect 56836 47104 56842 47116
rect 61197 47107 61255 47113
rect 56836 47076 56881 47104
rect 56836 47064 56842 47076
rect 61197 47073 61209 47107
rect 61243 47104 61255 47107
rect 62942 47104 62948 47116
rect 61243 47076 62948 47104
rect 61243 47073 61255 47076
rect 61197 47067 61255 47073
rect 62942 47064 62948 47076
rect 63000 47064 63006 47116
rect 47302 47036 47308 47048
rect 46339 47008 47308 47036
rect 46339 47005 46351 47008
rect 46293 46999 46351 47005
rect 47302 46996 47308 47008
rect 47360 46996 47366 47048
rect 47486 47036 47492 47048
rect 47447 47008 47492 47036
rect 47486 46996 47492 47008
rect 47544 46996 47550 47048
rect 51350 47036 51356 47048
rect 51311 47008 51356 47036
rect 51350 46996 51356 47008
rect 51408 46996 51414 47048
rect 57238 47036 57244 47048
rect 57199 47008 57244 47036
rect 57238 46996 57244 47008
rect 57296 46996 57302 47048
rect 61470 47036 61476 47048
rect 61431 47008 61476 47036
rect 61470 46996 61476 47008
rect 61528 46996 61534 47048
rect 47394 46968 47400 46980
rect 45572 46940 47400 46968
rect 47394 46928 47400 46940
rect 47452 46928 47458 46980
rect 50617 46971 50675 46977
rect 50617 46937 50629 46971
rect 50663 46968 50675 46971
rect 51445 46971 51503 46977
rect 51445 46968 51457 46971
rect 50663 46940 51457 46968
rect 50663 46937 50675 46940
rect 50617 46931 50675 46937
rect 51445 46937 51457 46940
rect 51491 46968 51503 46971
rect 56505 46971 56563 46977
rect 56505 46968 56517 46971
rect 51491 46940 56517 46968
rect 51491 46937 51503 46940
rect 51445 46931 51503 46937
rect 56505 46937 56517 46940
rect 56551 46968 56563 46971
rect 57333 46971 57391 46977
rect 57333 46968 57345 46971
rect 56551 46940 57345 46968
rect 56551 46937 56563 46940
rect 56505 46931 56563 46937
rect 57333 46937 57345 46940
rect 57379 46968 57391 46971
rect 59538 46968 59544 46980
rect 57379 46940 59544 46968
rect 57379 46937 57391 46940
rect 57333 46931 57391 46937
rect 59538 46928 59544 46940
rect 59596 46928 59602 46980
rect 46474 46900 46480 46912
rect 45480 46872 46480 46900
rect 46474 46860 46480 46872
rect 46532 46860 46538 46912
rect 47302 46860 47308 46912
rect 47360 46900 47366 46912
rect 47581 46903 47639 46909
rect 47581 46900 47593 46903
rect 47360 46872 47593 46900
rect 47360 46860 47366 46872
rect 47581 46869 47593 46872
rect 47627 46869 47639 46903
rect 47581 46863 47639 46869
rect 48682 46860 48688 46912
rect 48740 46900 48746 46912
rect 49513 46903 49571 46909
rect 49513 46900 49525 46903
rect 48740 46872 49525 46900
rect 48740 46860 48746 46872
rect 49513 46869 49525 46872
rect 49559 46869 49571 46903
rect 49513 46863 49571 46869
rect 51718 46860 51724 46912
rect 51776 46900 51782 46912
rect 52362 46900 52368 46912
rect 51776 46872 52368 46900
rect 51776 46860 51782 46872
rect 52362 46860 52368 46872
rect 52420 46860 52426 46912
rect 62114 46860 62120 46912
rect 62172 46900 62178 46912
rect 62577 46903 62635 46909
rect 62577 46900 62589 46903
rect 62172 46872 62589 46900
rect 62172 46860 62178 46872
rect 62577 46869 62589 46872
rect 62623 46869 62635 46903
rect 62942 46900 62948 46912
rect 62903 46872 62948 46900
rect 62577 46863 62635 46869
rect 62942 46860 62948 46872
rect 63000 46860 63006 46912
rect 1104 46810 108008 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 65686 46810
rect 65738 46758 65750 46810
rect 65802 46758 65814 46810
rect 65866 46758 65878 46810
rect 65930 46758 96406 46810
rect 96458 46758 96470 46810
rect 96522 46758 96534 46810
rect 96586 46758 96598 46810
rect 96650 46758 108008 46810
rect 1104 46736 108008 46758
rect 2501 46699 2559 46705
rect 2501 46665 2513 46699
rect 2547 46696 2559 46699
rect 2774 46696 2780 46708
rect 2547 46668 2780 46696
rect 2547 46665 2559 46668
rect 2501 46659 2559 46665
rect 2774 46656 2780 46668
rect 2832 46656 2838 46708
rect 22278 46656 22284 46708
rect 22336 46696 22342 46708
rect 24946 46696 24952 46708
rect 22336 46668 24952 46696
rect 22336 46656 22342 46668
rect 24946 46656 24952 46668
rect 25004 46656 25010 46708
rect 25317 46699 25375 46705
rect 25317 46665 25329 46699
rect 25363 46696 25375 46699
rect 25406 46696 25412 46708
rect 25363 46668 25412 46696
rect 25363 46665 25375 46668
rect 25317 46659 25375 46665
rect 25406 46656 25412 46668
rect 25464 46656 25470 46708
rect 37277 46699 37335 46705
rect 37277 46696 37289 46699
rect 26436 46668 37289 46696
rect 13998 46588 14004 46640
rect 14056 46628 14062 46640
rect 19981 46631 20039 46637
rect 19981 46628 19993 46631
rect 14056 46600 19993 46628
rect 14056 46588 14062 46600
rect 19981 46597 19993 46600
rect 20027 46628 20039 46631
rect 20027 46600 20852 46628
rect 20027 46597 20039 46600
rect 19981 46591 20039 46597
rect 2774 46520 2780 46572
rect 2832 46560 2838 46572
rect 2869 46563 2927 46569
rect 2869 46560 2881 46563
rect 2832 46532 2881 46560
rect 2832 46520 2838 46532
rect 2869 46529 2881 46532
rect 2915 46529 2927 46563
rect 2869 46523 2927 46529
rect 7561 46563 7619 46569
rect 7561 46529 7573 46563
rect 7607 46560 7619 46563
rect 8386 46560 8392 46572
rect 7607 46532 8392 46560
rect 7607 46529 7619 46532
rect 7561 46523 7619 46529
rect 8386 46520 8392 46532
rect 8444 46520 8450 46572
rect 9125 46563 9183 46569
rect 9125 46529 9137 46563
rect 9171 46560 9183 46563
rect 12437 46563 12495 46569
rect 12437 46560 12449 46563
rect 9171 46532 12449 46560
rect 9171 46529 9183 46532
rect 9125 46523 9183 46529
rect 12437 46529 12449 46532
rect 12483 46529 12495 46563
rect 12437 46523 12495 46529
rect 12713 46563 12771 46569
rect 12713 46529 12725 46563
rect 12759 46560 12771 46563
rect 13354 46560 13360 46572
rect 12759 46532 13360 46560
rect 12759 46529 12771 46532
rect 12713 46523 12771 46529
rect 2590 46492 2596 46504
rect 2551 46464 2596 46492
rect 2590 46452 2596 46464
rect 2648 46452 2654 46504
rect 7190 46452 7196 46504
rect 7248 46492 7254 46504
rect 7285 46495 7343 46501
rect 7285 46492 7297 46495
rect 7248 46464 7297 46492
rect 7248 46452 7254 46464
rect 7285 46461 7297 46464
rect 7331 46492 7343 46495
rect 9140 46492 9168 46523
rect 7331 46464 9168 46492
rect 12452 46492 12480 46523
rect 13354 46520 13360 46532
rect 13412 46520 13418 46572
rect 13722 46520 13728 46572
rect 13780 46560 13786 46572
rect 20824 46569 20852 46600
rect 20073 46563 20131 46569
rect 20073 46560 20085 46563
rect 13780 46532 20085 46560
rect 13780 46520 13786 46532
rect 20073 46529 20085 46532
rect 20119 46529 20131 46563
rect 20073 46523 20131 46529
rect 20809 46563 20867 46569
rect 20809 46529 20821 46563
rect 20855 46560 20867 46563
rect 26436 46560 26464 46668
rect 37277 46665 37289 46668
rect 37323 46696 37335 46699
rect 37461 46699 37519 46705
rect 37461 46696 37473 46699
rect 37323 46668 37473 46696
rect 37323 46665 37335 46668
rect 37277 46659 37335 46665
rect 37461 46665 37473 46668
rect 37507 46696 37519 46699
rect 40586 46696 40592 46708
rect 37507 46668 37688 46696
rect 40547 46668 40592 46696
rect 37507 46665 37519 46668
rect 37461 46659 37519 46665
rect 20855 46532 26464 46560
rect 20855 46529 20867 46532
rect 20809 46523 20867 46529
rect 30834 46520 30840 46572
rect 30892 46560 30898 46572
rect 37660 46569 37688 46668
rect 40586 46656 40592 46668
rect 40644 46656 40650 46708
rect 47394 46656 47400 46708
rect 47452 46696 47458 46708
rect 47581 46699 47639 46705
rect 47581 46696 47593 46699
rect 47452 46668 47593 46696
rect 47452 46656 47458 46668
rect 47581 46665 47593 46668
rect 47627 46665 47639 46699
rect 47581 46659 47639 46665
rect 48777 46699 48835 46705
rect 48777 46665 48789 46699
rect 48823 46696 48835 46699
rect 50890 46696 50896 46708
rect 48823 46668 50896 46696
rect 48823 46665 48835 46668
rect 48777 46659 48835 46665
rect 50890 46656 50896 46668
rect 50948 46656 50954 46708
rect 54941 46699 54999 46705
rect 54941 46696 54953 46699
rect 51736 46668 54953 46696
rect 45002 46588 45008 46640
rect 45060 46628 45066 46640
rect 51736 46628 51764 46668
rect 54941 46665 54953 46668
rect 54987 46665 54999 46699
rect 62114 46696 62120 46708
rect 62075 46668 62120 46696
rect 54941 46659 54999 46665
rect 45060 46600 51764 46628
rect 45060 46588 45066 46600
rect 31113 46563 31171 46569
rect 31113 46560 31125 46563
rect 30892 46532 31125 46560
rect 30892 46520 30898 46532
rect 31113 46529 31125 46532
rect 31159 46529 31171 46563
rect 31113 46523 31171 46529
rect 37645 46563 37703 46569
rect 37645 46529 37657 46563
rect 37691 46560 37703 46563
rect 42521 46563 42579 46569
rect 37691 46532 37964 46560
rect 37691 46529 37703 46532
rect 37645 46523 37703 46529
rect 13446 46492 13452 46504
rect 12452 46464 13452 46492
rect 7331 46461 7343 46464
rect 7285 46455 7343 46461
rect 13446 46452 13452 46464
rect 13504 46492 13510 46504
rect 14185 46495 14243 46501
rect 14185 46492 14197 46495
rect 13504 46464 14197 46492
rect 13504 46452 13510 46464
rect 14185 46461 14197 46464
rect 14231 46461 14243 46495
rect 14185 46455 14243 46461
rect 18049 46495 18107 46501
rect 18049 46461 18061 46495
rect 18095 46492 18107 46495
rect 18138 46492 18144 46504
rect 18095 46464 18144 46492
rect 18095 46461 18107 46464
rect 18049 46455 18107 46461
rect 18138 46452 18144 46464
rect 18196 46452 18202 46504
rect 19058 46492 19064 46504
rect 19019 46464 19064 46492
rect 19058 46452 19064 46464
rect 19116 46452 19122 46504
rect 20714 46492 20720 46504
rect 20675 46464 20720 46492
rect 20714 46452 20720 46464
rect 20772 46452 20778 46504
rect 21085 46495 21143 46501
rect 21085 46461 21097 46495
rect 21131 46461 21143 46495
rect 21085 46455 21143 46461
rect 21269 46495 21327 46501
rect 21269 46461 21281 46495
rect 21315 46492 21327 46495
rect 21453 46495 21511 46501
rect 21453 46492 21465 46495
rect 21315 46464 21465 46492
rect 21315 46461 21327 46464
rect 21269 46455 21327 46461
rect 21453 46461 21465 46464
rect 21499 46492 21511 46495
rect 23290 46492 23296 46504
rect 21499 46464 23296 46492
rect 21499 46461 21511 46464
rect 21453 46455 21511 46461
rect 21100 46424 21128 46455
rect 23290 46452 23296 46464
rect 23348 46452 23354 46504
rect 23937 46495 23995 46501
rect 23937 46492 23949 46495
rect 23768 46464 23949 46492
rect 21910 46424 21916 46436
rect 21100 46396 21916 46424
rect 21910 46384 21916 46396
rect 21968 46384 21974 46436
rect 4154 46356 4160 46368
rect 4115 46328 4160 46356
rect 4154 46316 4160 46328
rect 4212 46316 4218 46368
rect 4433 46359 4491 46365
rect 4433 46325 4445 46359
rect 4479 46356 4491 46359
rect 4706 46356 4712 46368
rect 4479 46328 4712 46356
rect 4479 46325 4491 46328
rect 4433 46319 4491 46325
rect 4706 46316 4712 46328
rect 4764 46316 4770 46368
rect 7926 46316 7932 46368
rect 7984 46356 7990 46368
rect 8665 46359 8723 46365
rect 8665 46356 8677 46359
rect 7984 46328 8677 46356
rect 7984 46316 7990 46328
rect 8665 46325 8677 46328
rect 8711 46325 8723 46359
rect 8665 46319 8723 46325
rect 13906 46316 13912 46368
rect 13964 46356 13970 46368
rect 14001 46359 14059 46365
rect 14001 46356 14013 46359
rect 13964 46328 14013 46356
rect 13964 46316 13970 46328
rect 14001 46325 14013 46328
rect 14047 46325 14059 46359
rect 18138 46356 18144 46368
rect 18099 46328 18144 46356
rect 14001 46319 14059 46325
rect 18138 46316 18144 46328
rect 18196 46316 18202 46368
rect 19150 46356 19156 46368
rect 19111 46328 19156 46356
rect 19150 46316 19156 46328
rect 19208 46316 19214 46368
rect 21818 46316 21824 46368
rect 21876 46356 21882 46368
rect 23768 46365 23796 46464
rect 23937 46461 23949 46464
rect 23983 46461 23995 46495
rect 23937 46455 23995 46461
rect 24026 46452 24032 46504
rect 24084 46492 24090 46504
rect 24213 46495 24271 46501
rect 24213 46492 24225 46495
rect 24084 46464 24225 46492
rect 24084 46452 24090 46464
rect 24213 46461 24225 46464
rect 24259 46461 24271 46495
rect 26421 46495 26479 46501
rect 26421 46492 26433 46495
rect 24213 46455 24271 46461
rect 26252 46464 26433 46492
rect 26252 46365 26280 46464
rect 26421 46461 26433 46464
rect 26467 46461 26479 46495
rect 26694 46492 26700 46504
rect 26655 46464 26700 46492
rect 26421 46455 26479 46461
rect 26694 46452 26700 46464
rect 26752 46452 26758 46504
rect 29178 46452 29184 46504
rect 29236 46492 29242 46504
rect 31297 46495 31355 46501
rect 31297 46492 31309 46495
rect 29236 46464 31309 46492
rect 29236 46452 29242 46464
rect 31297 46461 31309 46464
rect 31343 46461 31355 46495
rect 31297 46455 31355 46461
rect 31849 46495 31907 46501
rect 31849 46461 31861 46495
rect 31895 46492 31907 46495
rect 31938 46492 31944 46504
rect 31895 46464 31944 46492
rect 31895 46461 31907 46464
rect 31849 46455 31907 46461
rect 31938 46452 31944 46464
rect 31996 46452 32002 46504
rect 32030 46452 32036 46504
rect 32088 46492 32094 46504
rect 33778 46492 33784 46504
rect 32088 46464 32720 46492
rect 33739 46464 33784 46492
rect 32088 46452 32094 46464
rect 32692 46433 32720 46464
rect 33778 46452 33784 46464
rect 33836 46452 33842 46504
rect 34422 46452 34428 46504
rect 34480 46492 34486 46504
rect 34885 46495 34943 46501
rect 34885 46492 34897 46495
rect 34480 46464 34897 46492
rect 34480 46452 34486 46464
rect 34885 46461 34897 46464
rect 34931 46461 34943 46495
rect 34885 46455 34943 46461
rect 37829 46495 37887 46501
rect 37829 46461 37841 46495
rect 37875 46461 37887 46495
rect 37936 46492 37964 46532
rect 42521 46529 42533 46563
rect 42567 46560 42579 46563
rect 43438 46560 43444 46572
rect 42567 46532 43444 46560
rect 42567 46529 42579 46532
rect 42521 46523 42579 46529
rect 43438 46520 43444 46532
rect 43496 46520 43502 46572
rect 45370 46520 45376 46572
rect 45428 46560 45434 46572
rect 46661 46563 46719 46569
rect 45428 46532 46336 46560
rect 45428 46520 45434 46532
rect 38289 46495 38347 46501
rect 38289 46492 38301 46495
rect 37936 46464 38301 46492
rect 37829 46455 37887 46461
rect 38289 46461 38301 46464
rect 38335 46461 38347 46495
rect 38289 46455 38347 46461
rect 38381 46495 38439 46501
rect 38381 46461 38393 46495
rect 38427 46461 38439 46495
rect 38381 46455 38439 46461
rect 32677 46427 32735 46433
rect 32677 46393 32689 46427
rect 32723 46424 32735 46427
rect 37844 46424 37872 46455
rect 38396 46424 38424 46455
rect 38746 46452 38752 46504
rect 38804 46492 38810 46504
rect 40497 46495 40555 46501
rect 38804 46464 39068 46492
rect 38804 46452 38810 46464
rect 38930 46424 38936 46436
rect 32723 46396 35020 46424
rect 37844 46396 38424 46424
rect 38891 46396 38936 46424
rect 32723 46393 32735 46396
rect 32677 46387 32735 46393
rect 34992 46368 35020 46396
rect 23753 46359 23811 46365
rect 23753 46356 23765 46359
rect 21876 46328 23765 46356
rect 21876 46316 21882 46328
rect 23753 46325 23765 46328
rect 23799 46356 23811 46359
rect 26237 46359 26295 46365
rect 26237 46356 26249 46359
rect 23799 46328 26249 46356
rect 23799 46325 23811 46328
rect 23753 46319 23811 46325
rect 26237 46325 26249 46328
rect 26283 46325 26295 46359
rect 26237 46319 26295 46325
rect 27062 46316 27068 46368
rect 27120 46356 27126 46368
rect 27801 46359 27859 46365
rect 27801 46356 27813 46359
rect 27120 46328 27813 46356
rect 27120 46316 27126 46328
rect 27801 46325 27813 46328
rect 27847 46325 27859 46359
rect 27801 46319 27859 46325
rect 30834 46316 30840 46368
rect 30892 46356 30898 46368
rect 30929 46359 30987 46365
rect 30929 46356 30941 46359
rect 30892 46328 30941 46356
rect 30892 46316 30898 46328
rect 30929 46325 30941 46328
rect 30975 46325 30987 46359
rect 30929 46319 30987 46325
rect 31018 46316 31024 46368
rect 31076 46356 31082 46368
rect 32122 46356 32128 46368
rect 31076 46328 32128 46356
rect 31076 46316 31082 46328
rect 32122 46316 32128 46328
rect 32180 46316 32186 46368
rect 32306 46356 32312 46368
rect 32267 46328 32312 46356
rect 32306 46316 32312 46328
rect 32364 46316 32370 46368
rect 33870 46356 33876 46368
rect 33831 46328 33876 46356
rect 33870 46316 33876 46328
rect 33928 46316 33934 46368
rect 34974 46356 34980 46368
rect 34935 46328 34980 46356
rect 34974 46316 34980 46328
rect 35032 46316 35038 46368
rect 38396 46356 38424 46396
rect 38930 46384 38936 46396
rect 38988 46384 38994 46436
rect 39040 46424 39068 46464
rect 40497 46461 40509 46495
rect 40543 46492 40555 46495
rect 40678 46492 40684 46504
rect 40543 46464 40684 46492
rect 40543 46461 40555 46464
rect 40497 46455 40555 46461
rect 40678 46452 40684 46464
rect 40736 46452 40742 46504
rect 46308 46501 46336 46532
rect 46661 46529 46673 46563
rect 46707 46560 46719 46563
rect 50522 46560 50528 46572
rect 46707 46532 50108 46560
rect 50483 46532 50528 46560
rect 46707 46529 46719 46532
rect 46661 46523 46719 46529
rect 42245 46495 42303 46501
rect 42245 46461 42257 46495
rect 42291 46461 42303 46495
rect 46293 46495 46351 46501
rect 42245 46455 42303 46461
rect 43548 46464 46244 46492
rect 42061 46427 42119 46433
rect 42061 46424 42073 46427
rect 39040 46396 42073 46424
rect 42061 46393 42073 46396
rect 42107 46424 42119 46427
rect 42260 46424 42288 46455
rect 42107 46396 42288 46424
rect 42107 46393 42119 46396
rect 42061 46387 42119 46393
rect 38470 46356 38476 46368
rect 38383 46328 38476 46356
rect 38470 46316 38476 46328
rect 38528 46356 38534 46368
rect 39206 46356 39212 46368
rect 38528 46328 39212 46356
rect 38528 46316 38534 46328
rect 39206 46316 39212 46328
rect 39264 46356 39270 46368
rect 39393 46359 39451 46365
rect 39393 46356 39405 46359
rect 39264 46328 39405 46356
rect 39264 46316 39270 46328
rect 39393 46325 39405 46328
rect 39439 46356 39451 46359
rect 43548 46356 43576 46464
rect 43901 46427 43959 46433
rect 43901 46393 43913 46427
rect 43947 46424 43959 46427
rect 44450 46424 44456 46436
rect 43947 46396 44456 46424
rect 43947 46393 43959 46396
rect 43901 46387 43959 46393
rect 44450 46384 44456 46396
rect 44508 46384 44514 46436
rect 46106 46424 46112 46436
rect 46067 46396 46112 46424
rect 46106 46384 46112 46396
rect 46164 46384 46170 46436
rect 46216 46424 46244 46464
rect 46293 46461 46305 46495
rect 46339 46492 46351 46495
rect 46753 46495 46811 46501
rect 46753 46492 46765 46495
rect 46339 46464 46765 46492
rect 46339 46461 46351 46464
rect 46293 46455 46351 46461
rect 46753 46461 46765 46464
rect 46799 46461 46811 46495
rect 47486 46492 47492 46504
rect 47447 46464 47492 46492
rect 46753 46455 46811 46461
rect 47486 46452 47492 46464
rect 47544 46492 47550 46504
rect 48501 46495 48559 46501
rect 48501 46492 48513 46495
rect 47544 46464 48513 46492
rect 47544 46452 47550 46464
rect 48501 46461 48513 46464
rect 48547 46461 48559 46495
rect 48682 46492 48688 46504
rect 48643 46464 48688 46492
rect 48501 46455 48559 46461
rect 48682 46452 48688 46464
rect 48740 46452 48746 46504
rect 46934 46424 46940 46436
rect 46216 46396 46940 46424
rect 46934 46384 46940 46396
rect 46992 46384 46998 46436
rect 47394 46384 47400 46436
rect 47452 46424 47458 46436
rect 49973 46427 50031 46433
rect 49973 46424 49985 46427
rect 47452 46396 49985 46424
rect 47452 46384 47458 46396
rect 49973 46393 49985 46396
rect 50019 46393 50031 46427
rect 50080 46424 50108 46532
rect 50522 46520 50528 46532
rect 50580 46520 50586 46572
rect 51350 46520 51356 46572
rect 51408 46560 51414 46572
rect 51997 46563 52055 46569
rect 51997 46560 52009 46563
rect 51408 46532 52009 46560
rect 51408 46520 51414 46532
rect 51997 46529 52009 46532
rect 52043 46529 52055 46563
rect 51997 46523 52055 46529
rect 50154 46452 50160 46504
rect 50212 46492 50218 46504
rect 51166 46492 51172 46504
rect 50212 46464 51172 46492
rect 50212 46452 50218 46464
rect 51166 46452 51172 46464
rect 51224 46452 51230 46504
rect 51442 46452 51448 46504
rect 51500 46492 51506 46504
rect 51721 46495 51779 46501
rect 51721 46492 51733 46495
rect 51500 46464 51733 46492
rect 51500 46452 51506 46464
rect 51721 46461 51733 46464
rect 51767 46461 51779 46495
rect 54846 46492 54852 46504
rect 51721 46455 51779 46461
rect 51828 46464 54852 46492
rect 51828 46424 51856 46464
rect 54846 46452 54852 46464
rect 54904 46452 54910 46504
rect 54956 46492 54984 46659
rect 62114 46656 62120 46668
rect 62172 46656 62178 46708
rect 56413 46563 56471 46569
rect 56413 46529 56425 46563
rect 56459 46560 56471 46563
rect 56686 46560 56692 46572
rect 56459 46532 56692 46560
rect 56459 46529 56471 46532
rect 56413 46523 56471 46529
rect 56686 46520 56692 46532
rect 56744 46520 56750 46572
rect 57238 46520 57244 46572
rect 57296 46560 57302 46572
rect 57609 46563 57667 46569
rect 57609 46560 57621 46563
rect 57296 46532 57621 46560
rect 57296 46520 57302 46532
rect 57609 46529 57621 46532
rect 57655 46529 57667 46563
rect 57609 46523 57667 46529
rect 55861 46495 55919 46501
rect 55861 46492 55873 46495
rect 54956 46464 55873 46492
rect 55861 46461 55873 46464
rect 55907 46461 55919 46495
rect 55861 46455 55919 46461
rect 56045 46495 56103 46501
rect 56045 46461 56057 46495
rect 56091 46492 56103 46495
rect 57330 46492 57336 46504
rect 56091 46464 56640 46492
rect 57291 46464 57336 46492
rect 56091 46461 56103 46464
rect 56045 46455 56103 46461
rect 50080 46396 51856 46424
rect 49973 46387 50031 46393
rect 56612 46368 56640 46464
rect 57330 46452 57336 46464
rect 57388 46452 57394 46504
rect 57422 46452 57428 46504
rect 57480 46492 57486 46504
rect 61749 46495 61807 46501
rect 61749 46492 61761 46495
rect 57480 46464 61761 46492
rect 57480 46452 57486 46464
rect 61749 46461 61761 46464
rect 61795 46492 61807 46495
rect 62114 46492 62120 46504
rect 61795 46464 62120 46492
rect 61795 46461 61807 46464
rect 61749 46455 61807 46461
rect 62114 46452 62120 46464
rect 62172 46452 62178 46504
rect 39439 46328 43576 46356
rect 39439 46325 39451 46328
rect 39393 46319 39451 46325
rect 51350 46316 51356 46368
rect 51408 46356 51414 46368
rect 51445 46359 51503 46365
rect 51445 46356 51457 46359
rect 51408 46328 51457 46356
rect 51408 46316 51414 46328
rect 51445 46325 51457 46328
rect 51491 46325 51503 46359
rect 51445 46319 51503 46325
rect 51994 46316 52000 46368
rect 52052 46356 52058 46368
rect 53101 46359 53159 46365
rect 53101 46356 53113 46359
rect 52052 46328 53113 46356
rect 52052 46316 52058 46328
rect 53101 46325 53113 46328
rect 53147 46325 53159 46359
rect 56594 46356 56600 46368
rect 56555 46328 56600 46356
rect 53101 46319 53159 46325
rect 56594 46316 56600 46328
rect 56652 46356 56658 46368
rect 58713 46359 58771 46365
rect 58713 46356 58725 46359
rect 56652 46328 58725 46356
rect 56652 46316 56658 46328
rect 58713 46325 58725 46328
rect 58759 46325 58771 46359
rect 59170 46356 59176 46368
rect 59131 46328 59176 46356
rect 58713 46319 58771 46325
rect 59170 46316 59176 46328
rect 59228 46316 59234 46368
rect 61841 46359 61899 46365
rect 61841 46325 61853 46359
rect 61887 46356 61899 46359
rect 62022 46356 62028 46368
rect 61887 46328 62028 46356
rect 61887 46325 61899 46328
rect 61841 46319 61899 46325
rect 62022 46316 62028 46328
rect 62080 46316 62086 46368
rect 83826 46316 83832 46368
rect 83884 46356 83890 46368
rect 90818 46356 90824 46368
rect 83884 46328 90824 46356
rect 83884 46316 83890 46328
rect 90818 46316 90824 46328
rect 90876 46316 90882 46368
rect 1104 46266 108008 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 50326 46266
rect 50378 46214 50390 46266
rect 50442 46214 50454 46266
rect 50506 46214 50518 46266
rect 50570 46214 81046 46266
rect 81098 46214 81110 46266
rect 81162 46214 81174 46266
rect 81226 46214 81238 46266
rect 81290 46214 108008 46266
rect 1104 46192 108008 46214
rect 4614 46112 4620 46164
rect 4672 46152 4678 46164
rect 8021 46155 8079 46161
rect 8021 46152 8033 46155
rect 4672 46124 8033 46152
rect 4672 46112 4678 46124
rect 8021 46121 8033 46124
rect 8067 46121 8079 46155
rect 13998 46152 14004 46164
rect 13959 46124 14004 46152
rect 8021 46115 8079 46121
rect 13998 46112 14004 46124
rect 14056 46112 14062 46164
rect 18601 46155 18659 46161
rect 18601 46152 18613 46155
rect 17512 46124 18613 46152
rect 7098 45976 7104 46028
rect 7156 46016 7162 46028
rect 8018 46016 8024 46028
rect 7156 45988 8024 46016
rect 7156 45976 7162 45988
rect 8018 45976 8024 45988
rect 8076 45976 8082 46028
rect 8389 46019 8447 46025
rect 8389 45985 8401 46019
rect 8435 45985 8447 46019
rect 13906 46016 13912 46028
rect 13867 45988 13912 46016
rect 8389 45979 8447 45985
rect 8404 45812 8432 45979
rect 13906 45976 13912 45988
rect 13964 45976 13970 46028
rect 14182 45976 14188 46028
rect 14240 46016 14246 46028
rect 17037 46019 17095 46025
rect 17037 46016 17049 46019
rect 14240 45988 17049 46016
rect 14240 45976 14246 45988
rect 17037 45985 17049 45988
rect 17083 46016 17095 46019
rect 17512 46016 17540 46124
rect 18601 46121 18613 46124
rect 18647 46152 18659 46155
rect 18785 46155 18843 46161
rect 18785 46152 18797 46155
rect 18647 46124 18797 46152
rect 18647 46121 18659 46124
rect 18601 46115 18659 46121
rect 18785 46121 18797 46124
rect 18831 46152 18843 46155
rect 23382 46152 23388 46164
rect 18831 46124 23388 46152
rect 18831 46121 18843 46124
rect 18785 46115 18843 46121
rect 23382 46112 23388 46124
rect 23440 46112 23446 46164
rect 24949 46155 25007 46161
rect 24949 46121 24961 46155
rect 24995 46152 25007 46155
rect 26694 46152 26700 46164
rect 24995 46124 26700 46152
rect 24995 46121 25007 46124
rect 24949 46115 25007 46121
rect 26694 46112 26700 46124
rect 26752 46112 26758 46164
rect 31941 46155 31999 46161
rect 31941 46152 31953 46155
rect 26804 46124 31953 46152
rect 22646 46084 22652 46096
rect 21560 46056 22652 46084
rect 17589 46019 17647 46025
rect 17589 46016 17601 46019
rect 17083 45988 17601 46016
rect 17083 45985 17095 45988
rect 17037 45979 17095 45985
rect 17589 45985 17601 45988
rect 17635 45985 17647 46019
rect 17589 45979 17647 45985
rect 17773 46019 17831 46025
rect 17773 45985 17785 46019
rect 17819 46016 17831 46019
rect 18325 46019 18383 46025
rect 18325 46016 18337 46019
rect 17819 45988 18337 46016
rect 17819 45985 17831 45988
rect 17773 45979 17831 45985
rect 18325 45985 18337 45988
rect 18371 46016 18383 46019
rect 19150 46016 19156 46028
rect 18371 45988 19156 46016
rect 18371 45985 18383 45988
rect 18325 45979 18383 45985
rect 19150 45976 19156 45988
rect 19208 46016 19214 46028
rect 20625 46019 20683 46025
rect 20625 46016 20637 46019
rect 19208 45988 20637 46016
rect 19208 45976 19214 45988
rect 20625 45985 20637 45988
rect 20671 45985 20683 46019
rect 20625 45979 20683 45985
rect 16945 45951 17003 45957
rect 16945 45917 16957 45951
rect 16991 45917 17003 45951
rect 18046 45948 18052 45960
rect 18007 45920 18052 45948
rect 16945 45911 17003 45917
rect 16758 45880 16764 45892
rect 16671 45852 16764 45880
rect 16758 45840 16764 45852
rect 16816 45880 16822 45892
rect 16960 45880 16988 45911
rect 18046 45908 18052 45920
rect 18104 45908 18110 45960
rect 20640 45948 20668 45979
rect 20714 45976 20720 46028
rect 20772 46016 20778 46028
rect 21560 46025 21588 46056
rect 22646 46044 22652 46056
rect 22704 46044 22710 46096
rect 26804 46084 26832 46124
rect 31941 46121 31953 46124
rect 31987 46121 31999 46155
rect 31941 46115 31999 46121
rect 32122 46112 32128 46164
rect 32180 46152 32186 46164
rect 34422 46152 34428 46164
rect 32180 46124 34284 46152
rect 34383 46124 34428 46152
rect 32180 46112 32186 46124
rect 29457 46087 29515 46093
rect 29457 46084 29469 46087
rect 23676 46056 26832 46084
rect 29288 46056 29469 46084
rect 21545 46019 21603 46025
rect 21545 46016 21557 46019
rect 20772 45988 21557 46016
rect 20772 45976 20778 45988
rect 21545 45985 21557 45988
rect 21591 45985 21603 46019
rect 21910 46016 21916 46028
rect 21871 45988 21916 46016
rect 21545 45979 21603 45985
rect 21910 45976 21916 45988
rect 21968 45976 21974 46028
rect 22097 46019 22155 46025
rect 22097 45985 22109 46019
rect 22143 46016 22155 46019
rect 22186 46016 22192 46028
rect 22143 45988 22192 46016
rect 22143 45985 22155 45988
rect 22097 45979 22155 45985
rect 22186 45976 22192 45988
rect 22244 45976 22250 46028
rect 21361 45951 21419 45957
rect 21361 45948 21373 45951
rect 20640 45920 21373 45948
rect 21361 45917 21373 45920
rect 21407 45948 21419 45951
rect 23676 45948 23704 46056
rect 23934 46016 23940 46028
rect 23847 45988 23940 46016
rect 23934 45976 23940 45988
rect 23992 46016 23998 46028
rect 24486 46016 24492 46028
rect 23992 45988 24492 46016
rect 23992 45976 23998 45988
rect 24486 45976 24492 45988
rect 24544 45976 24550 46028
rect 24670 46016 24676 46028
rect 24631 45988 24676 46016
rect 24670 45976 24676 45988
rect 24728 45976 24734 46028
rect 27062 46016 27068 46028
rect 27023 45988 27068 46016
rect 27062 45976 27068 45988
rect 27120 45976 27126 46028
rect 27798 45976 27804 46028
rect 27856 46016 27862 46028
rect 28721 46019 28779 46025
rect 28721 46016 28733 46019
rect 27856 45988 28733 46016
rect 27856 45976 27862 45988
rect 28721 45985 28733 45988
rect 28767 45985 28779 46019
rect 29086 46016 29092 46028
rect 29047 45988 29092 46016
rect 28721 45979 28779 45985
rect 29086 45976 29092 45988
rect 29144 45976 29150 46028
rect 29288 46025 29316 46056
rect 29457 46053 29469 46056
rect 29503 46084 29515 46087
rect 32030 46084 32036 46096
rect 29503 46056 32036 46084
rect 29503 46053 29515 46056
rect 29457 46047 29515 46053
rect 32030 46044 32036 46056
rect 32088 46044 32094 46096
rect 34256 46084 34284 46124
rect 34422 46112 34428 46124
rect 34480 46112 34486 46164
rect 39206 46152 39212 46164
rect 37752 46124 38608 46152
rect 39167 46124 39212 46152
rect 37277 46087 37335 46093
rect 37277 46084 37289 46087
rect 34256 46056 37289 46084
rect 37277 46053 37289 46056
rect 37323 46084 37335 46087
rect 37461 46087 37519 46093
rect 37461 46084 37473 46087
rect 37323 46056 37473 46084
rect 37323 46053 37335 46056
rect 37277 46047 37335 46053
rect 37461 46053 37473 46056
rect 37507 46084 37519 46087
rect 37752 46084 37780 46124
rect 37507 46056 37780 46084
rect 37507 46053 37519 46056
rect 37461 46047 37519 46053
rect 29273 46019 29331 46025
rect 29273 45985 29285 46019
rect 29319 45985 29331 46019
rect 29273 45979 29331 45985
rect 32306 45976 32312 46028
rect 32364 46016 32370 46028
rect 37752 46025 37780 46056
rect 33137 46019 33195 46025
rect 33137 46016 33149 46019
rect 32364 45988 33149 46016
rect 32364 45976 32370 45988
rect 33137 45985 33149 45988
rect 33183 45985 33195 46019
rect 33137 45979 33195 45985
rect 37737 46019 37795 46025
rect 37737 45985 37749 46019
rect 37783 45985 37795 46019
rect 37737 45979 37795 45985
rect 37921 46019 37979 46025
rect 37921 45985 37933 46019
rect 37967 46016 37979 46019
rect 38470 46016 38476 46028
rect 37967 45988 38476 46016
rect 37967 45985 37979 45988
rect 37921 45979 37979 45985
rect 38470 45976 38476 45988
rect 38528 45976 38534 46028
rect 38580 46016 38608 46124
rect 39206 46112 39212 46124
rect 39264 46152 39270 46164
rect 39393 46155 39451 46161
rect 39393 46152 39405 46155
rect 39264 46124 39405 46152
rect 39264 46112 39270 46124
rect 39393 46121 39405 46124
rect 39439 46121 39451 46155
rect 39393 46115 39451 46121
rect 46106 46112 46112 46164
rect 46164 46152 46170 46164
rect 46845 46155 46903 46161
rect 46845 46152 46857 46155
rect 46164 46124 46857 46152
rect 46164 46112 46170 46124
rect 46845 46121 46857 46124
rect 46891 46121 46903 46155
rect 46845 46115 46903 46121
rect 46934 46112 46940 46164
rect 46992 46152 46998 46164
rect 57422 46152 57428 46164
rect 46992 46124 57428 46152
rect 46992 46112 46998 46124
rect 57422 46112 57428 46124
rect 57480 46112 57486 46164
rect 39025 46087 39083 46093
rect 39025 46053 39037 46087
rect 39071 46084 39083 46087
rect 40770 46084 40776 46096
rect 39071 46056 40776 46084
rect 39071 46053 39083 46056
rect 39025 46047 39083 46053
rect 40770 46044 40776 46056
rect 40828 46044 40834 46096
rect 44358 46084 44364 46096
rect 44319 46056 44364 46084
rect 44358 46044 44364 46056
rect 44416 46044 44422 46096
rect 45649 46087 45707 46093
rect 45649 46084 45661 46087
rect 45388 46056 45661 46084
rect 45388 46028 45416 46056
rect 45649 46053 45661 46056
rect 45695 46053 45707 46087
rect 45649 46047 45707 46053
rect 38657 46019 38715 46025
rect 38657 46016 38669 46019
rect 38580 45988 38669 46016
rect 38657 45985 38669 45988
rect 38703 45985 38715 46019
rect 45002 46016 45008 46028
rect 44963 45988 45008 46016
rect 38657 45979 38715 45985
rect 45002 45976 45008 45988
rect 45060 45976 45066 46028
rect 45370 45976 45376 46028
rect 45428 46016 45434 46028
rect 45557 46019 45615 46025
rect 45428 45988 45473 46016
rect 45428 45976 45434 45988
rect 45557 45985 45569 46019
rect 45603 46016 45615 46019
rect 46124 46016 46152 46112
rect 47302 46084 47308 46096
rect 46400 46056 47308 46084
rect 46400 46025 46428 46056
rect 47302 46044 47308 46056
rect 47360 46044 47366 46096
rect 51000 46056 51948 46084
rect 45603 45988 46152 46016
rect 46385 46019 46443 46025
rect 45603 45985 45615 45988
rect 45557 45979 45615 45985
rect 46385 45985 46397 46019
rect 46431 45985 46443 46019
rect 46658 46016 46664 46028
rect 46619 45988 46664 46016
rect 46385 45979 46443 45985
rect 46658 45976 46664 45988
rect 46716 45976 46722 46028
rect 21407 45920 23704 45948
rect 23753 45951 23811 45957
rect 21407 45917 21419 45920
rect 21361 45911 21419 45917
rect 23753 45917 23765 45951
rect 23799 45917 23811 45951
rect 23753 45911 23811 45917
rect 23569 45883 23627 45889
rect 23569 45880 23581 45883
rect 16816 45852 23581 45880
rect 16816 45840 16822 45852
rect 23569 45849 23581 45852
rect 23615 45880 23627 45883
rect 23768 45880 23796 45911
rect 24946 45908 24952 45960
rect 25004 45948 25010 45960
rect 28077 45951 28135 45957
rect 28077 45948 28089 45951
rect 25004 45920 28089 45948
rect 25004 45908 25010 45920
rect 28077 45917 28089 45920
rect 28123 45917 28135 45951
rect 28077 45911 28135 45917
rect 28813 45951 28871 45957
rect 28813 45917 28825 45951
rect 28859 45948 28871 45951
rect 28859 45920 29684 45948
rect 28859 45917 28871 45920
rect 28813 45911 28871 45917
rect 23615 45852 23796 45880
rect 23615 45849 23627 45852
rect 23569 45843 23627 45849
rect 24486 45840 24492 45892
rect 24544 45880 24550 45892
rect 29178 45880 29184 45892
rect 24544 45852 29184 45880
rect 24544 45840 24550 45852
rect 29178 45840 29184 45852
rect 29236 45840 29242 45892
rect 21177 45815 21235 45821
rect 21177 45812 21189 45815
rect 8404 45784 21189 45812
rect 21177 45781 21189 45784
rect 21223 45781 21235 45815
rect 21177 45775 21235 45781
rect 22186 45772 22192 45824
rect 22244 45812 22250 45824
rect 22281 45815 22339 45821
rect 22281 45812 22293 45815
rect 22244 45784 22293 45812
rect 22244 45772 22250 45784
rect 22281 45781 22293 45784
rect 22327 45812 22339 45815
rect 24670 45812 24676 45824
rect 22327 45784 24676 45812
rect 22327 45781 22339 45784
rect 22281 45775 22339 45781
rect 24670 45772 24676 45784
rect 24728 45812 24734 45824
rect 25317 45815 25375 45821
rect 25317 45812 25329 45815
rect 24728 45784 25329 45812
rect 24728 45772 24734 45784
rect 25317 45781 25329 45784
rect 25363 45812 25375 45815
rect 27154 45812 27160 45824
rect 25363 45784 27160 45812
rect 25363 45781 25375 45784
rect 25317 45775 25375 45781
rect 27154 45772 27160 45784
rect 27212 45772 27218 45824
rect 29656 45821 29684 45920
rect 32582 45908 32588 45960
rect 32640 45948 32646 45960
rect 32861 45951 32919 45957
rect 32861 45948 32873 45951
rect 32640 45920 32873 45948
rect 32640 45908 32646 45920
rect 32861 45917 32873 45920
rect 32907 45948 32919 45951
rect 34609 45951 34667 45957
rect 34609 45948 34621 45951
rect 32907 45920 34621 45948
rect 32907 45917 32919 45920
rect 32861 45911 32919 45917
rect 34609 45917 34621 45920
rect 34655 45948 34667 45951
rect 35434 45948 35440 45960
rect 34655 45920 35440 45948
rect 34655 45917 34667 45920
rect 34609 45911 34667 45917
rect 35434 45908 35440 45920
rect 35492 45908 35498 45960
rect 45097 45951 45155 45957
rect 38856 45920 40264 45948
rect 34974 45840 34980 45892
rect 35032 45880 35038 45892
rect 38856 45880 38884 45920
rect 40126 45880 40132 45892
rect 35032 45852 38884 45880
rect 38948 45852 40132 45880
rect 35032 45840 35038 45852
rect 29641 45815 29699 45821
rect 29641 45781 29653 45815
rect 29687 45812 29699 45815
rect 30374 45812 30380 45824
rect 29687 45784 30380 45812
rect 29687 45781 29699 45784
rect 29641 45775 29699 45781
rect 30374 45772 30380 45784
rect 30432 45772 30438 45824
rect 31941 45815 31999 45821
rect 31941 45781 31953 45815
rect 31987 45812 31999 45815
rect 38948 45812 38976 45852
rect 40126 45840 40132 45852
rect 40184 45840 40190 45892
rect 40236 45880 40264 45920
rect 45097 45917 45109 45951
rect 45143 45948 45155 45951
rect 45922 45948 45928 45960
rect 45143 45920 45928 45948
rect 45143 45917 45155 45920
rect 45097 45911 45155 45917
rect 45922 45908 45928 45920
rect 45980 45908 45986 45960
rect 46477 45951 46535 45957
rect 46477 45917 46489 45951
rect 46523 45948 46535 45951
rect 48682 45948 48688 45960
rect 46523 45920 48688 45948
rect 46523 45917 46535 45920
rect 46477 45911 46535 45917
rect 48682 45908 48688 45920
rect 48740 45908 48746 45960
rect 51000 45957 51028 46056
rect 51166 46016 51172 46028
rect 51079 45988 51172 46016
rect 51166 45976 51172 45988
rect 51224 46016 51230 46028
rect 51626 46016 51632 46028
rect 51224 45988 51632 46016
rect 51224 45976 51230 45988
rect 51626 45976 51632 45988
rect 51684 45976 51690 46028
rect 51718 45976 51724 46028
rect 51776 46016 51782 46028
rect 51920 46025 51948 46056
rect 54846 46044 54852 46096
rect 54904 46084 54910 46096
rect 55677 46087 55735 46093
rect 55677 46084 55689 46087
rect 54904 46056 55689 46084
rect 54904 46044 54910 46056
rect 55677 46053 55689 46056
rect 55723 46053 55735 46087
rect 55677 46047 55735 46053
rect 56229 46087 56287 46093
rect 56229 46053 56241 46087
rect 56275 46084 56287 46087
rect 56778 46084 56784 46096
rect 56275 46056 56784 46084
rect 56275 46053 56287 46056
rect 56229 46047 56287 46053
rect 56778 46044 56784 46056
rect 56836 46044 56842 46096
rect 61470 46044 61476 46096
rect 61528 46084 61534 46096
rect 61749 46087 61807 46093
rect 61749 46084 61761 46087
rect 61528 46056 61761 46084
rect 61528 46044 61534 46056
rect 61749 46053 61761 46056
rect 61795 46053 61807 46087
rect 61749 46047 61807 46053
rect 51905 46019 51963 46025
rect 51776 45988 51821 46016
rect 51776 45976 51782 45988
rect 51905 45985 51917 46019
rect 51951 45985 51963 46019
rect 51905 45979 51963 45985
rect 55861 46019 55919 46025
rect 55861 45985 55873 46019
rect 55907 46016 55919 46019
rect 55950 46016 55956 46028
rect 55907 45988 55956 46016
rect 55907 45985 55919 45988
rect 55861 45979 55919 45985
rect 55950 45976 55956 45988
rect 56008 45976 56014 46028
rect 62577 46019 62635 46025
rect 62577 45985 62589 46019
rect 62623 46016 62635 46019
rect 63218 46016 63224 46028
rect 62623 45988 63224 46016
rect 62623 45985 62635 45988
rect 62577 45979 62635 45985
rect 63218 45976 63224 45988
rect 63276 45976 63282 46028
rect 50985 45951 51043 45957
rect 50985 45917 50997 45951
rect 51031 45917 51043 45951
rect 62298 45948 62304 45960
rect 62259 45920 62304 45948
rect 50985 45911 51043 45917
rect 50617 45883 50675 45889
rect 50617 45880 50629 45883
rect 40236 45852 50629 45880
rect 50617 45849 50629 45852
rect 50663 45880 50675 45883
rect 50801 45883 50859 45889
rect 50801 45880 50813 45883
rect 50663 45852 50813 45880
rect 50663 45849 50675 45852
rect 50617 45843 50675 45849
rect 50801 45849 50813 45852
rect 50847 45880 50859 45883
rect 51000 45880 51028 45911
rect 62298 45908 62304 45920
rect 62356 45908 62362 45960
rect 62761 45951 62819 45957
rect 62761 45917 62773 45951
rect 62807 45917 62819 45951
rect 62761 45911 62819 45917
rect 50847 45852 51028 45880
rect 50847 45849 50859 45852
rect 50801 45843 50859 45849
rect 62022 45840 62028 45892
rect 62080 45880 62086 45892
rect 62776 45880 62804 45911
rect 62080 45852 62804 45880
rect 62080 45840 62086 45852
rect 45922 45812 45928 45824
rect 31987 45784 38976 45812
rect 45835 45784 45928 45812
rect 31987 45781 31999 45784
rect 31941 45775 31999 45781
rect 45922 45772 45928 45784
rect 45980 45812 45986 45824
rect 46474 45812 46480 45824
rect 45980 45784 46480 45812
rect 45980 45772 45986 45784
rect 46474 45772 46480 45784
rect 46532 45772 46538 45824
rect 47302 45812 47308 45824
rect 47263 45784 47308 45812
rect 47302 45772 47308 45784
rect 47360 45772 47366 45824
rect 52181 45815 52239 45821
rect 52181 45781 52193 45815
rect 52227 45812 52239 45815
rect 52638 45812 52644 45824
rect 52227 45784 52644 45812
rect 52227 45781 52239 45784
rect 52181 45775 52239 45781
rect 52638 45772 52644 45784
rect 52696 45772 52702 45824
rect 1104 45722 108008 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 65686 45722
rect 65738 45670 65750 45722
rect 65802 45670 65814 45722
rect 65866 45670 65878 45722
rect 65930 45670 96406 45722
rect 96458 45670 96470 45722
rect 96522 45670 96534 45722
rect 96586 45670 96598 45722
rect 96650 45670 108008 45722
rect 1104 45648 108008 45670
rect 27154 45568 27160 45620
rect 27212 45608 27218 45620
rect 38562 45608 38568 45620
rect 27212 45580 38568 45608
rect 27212 45568 27218 45580
rect 38562 45568 38568 45580
rect 38620 45568 38626 45620
rect 46201 45611 46259 45617
rect 46201 45577 46213 45611
rect 46247 45608 46259 45611
rect 46658 45608 46664 45620
rect 46247 45580 46664 45608
rect 46247 45577 46259 45580
rect 46201 45571 46259 45577
rect 46658 45568 46664 45580
rect 46716 45568 46722 45620
rect 54478 45568 54484 45620
rect 54536 45608 54542 45620
rect 55122 45608 55128 45620
rect 54536 45580 55128 45608
rect 54536 45568 54542 45580
rect 55122 45568 55128 45580
rect 55180 45568 55186 45620
rect 15013 45543 15071 45549
rect 15013 45509 15025 45543
rect 15059 45540 15071 45543
rect 15654 45540 15660 45552
rect 15059 45512 15660 45540
rect 15059 45509 15071 45512
rect 15013 45503 15071 45509
rect 15654 45500 15660 45512
rect 15712 45540 15718 45552
rect 44542 45540 44548 45552
rect 15712 45512 44548 45540
rect 15712 45500 15718 45512
rect 44542 45500 44548 45512
rect 44600 45500 44606 45552
rect 47670 45500 47676 45552
rect 47728 45540 47734 45552
rect 65058 45540 65064 45552
rect 47728 45512 65064 45540
rect 47728 45500 47734 45512
rect 65058 45500 65064 45512
rect 65116 45500 65122 45552
rect 2869 45475 2927 45481
rect 2869 45441 2881 45475
rect 2915 45472 2927 45475
rect 4614 45472 4620 45484
rect 2915 45444 4620 45472
rect 2915 45441 2927 45444
rect 2869 45435 2927 45441
rect 4614 45432 4620 45444
rect 4672 45432 4678 45484
rect 13446 45472 13452 45484
rect 13407 45444 13452 45472
rect 13446 45432 13452 45444
rect 13504 45472 13510 45484
rect 15197 45475 15255 45481
rect 15197 45472 15209 45475
rect 13504 45444 15209 45472
rect 13504 45432 13510 45444
rect 15197 45441 15209 45444
rect 15243 45472 15255 45475
rect 15470 45472 15476 45484
rect 15243 45444 15476 45472
rect 15243 45441 15255 45444
rect 15197 45435 15255 45441
rect 15470 45432 15476 45444
rect 15528 45432 15534 45484
rect 30834 45432 30840 45484
rect 30892 45472 30898 45484
rect 31021 45475 31079 45481
rect 31021 45472 31033 45475
rect 30892 45444 31033 45472
rect 30892 45432 30898 45444
rect 31021 45441 31033 45444
rect 31067 45441 31079 45475
rect 31021 45435 31079 45441
rect 32309 45475 32367 45481
rect 32309 45441 32321 45475
rect 32355 45472 32367 45475
rect 32858 45472 32864 45484
rect 32355 45444 32864 45472
rect 32355 45441 32367 45444
rect 32309 45435 32367 45441
rect 32858 45432 32864 45444
rect 32916 45432 32922 45484
rect 2590 45404 2596 45416
rect 2551 45376 2596 45404
rect 2590 45364 2596 45376
rect 2648 45364 2654 45416
rect 13725 45407 13783 45413
rect 13725 45373 13737 45407
rect 13771 45404 13783 45407
rect 13814 45404 13820 45416
rect 13771 45376 13820 45404
rect 13771 45373 13783 45376
rect 13725 45367 13783 45373
rect 13814 45364 13820 45376
rect 13872 45364 13878 45416
rect 23382 45364 23388 45416
rect 23440 45404 23446 45416
rect 30653 45407 30711 45413
rect 30653 45404 30665 45407
rect 23440 45376 30665 45404
rect 23440 45364 23446 45376
rect 30653 45373 30665 45376
rect 30699 45404 30711 45407
rect 31205 45407 31263 45413
rect 31205 45404 31217 45407
rect 30699 45376 31217 45404
rect 30699 45373 30711 45376
rect 30653 45367 30711 45373
rect 31205 45373 31217 45376
rect 31251 45373 31263 45407
rect 31205 45367 31263 45373
rect 31757 45407 31815 45413
rect 31757 45373 31769 45407
rect 31803 45404 31815 45407
rect 31846 45404 31852 45416
rect 31803 45376 31852 45404
rect 31803 45373 31815 45376
rect 31757 45367 31815 45373
rect 31846 45364 31852 45376
rect 31904 45364 31910 45416
rect 31941 45407 31999 45413
rect 31941 45373 31953 45407
rect 31987 45404 31999 45407
rect 44450 45404 44456 45416
rect 31987 45376 32628 45404
rect 44411 45376 44456 45404
rect 31987 45373 31999 45376
rect 31941 45367 31999 45373
rect 30374 45296 30380 45348
rect 30432 45336 30438 45348
rect 31956 45336 31984 45367
rect 30432 45308 31984 45336
rect 30432 45296 30438 45308
rect 2958 45228 2964 45280
rect 3016 45268 3022 45280
rect 3973 45271 4031 45277
rect 3973 45268 3985 45271
rect 3016 45240 3985 45268
rect 3016 45228 3022 45240
rect 3973 45237 3985 45240
rect 4019 45237 4031 45271
rect 4430 45268 4436 45280
rect 4391 45240 4436 45268
rect 3973 45231 4031 45237
rect 4430 45228 4436 45240
rect 4488 45228 4494 45280
rect 30834 45268 30840 45280
rect 30795 45240 30840 45268
rect 30834 45228 30840 45240
rect 30892 45228 30898 45280
rect 32600 45277 32628 45376
rect 44450 45364 44456 45376
rect 44508 45364 44514 45416
rect 46106 45404 46112 45416
rect 46067 45376 46112 45404
rect 46106 45364 46112 45376
rect 46164 45364 46170 45416
rect 51902 45404 51908 45416
rect 51863 45376 51908 45404
rect 51902 45364 51908 45376
rect 51960 45364 51966 45416
rect 51997 45407 52055 45413
rect 51997 45373 52009 45407
rect 52043 45404 52055 45407
rect 52365 45407 52423 45413
rect 52365 45404 52377 45407
rect 52043 45376 52377 45404
rect 52043 45373 52055 45376
rect 51997 45367 52055 45373
rect 52365 45373 52377 45376
rect 52411 45373 52423 45407
rect 52365 45367 52423 45373
rect 51353 45339 51411 45345
rect 51353 45336 51365 45339
rect 43456 45308 51365 45336
rect 32585 45271 32643 45277
rect 32585 45237 32597 45271
rect 32631 45268 32643 45271
rect 33870 45268 33876 45280
rect 32631 45240 33876 45268
rect 32631 45237 32643 45240
rect 32585 45231 32643 45237
rect 33870 45228 33876 45240
rect 33928 45268 33934 45280
rect 43456 45268 43484 45308
rect 51353 45305 51365 45308
rect 51399 45336 51411 45339
rect 51537 45339 51595 45345
rect 51537 45336 51549 45339
rect 51399 45308 51549 45336
rect 51399 45305 51411 45308
rect 51353 45299 51411 45305
rect 51537 45305 51549 45308
rect 51583 45336 51595 45339
rect 52012 45336 52040 45367
rect 52454 45364 52460 45416
rect 52512 45404 52518 45416
rect 56045 45407 56103 45413
rect 52512 45376 52557 45404
rect 52512 45364 52518 45376
rect 56045 45373 56057 45407
rect 56091 45404 56103 45407
rect 56594 45404 56600 45416
rect 56091 45376 56600 45404
rect 56091 45373 56103 45376
rect 56045 45367 56103 45373
rect 56594 45364 56600 45376
rect 56652 45364 56658 45416
rect 58069 45407 58127 45413
rect 58069 45373 58081 45407
rect 58115 45404 58127 45407
rect 58526 45404 58532 45416
rect 58115 45376 58532 45404
rect 58115 45373 58127 45376
rect 58069 45367 58127 45373
rect 58526 45364 58532 45376
rect 58584 45364 58590 45416
rect 51583 45308 52040 45336
rect 53009 45339 53067 45345
rect 51583 45305 51595 45308
rect 51537 45299 51595 45305
rect 53009 45305 53021 45339
rect 53055 45336 53067 45339
rect 54938 45336 54944 45348
rect 53055 45308 54944 45336
rect 53055 45305 53067 45308
rect 53009 45299 53067 45305
rect 54938 45296 54944 45308
rect 54996 45296 55002 45348
rect 55858 45296 55864 45348
rect 55916 45336 55922 45348
rect 65242 45336 65248 45348
rect 55916 45308 65248 45336
rect 55916 45296 55922 45308
rect 65242 45296 65248 45308
rect 65300 45296 65306 45348
rect 33928 45240 43484 45268
rect 33928 45228 33934 45240
rect 43806 45228 43812 45280
rect 43864 45268 43870 45280
rect 44545 45271 44603 45277
rect 44545 45268 44557 45271
rect 43864 45240 44557 45268
rect 43864 45228 43870 45240
rect 44545 45237 44557 45240
rect 44591 45268 44603 45271
rect 45370 45268 45376 45280
rect 44591 45240 45376 45268
rect 44591 45237 44603 45240
rect 44545 45231 44603 45237
rect 45370 45228 45376 45240
rect 45428 45228 45434 45280
rect 51902 45228 51908 45280
rect 51960 45268 51966 45280
rect 55950 45268 55956 45280
rect 51960 45240 55956 45268
rect 51960 45228 51966 45240
rect 55950 45228 55956 45240
rect 56008 45268 56014 45280
rect 56137 45271 56195 45277
rect 56137 45268 56149 45271
rect 56008 45240 56149 45268
rect 56008 45228 56014 45240
rect 56137 45237 56149 45240
rect 56183 45237 56195 45271
rect 56137 45231 56195 45237
rect 56413 45271 56471 45277
rect 56413 45237 56425 45271
rect 56459 45268 56471 45271
rect 56594 45268 56600 45280
rect 56459 45240 56600 45268
rect 56459 45237 56471 45240
rect 56413 45231 56471 45237
rect 56594 45228 56600 45240
rect 56652 45268 56658 45280
rect 57514 45268 57520 45280
rect 56652 45240 57520 45268
rect 56652 45228 56658 45240
rect 57514 45228 57520 45240
rect 57572 45228 57578 45280
rect 57698 45228 57704 45280
rect 57756 45268 57762 45280
rect 58161 45271 58219 45277
rect 58161 45268 58173 45271
rect 57756 45240 58173 45268
rect 57756 45228 57762 45240
rect 58161 45237 58173 45240
rect 58207 45237 58219 45271
rect 58161 45231 58219 45237
rect 1104 45178 108008 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 50326 45178
rect 50378 45126 50390 45178
rect 50442 45126 50454 45178
rect 50506 45126 50518 45178
rect 50570 45126 81046 45178
rect 81098 45126 81110 45178
rect 81162 45126 81174 45178
rect 81226 45126 81238 45178
rect 81290 45126 108008 45178
rect 1104 45104 108008 45126
rect 4430 45024 4436 45076
rect 4488 45064 4494 45076
rect 4706 45064 4712 45076
rect 4488 45036 4712 45064
rect 4488 45024 4494 45036
rect 4706 45024 4712 45036
rect 4764 45064 4770 45076
rect 7190 45064 7196 45076
rect 4764 45036 7196 45064
rect 4764 45024 4770 45036
rect 5368 44937 5396 45036
rect 7190 45024 7196 45036
rect 7248 45024 7254 45076
rect 15286 45024 15292 45076
rect 15344 45064 15350 45076
rect 15344 45036 23336 45064
rect 15344 45024 15350 45036
rect 5353 44931 5411 44937
rect 5353 44897 5365 44931
rect 5399 44897 5411 44931
rect 5353 44891 5411 44897
rect 5629 44863 5687 44869
rect 5629 44829 5641 44863
rect 5675 44860 5687 44863
rect 6914 44860 6920 44872
rect 5675 44832 6920 44860
rect 5675 44829 5687 44832
rect 5629 44823 5687 44829
rect 6914 44820 6920 44832
rect 6972 44820 6978 44872
rect 23308 44860 23336 45036
rect 23382 45024 23388 45076
rect 23440 45064 23446 45076
rect 24397 45067 24455 45073
rect 24397 45064 24409 45067
rect 23440 45036 24409 45064
rect 23440 45024 23446 45036
rect 24397 45033 24409 45036
rect 24443 45033 24455 45067
rect 29178 45064 29184 45076
rect 29139 45036 29184 45064
rect 24397 45027 24455 45033
rect 29178 45024 29184 45036
rect 29236 45024 29242 45076
rect 44542 45064 44548 45076
rect 44503 45036 44548 45064
rect 44542 45024 44548 45036
rect 44600 45024 44606 45076
rect 44726 45064 44732 45076
rect 44639 45036 44732 45064
rect 44726 45024 44732 45036
rect 44784 45064 44790 45076
rect 45462 45064 45468 45076
rect 44784 45036 45468 45064
rect 44784 45024 44790 45036
rect 45462 45024 45468 45036
rect 45520 45024 45526 45076
rect 47302 45024 47308 45076
rect 47360 45064 47366 45076
rect 60918 45064 60924 45076
rect 47360 45036 60924 45064
rect 47360 45024 47366 45036
rect 60918 45024 60924 45036
rect 60976 45024 60982 45076
rect 62298 45024 62304 45076
rect 62356 45064 62362 45076
rect 62485 45067 62543 45073
rect 62485 45064 62497 45067
rect 62356 45036 62497 45064
rect 62356 45024 62362 45036
rect 62485 45033 62497 45036
rect 62531 45033 62543 45067
rect 62485 45027 62543 45033
rect 44450 44956 44456 45008
rect 44508 44996 44514 45008
rect 46109 44999 46167 45005
rect 44508 44968 45600 44996
rect 44508 44956 44514 44968
rect 23842 44888 23848 44940
rect 23900 44928 23906 44940
rect 24213 44931 24271 44937
rect 24213 44928 24225 44931
rect 23900 44900 24225 44928
rect 23900 44888 23906 44900
rect 24213 44897 24225 44900
rect 24259 44897 24271 44931
rect 24213 44891 24271 44897
rect 28997 44931 29055 44937
rect 28997 44897 29009 44931
rect 29043 44928 29055 44931
rect 29178 44928 29184 44940
rect 29043 44900 29184 44928
rect 29043 44897 29055 44900
rect 28997 44891 29055 44897
rect 29178 44888 29184 44900
rect 29236 44928 29242 44940
rect 29365 44931 29423 44937
rect 29365 44928 29377 44931
rect 29236 44900 29377 44928
rect 29236 44888 29242 44900
rect 29365 44897 29377 44900
rect 29411 44897 29423 44931
rect 44358 44928 44364 44940
rect 29365 44891 29423 44897
rect 33704 44900 44364 44928
rect 33704 44860 33732 44900
rect 44358 44888 44364 44900
rect 44416 44888 44422 44940
rect 44542 44888 44548 44940
rect 44600 44928 44606 44940
rect 44821 44931 44879 44937
rect 44821 44928 44833 44931
rect 44600 44900 44833 44928
rect 44600 44888 44606 44900
rect 44821 44897 44833 44900
rect 44867 44897 44879 44931
rect 44821 44891 44879 44897
rect 44990 44931 45048 44937
rect 44990 44897 45002 44931
rect 45036 44897 45048 44931
rect 45462 44928 45468 44940
rect 45423 44900 45468 44928
rect 44990 44891 45048 44897
rect 23308 44832 33732 44860
rect 38746 44820 38752 44872
rect 38804 44860 38810 44872
rect 38933 44863 38991 44869
rect 38933 44860 38945 44863
rect 38804 44832 38945 44860
rect 38804 44820 38810 44832
rect 38933 44829 38945 44832
rect 38979 44829 38991 44863
rect 39206 44860 39212 44872
rect 39167 44832 39212 44860
rect 38933 44823 38991 44829
rect 39206 44820 39212 44832
rect 39264 44820 39270 44872
rect 45020 44792 45048 44891
rect 45462 44888 45468 44900
rect 45520 44888 45526 44940
rect 45572 44937 45600 44968
rect 46109 44965 46121 44999
rect 46155 44996 46167 44999
rect 52273 44999 52331 45005
rect 52273 44996 52285 44999
rect 46155 44968 52285 44996
rect 46155 44965 46167 44968
rect 46109 44959 46167 44965
rect 52273 44965 52285 44968
rect 52319 44965 52331 44999
rect 52273 44959 52331 44965
rect 60185 44999 60243 45005
rect 60185 44965 60197 44999
rect 60231 44996 60243 44999
rect 61562 44996 61568 45008
rect 60231 44968 61568 44996
rect 60231 44965 60243 44968
rect 60185 44959 60243 44965
rect 61562 44956 61568 44968
rect 61620 44956 61626 45008
rect 63589 44999 63647 45005
rect 63589 44996 63601 44999
rect 62592 44968 63601 44996
rect 45557 44931 45615 44937
rect 45557 44897 45569 44931
rect 45603 44928 45615 44931
rect 46842 44928 46848 44940
rect 45603 44900 46848 44928
rect 45603 44897 45615 44900
rect 45557 44891 45615 44897
rect 46842 44888 46848 44900
rect 46900 44888 46906 44940
rect 55858 44928 55864 44940
rect 46952 44900 55864 44928
rect 46385 44863 46443 44869
rect 46385 44829 46397 44863
rect 46431 44860 46443 44863
rect 46566 44860 46572 44872
rect 46431 44832 46572 44860
rect 46431 44829 46443 44832
rect 46385 44823 46443 44829
rect 46400 44792 46428 44823
rect 46566 44820 46572 44832
rect 46624 44860 46630 44872
rect 46952 44860 46980 44900
rect 55858 44888 55864 44900
rect 55916 44888 55922 44940
rect 57698 44928 57704 44940
rect 57659 44900 57704 44928
rect 57698 44888 57704 44900
rect 57756 44888 57762 44940
rect 60366 44928 60372 44940
rect 60327 44900 60372 44928
rect 60366 44888 60372 44900
rect 60424 44888 60430 44940
rect 61746 44928 61752 44940
rect 61707 44900 61752 44928
rect 61746 44888 61752 44900
rect 61804 44888 61810 44940
rect 62592 44937 62620 44968
rect 63589 44965 63601 44968
rect 63635 44996 63647 44999
rect 65518 44996 65524 45008
rect 63635 44968 65524 44996
rect 63635 44965 63647 44968
rect 63589 44959 63647 44965
rect 65518 44956 65524 44968
rect 65576 44956 65582 45008
rect 62577 44931 62635 44937
rect 62577 44897 62589 44931
rect 62623 44897 62635 44931
rect 62577 44891 62635 44897
rect 62945 44931 63003 44937
rect 62945 44897 62957 44931
rect 62991 44897 63003 44931
rect 62945 44891 63003 44897
rect 52638 44860 52644 44872
rect 46624 44832 46980 44860
rect 47044 44832 52500 44860
rect 52599 44832 52644 44860
rect 46624 44820 46630 44832
rect 45020 44764 46428 44792
rect 46474 44752 46480 44804
rect 46532 44792 46538 44804
rect 47044 44792 47072 44832
rect 46532 44764 47072 44792
rect 46532 44752 46538 44764
rect 47118 44752 47124 44804
rect 47176 44792 47182 44804
rect 51718 44792 51724 44804
rect 47176 44764 51724 44792
rect 47176 44752 47182 44764
rect 51718 44752 51724 44764
rect 51776 44752 51782 44804
rect 52472 44792 52500 44832
rect 52638 44820 52644 44832
rect 52696 44820 52702 44872
rect 57330 44820 57336 44872
rect 57388 44860 57394 44872
rect 57425 44863 57483 44869
rect 57425 44860 57437 44863
rect 57388 44832 57437 44860
rect 57388 44820 57394 44832
rect 57425 44829 57437 44832
rect 57471 44860 57483 44863
rect 59170 44860 59176 44872
rect 57471 44832 59176 44860
rect 57471 44829 57483 44832
rect 57425 44823 57483 44829
rect 59170 44820 59176 44832
rect 59228 44860 59234 44872
rect 59228 44832 59308 44860
rect 59228 44820 59234 44832
rect 57238 44792 57244 44804
rect 52472 44764 57244 44792
rect 57238 44752 57244 44764
rect 57296 44752 57302 44804
rect 59280 44801 59308 44832
rect 60734 44820 60740 44872
rect 60792 44860 60798 44872
rect 62022 44860 62028 44872
rect 60792 44832 62028 44860
rect 60792 44820 60798 44832
rect 62022 44820 62028 44832
rect 62080 44860 62086 44872
rect 62960 44860 62988 44891
rect 63218 44860 63224 44872
rect 62080 44832 62988 44860
rect 63179 44832 63224 44860
rect 62080 44820 62086 44832
rect 63218 44820 63224 44832
rect 63276 44820 63282 44872
rect 64322 44820 64328 44872
rect 64380 44860 64386 44872
rect 66625 44863 66683 44869
rect 66625 44860 66637 44863
rect 64380 44832 66637 44860
rect 64380 44820 64386 44832
rect 66625 44829 66637 44832
rect 66671 44860 66683 44863
rect 66717 44863 66775 44869
rect 66717 44860 66729 44863
rect 66671 44832 66729 44860
rect 66671 44829 66683 44832
rect 66625 44823 66683 44829
rect 66717 44829 66729 44832
rect 66763 44829 66775 44863
rect 66717 44823 66775 44829
rect 66898 44820 66904 44872
rect 66956 44860 66962 44872
rect 66993 44863 67051 44869
rect 66993 44860 67005 44863
rect 66956 44832 67005 44860
rect 66956 44820 66962 44832
rect 66993 44829 67005 44832
rect 67039 44829 67051 44863
rect 66993 44823 67051 44829
rect 59265 44795 59323 44801
rect 59265 44761 59277 44795
rect 59311 44792 59323 44795
rect 61565 44795 61623 44801
rect 61565 44792 61577 44795
rect 59311 44764 61577 44792
rect 59311 44761 59323 44764
rect 59265 44755 59323 44761
rect 61565 44761 61577 44764
rect 61611 44792 61623 44795
rect 62942 44792 62948 44804
rect 61611 44764 62948 44792
rect 61611 44761 61623 44764
rect 61565 44755 61623 44761
rect 62942 44752 62948 44764
rect 63000 44792 63006 44804
rect 64340 44792 64368 44820
rect 63000 44764 64368 44792
rect 63000 44752 63006 44764
rect 6917 44727 6975 44733
rect 6917 44693 6929 44727
rect 6963 44724 6975 44727
rect 7006 44724 7012 44736
rect 6963 44696 7012 44724
rect 6963 44693 6975 44696
rect 6917 44687 6975 44693
rect 7006 44684 7012 44696
rect 7064 44684 7070 44736
rect 23842 44684 23848 44736
rect 23900 44724 23906 44736
rect 24029 44727 24087 44733
rect 24029 44724 24041 44727
rect 23900 44696 24041 44724
rect 23900 44684 23906 44696
rect 24029 44693 24041 44696
rect 24075 44693 24087 44727
rect 38746 44724 38752 44736
rect 38707 44696 38752 44724
rect 24029 44687 24087 44693
rect 38746 44684 38752 44696
rect 38804 44684 38810 44736
rect 40494 44724 40500 44736
rect 40455 44696 40500 44724
rect 40494 44684 40500 44696
rect 40552 44684 40558 44736
rect 52454 44733 52460 44736
rect 52438 44727 52460 44733
rect 52438 44693 52450 44727
rect 52438 44687 52460 44693
rect 52454 44684 52460 44687
rect 52512 44684 52518 44736
rect 52546 44684 52552 44736
rect 52604 44724 52610 44736
rect 52917 44727 52975 44733
rect 52604 44696 52649 44724
rect 52604 44684 52610 44696
rect 52917 44693 52929 44727
rect 52963 44724 52975 44727
rect 54570 44724 54576 44736
rect 52963 44696 54576 44724
rect 52963 44693 52975 44696
rect 52917 44687 52975 44693
rect 54570 44684 54576 44696
rect 54628 44684 54634 44736
rect 58989 44727 59047 44733
rect 58989 44693 59001 44727
rect 59035 44724 59047 44727
rect 59078 44724 59084 44736
rect 59035 44696 59084 44724
rect 59035 44693 59047 44696
rect 58989 44687 59047 44693
rect 59078 44684 59084 44696
rect 59136 44684 59142 44736
rect 60458 44724 60464 44736
rect 60419 44696 60464 44724
rect 60458 44684 60464 44696
rect 60516 44684 60522 44736
rect 68281 44727 68339 44733
rect 68281 44693 68293 44727
rect 68327 44724 68339 44727
rect 68554 44724 68560 44736
rect 68327 44696 68560 44724
rect 68327 44693 68339 44696
rect 68281 44687 68339 44693
rect 68554 44684 68560 44696
rect 68612 44684 68618 44736
rect 1104 44634 108008 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 65686 44634
rect 65738 44582 65750 44634
rect 65802 44582 65814 44634
rect 65866 44582 65878 44634
rect 65930 44582 96406 44634
rect 96458 44582 96470 44634
rect 96522 44582 96534 44634
rect 96586 44582 96598 44634
rect 96650 44582 108008 44634
rect 1104 44560 108008 44582
rect 4433 44523 4491 44529
rect 4433 44489 4445 44523
rect 4479 44520 4491 44523
rect 4706 44520 4712 44532
rect 4479 44492 4712 44520
rect 4479 44489 4491 44492
rect 4433 44483 4491 44489
rect 4706 44480 4712 44492
rect 4764 44480 4770 44532
rect 7834 44480 7840 44532
rect 7892 44520 7898 44532
rect 27433 44523 27491 44529
rect 27433 44520 27445 44523
rect 7892 44492 27445 44520
rect 7892 44480 7898 44492
rect 27433 44489 27445 44492
rect 27479 44489 27491 44523
rect 27433 44483 27491 44489
rect 33689 44523 33747 44529
rect 33689 44489 33701 44523
rect 33735 44520 33747 44523
rect 39206 44520 39212 44532
rect 33735 44492 39212 44520
rect 33735 44489 33747 44492
rect 33689 44483 33747 44489
rect 39206 44480 39212 44492
rect 39264 44480 39270 44532
rect 41509 44523 41567 44529
rect 41509 44489 41521 44523
rect 41555 44520 41567 44523
rect 56778 44520 56784 44532
rect 41555 44492 56784 44520
rect 41555 44489 41567 44492
rect 41509 44483 41567 44489
rect 15286 44452 15292 44464
rect 15247 44424 15292 44452
rect 15286 44412 15292 44424
rect 15344 44412 15350 44464
rect 15470 44452 15476 44464
rect 15431 44424 15476 44452
rect 15470 44412 15476 44424
rect 15528 44412 15534 44464
rect 32309 44455 32367 44461
rect 32309 44452 32321 44455
rect 24780 44424 32321 44452
rect 24780 44396 24808 44424
rect 31956 44396 31984 44424
rect 32309 44421 32321 44424
rect 32355 44452 32367 44455
rect 32355 44424 32536 44452
rect 32355 44421 32367 44424
rect 32309 44415 32367 44421
rect 24762 44384 24768 44396
rect 13372 44356 24768 44384
rect 2590 44316 2596 44328
rect 2551 44288 2596 44316
rect 2590 44276 2596 44288
rect 2648 44276 2654 44328
rect 2869 44319 2927 44325
rect 2869 44285 2881 44319
rect 2915 44316 2927 44319
rect 6730 44316 6736 44328
rect 2915 44288 6736 44316
rect 2915 44285 2927 44288
rect 2869 44279 2927 44285
rect 6730 44276 6736 44288
rect 6788 44276 6794 44328
rect 7653 44319 7711 44325
rect 7653 44285 7665 44319
rect 7699 44285 7711 44319
rect 7653 44279 7711 44285
rect 7929 44319 7987 44325
rect 7929 44285 7941 44319
rect 7975 44316 7987 44319
rect 8938 44316 8944 44328
rect 7975 44288 8944 44316
rect 7975 44285 7987 44288
rect 7929 44279 7987 44285
rect 2866 44140 2872 44192
rect 2924 44180 2930 44192
rect 3973 44183 4031 44189
rect 3973 44180 3985 44183
rect 2924 44152 3985 44180
rect 2924 44140 2930 44152
rect 3973 44149 3985 44152
rect 4019 44149 4031 44183
rect 3973 44143 4031 44149
rect 4614 44140 4620 44192
rect 4672 44180 4678 44192
rect 7668 44180 7696 44279
rect 8938 44276 8944 44288
rect 8996 44276 9002 44328
rect 9030 44276 9036 44328
rect 9088 44316 9094 44328
rect 13372 44316 13400 44356
rect 24762 44344 24768 44356
rect 24820 44344 24826 44396
rect 27893 44387 27951 44393
rect 27893 44353 27905 44387
rect 27939 44384 27951 44387
rect 28721 44387 28779 44393
rect 28721 44384 28733 44387
rect 27939 44356 28733 44384
rect 27939 44353 27951 44356
rect 27893 44347 27951 44353
rect 28721 44353 28733 44356
rect 28767 44384 28779 44387
rect 28767 44356 31800 44384
rect 28767 44353 28779 44356
rect 28721 44347 28779 44353
rect 9088 44288 13400 44316
rect 9088 44276 9094 44288
rect 13446 44276 13452 44328
rect 13504 44316 13510 44328
rect 13725 44319 13783 44325
rect 13725 44316 13737 44319
rect 13504 44288 13737 44316
rect 13504 44276 13510 44288
rect 13725 44285 13737 44288
rect 13771 44285 13783 44319
rect 13998 44316 14004 44328
rect 13959 44288 14004 44316
rect 13725 44279 13783 44285
rect 13998 44276 14004 44288
rect 14056 44276 14062 44328
rect 18693 44319 18751 44325
rect 18693 44285 18705 44319
rect 18739 44285 18751 44319
rect 18966 44316 18972 44328
rect 18927 44288 18972 44316
rect 18693 44279 18751 44285
rect 9309 44251 9367 44257
rect 9309 44217 9321 44251
rect 9355 44248 9367 44251
rect 9674 44248 9680 44260
rect 9355 44220 9680 44248
rect 9355 44217 9367 44220
rect 9309 44211 9367 44217
rect 9674 44208 9680 44220
rect 9732 44208 9738 44260
rect 9401 44183 9459 44189
rect 9401 44180 9413 44183
rect 4672 44152 9413 44180
rect 4672 44140 4678 44152
rect 9401 44149 9413 44152
rect 9447 44149 9459 44183
rect 18708 44180 18736 44279
rect 18966 44276 18972 44288
rect 19024 44276 19030 44328
rect 22646 44276 22652 44328
rect 22704 44316 22710 44328
rect 27798 44316 27804 44328
rect 22704 44288 27804 44316
rect 22704 44276 22710 44288
rect 27798 44276 27804 44288
rect 27856 44276 27862 44328
rect 28169 44319 28227 44325
rect 28169 44285 28181 44319
rect 28215 44285 28227 44319
rect 28169 44279 28227 44285
rect 28353 44319 28411 44325
rect 28353 44285 28365 44319
rect 28399 44285 28411 44319
rect 28353 44279 28411 44285
rect 20349 44251 20407 44257
rect 20349 44217 20361 44251
rect 20395 44248 20407 44251
rect 20898 44248 20904 44260
rect 20395 44220 20904 44248
rect 20395 44217 20407 44220
rect 20349 44211 20407 44217
rect 20898 44208 20904 44220
rect 20956 44208 20962 44260
rect 21082 44208 21088 44260
rect 21140 44248 21146 44260
rect 21910 44248 21916 44260
rect 21140 44220 21916 44248
rect 21140 44208 21146 44220
rect 21910 44208 21916 44220
rect 21968 44248 21974 44260
rect 28184 44248 28212 44279
rect 28258 44248 28264 44260
rect 21968 44220 28264 44248
rect 21968 44208 21974 44220
rect 28258 44208 28264 44220
rect 28316 44208 28322 44260
rect 28368 44248 28396 44279
rect 28537 44251 28595 44257
rect 28537 44248 28549 44251
rect 28368 44220 28549 44248
rect 28537 44217 28549 44220
rect 28583 44248 28595 44251
rect 28994 44248 29000 44260
rect 28583 44220 29000 44248
rect 28583 44217 28595 44220
rect 28537 44211 28595 44217
rect 28994 44208 29000 44220
rect 29052 44208 29058 44260
rect 31772 44248 31800 44356
rect 31938 44344 31944 44396
rect 31996 44344 32002 44396
rect 32508 44393 32536 44424
rect 32493 44387 32551 44393
rect 32493 44353 32505 44387
rect 32539 44353 32551 44387
rect 32493 44347 32551 44353
rect 34057 44387 34115 44393
rect 34057 44353 34069 44387
rect 34103 44384 34115 44387
rect 41524 44384 41552 44483
rect 56778 44480 56784 44492
rect 56836 44480 56842 44532
rect 58526 44520 58532 44532
rect 58487 44492 58532 44520
rect 58526 44480 58532 44492
rect 58584 44480 58590 44532
rect 60458 44480 60464 44532
rect 60516 44520 60522 44532
rect 60599 44523 60657 44529
rect 60599 44520 60611 44523
rect 60516 44492 60611 44520
rect 60516 44480 60522 44492
rect 60599 44489 60611 44492
rect 60645 44489 60657 44523
rect 60599 44483 60657 44489
rect 60734 44480 60740 44532
rect 60792 44520 60798 44532
rect 60918 44520 60924 44532
rect 60792 44492 60837 44520
rect 60879 44492 60924 44520
rect 60792 44480 60798 44492
rect 60918 44480 60924 44492
rect 60976 44480 60982 44532
rect 65242 44520 65248 44532
rect 65203 44492 65248 44520
rect 65242 44480 65248 44492
rect 65300 44520 65306 44532
rect 65978 44520 65984 44532
rect 65300 44492 65984 44520
rect 65300 44480 65306 44492
rect 65978 44480 65984 44492
rect 66036 44480 66042 44532
rect 71314 44480 71320 44532
rect 71372 44520 71378 44532
rect 73614 44520 73620 44532
rect 71372 44492 73620 44520
rect 71372 44480 71378 44492
rect 73614 44480 73620 44492
rect 73672 44480 73678 44532
rect 44358 44412 44364 44464
rect 44416 44452 44422 44464
rect 45462 44452 45468 44464
rect 44416 44424 45468 44452
rect 44416 44412 44422 44424
rect 45462 44412 45468 44424
rect 45520 44452 45526 44464
rect 45741 44455 45799 44461
rect 45741 44452 45753 44455
rect 45520 44424 45753 44452
rect 45520 44412 45526 44424
rect 45741 44421 45753 44424
rect 45787 44452 45799 44455
rect 47670 44452 47676 44464
rect 45787 44424 46152 44452
rect 45787 44421 45799 44424
rect 45741 44415 45799 44421
rect 46124 44393 46152 44424
rect 46308 44424 47676 44452
rect 34103 44356 41552 44384
rect 46109 44387 46167 44393
rect 34103 44353 34115 44356
rect 34057 44347 34115 44353
rect 46109 44353 46121 44387
rect 46155 44353 46167 44387
rect 46109 44347 46167 44353
rect 31846 44276 31852 44328
rect 31904 44316 31910 44328
rect 32677 44319 32735 44325
rect 32677 44316 32689 44319
rect 31904 44288 32689 44316
rect 31904 44276 31910 44288
rect 32677 44285 32689 44288
rect 32723 44316 32735 44319
rect 32858 44316 32864 44328
rect 32723 44288 32864 44316
rect 32723 44285 32735 44288
rect 32677 44279 32735 44285
rect 32858 44276 32864 44288
rect 32916 44316 32922 44328
rect 33229 44319 33287 44325
rect 33229 44316 33241 44319
rect 32916 44288 33241 44316
rect 32916 44276 32922 44288
rect 33229 44285 33241 44288
rect 33275 44285 33287 44319
rect 33229 44279 33287 44285
rect 33413 44319 33471 44325
rect 33413 44285 33425 44319
rect 33459 44316 33471 44319
rect 34072 44316 34100 44347
rect 33459 44288 34100 44316
rect 33459 44285 33471 44288
rect 33413 44279 33471 44285
rect 33428 44248 33456 44279
rect 40494 44276 40500 44328
rect 40552 44316 40558 44328
rect 46308 44325 46336 44424
rect 47670 44412 47676 44424
rect 47728 44412 47734 44464
rect 52822 44452 52828 44464
rect 52104 44424 52828 44452
rect 51718 44384 51724 44396
rect 51679 44356 51724 44384
rect 51718 44344 51724 44356
rect 51776 44344 51782 44396
rect 41417 44319 41475 44325
rect 41417 44316 41429 44319
rect 40552 44288 41429 44316
rect 40552 44276 40558 44288
rect 41417 44285 41429 44288
rect 41463 44316 41475 44319
rect 45925 44319 45983 44325
rect 45925 44316 45937 44319
rect 41463 44288 45937 44316
rect 41463 44285 41475 44288
rect 41417 44279 41475 44285
rect 45925 44285 45937 44288
rect 45971 44285 45983 44319
rect 45925 44279 45983 44285
rect 46293 44319 46351 44325
rect 46293 44285 46305 44319
rect 46339 44285 46351 44319
rect 46293 44279 46351 44285
rect 46753 44319 46811 44325
rect 46753 44285 46765 44319
rect 46799 44285 46811 44319
rect 46753 44279 46811 44285
rect 46768 44248 46796 44279
rect 46842 44276 46848 44328
rect 46900 44316 46906 44328
rect 46900 44288 46945 44316
rect 46900 44276 46906 44288
rect 51258 44276 51264 44328
rect 51316 44316 51322 44328
rect 51902 44316 51908 44328
rect 51316 44288 51908 44316
rect 51316 44276 51322 44288
rect 51902 44276 51908 44288
rect 51960 44276 51966 44328
rect 31772 44220 33456 44248
rect 45572 44220 46796 44248
rect 47397 44251 47455 44257
rect 20533 44183 20591 44189
rect 20533 44180 20545 44183
rect 18708 44152 20545 44180
rect 9401 44143 9459 44149
rect 20533 44149 20545 44152
rect 20579 44180 20591 44183
rect 21818 44180 21824 44192
rect 20579 44152 21824 44180
rect 20579 44149 20591 44152
rect 20533 44143 20591 44149
rect 21818 44140 21824 44152
rect 21876 44140 21882 44192
rect 28276 44180 28304 44208
rect 45572 44192 45600 44220
rect 47397 44217 47409 44251
rect 47443 44248 47455 44251
rect 52104 44248 52132 44424
rect 52822 44412 52828 44424
rect 52880 44412 52886 44464
rect 59817 44455 59875 44461
rect 59817 44421 59829 44455
rect 59863 44452 59875 44455
rect 66070 44452 66076 44464
rect 59863 44424 66076 44452
rect 59863 44421 59875 44424
rect 59817 44415 59875 44421
rect 57238 44344 57244 44396
rect 57296 44384 57302 44396
rect 58989 44387 59047 44393
rect 58989 44384 59001 44387
rect 57296 44356 59001 44384
rect 57296 44344 57302 44356
rect 58989 44353 59001 44356
rect 59035 44384 59047 44387
rect 59832 44384 59860 44415
rect 66070 44412 66076 44424
rect 66128 44412 66134 44464
rect 66162 44412 66168 44464
rect 66220 44452 66226 44464
rect 71406 44452 71412 44464
rect 66220 44424 71412 44452
rect 66220 44412 66226 44424
rect 71406 44412 71412 44424
rect 71464 44412 71470 44464
rect 59035 44356 59860 44384
rect 59035 44353 59047 44356
rect 58989 44347 59047 44353
rect 60734 44344 60740 44396
rect 60792 44384 60798 44396
rect 60829 44387 60887 44393
rect 60829 44384 60841 44387
rect 60792 44356 60841 44384
rect 60792 44344 60798 44356
rect 60829 44353 60841 44356
rect 60875 44353 60887 44387
rect 60829 44347 60887 44353
rect 65978 44344 65984 44396
rect 66036 44384 66042 44396
rect 66036 44356 66760 44384
rect 66036 44344 66042 44356
rect 52365 44319 52423 44325
rect 52365 44285 52377 44319
rect 52411 44285 52423 44319
rect 52365 44279 52423 44285
rect 52457 44319 52515 44325
rect 52457 44285 52469 44319
rect 52503 44285 52515 44319
rect 52457 44279 52515 44285
rect 59081 44319 59139 44325
rect 59081 44285 59093 44319
rect 59127 44316 59139 44319
rect 59170 44316 59176 44328
rect 59127 44288 59176 44316
rect 59127 44285 59139 44288
rect 59081 44279 59139 44285
rect 47443 44220 52132 44248
rect 47443 44217 47455 44220
rect 47397 44211 47455 44217
rect 29086 44180 29092 44192
rect 28276 44152 29092 44180
rect 29086 44140 29092 44152
rect 29144 44140 29150 44192
rect 45554 44180 45560 44192
rect 45515 44152 45560 44180
rect 45554 44140 45560 44152
rect 45612 44140 45618 44192
rect 45925 44183 45983 44189
rect 45925 44149 45937 44183
rect 45971 44180 45983 44183
rect 47118 44180 47124 44192
rect 45971 44152 47124 44180
rect 45971 44149 45983 44152
rect 45925 44143 45983 44149
rect 47118 44140 47124 44152
rect 47176 44140 47182 44192
rect 50706 44140 50712 44192
rect 50764 44180 50770 44192
rect 52380 44180 52408 44279
rect 50764 44152 52408 44180
rect 52472 44180 52500 44279
rect 59170 44276 59176 44288
rect 59228 44276 59234 44328
rect 59446 44316 59452 44328
rect 59407 44288 59452 44316
rect 59446 44276 59452 44288
rect 59504 44276 59510 44328
rect 59633 44319 59691 44325
rect 59633 44285 59645 44319
rect 59679 44316 59691 44319
rect 65058 44316 65064 44328
rect 59679 44288 60228 44316
rect 65019 44288 65064 44316
rect 59679 44285 59691 44288
rect 59633 44279 59691 44285
rect 60200 44260 60228 44288
rect 65058 44276 65064 44288
rect 65116 44316 65122 44328
rect 65429 44319 65487 44325
rect 65429 44316 65441 44319
rect 65116 44288 65441 44316
rect 65116 44276 65122 44288
rect 65429 44285 65441 44288
rect 65475 44285 65487 44319
rect 65429 44279 65487 44285
rect 53009 44251 53067 44257
rect 53009 44217 53021 44251
rect 53055 44248 53067 44251
rect 54662 44248 54668 44260
rect 53055 44220 54668 44248
rect 53055 44217 53067 44220
rect 53009 44211 53067 44217
rect 54662 44208 54668 44220
rect 54720 44208 54726 44260
rect 60182 44208 60188 44260
rect 60240 44248 60246 44260
rect 60461 44251 60519 44257
rect 60461 44248 60473 44251
rect 60240 44220 60473 44248
rect 60240 44208 60246 44220
rect 60461 44217 60473 44220
rect 60507 44217 60519 44251
rect 65444 44248 65472 44279
rect 65518 44276 65524 44328
rect 65576 44316 65582 44328
rect 66732 44325 66760 44356
rect 66165 44319 66223 44325
rect 66165 44316 66177 44319
rect 65576 44288 66177 44316
rect 65576 44276 65582 44288
rect 66165 44285 66177 44288
rect 66211 44316 66223 44319
rect 66717 44319 66775 44325
rect 66211 44288 66484 44316
rect 66211 44285 66223 44288
rect 66165 44279 66223 44285
rect 66456 44248 66484 44288
rect 66717 44285 66729 44319
rect 66763 44285 66775 44319
rect 66990 44316 66996 44328
rect 66951 44288 66996 44316
rect 66717 44279 66775 44285
rect 66990 44276 66996 44288
rect 67048 44276 67054 44328
rect 68554 44316 68560 44328
rect 68515 44288 68560 44316
rect 68554 44276 68560 44288
rect 68612 44276 68618 44328
rect 71409 44319 71467 44325
rect 71409 44285 71421 44319
rect 71455 44285 71467 44319
rect 71409 44279 71467 44285
rect 71685 44319 71743 44325
rect 71685 44285 71697 44319
rect 71731 44316 71743 44319
rect 72878 44316 72884 44328
rect 71731 44288 72884 44316
rect 71731 44285 71743 44288
rect 71685 44279 71743 44285
rect 67361 44251 67419 44257
rect 67361 44248 67373 44251
rect 65444 44220 66392 44248
rect 66456 44220 67373 44248
rect 60461 44211 60519 44217
rect 53282 44180 53288 44192
rect 52472 44152 53288 44180
rect 50764 44140 50770 44152
rect 53282 44140 53288 44152
rect 53340 44140 53346 44192
rect 66162 44140 66168 44192
rect 66220 44180 66226 44192
rect 66257 44183 66315 44189
rect 66257 44180 66269 44183
rect 66220 44152 66269 44180
rect 66220 44140 66226 44152
rect 66257 44149 66269 44152
rect 66303 44149 66315 44183
rect 66364 44180 66392 44220
rect 67361 44217 67373 44220
rect 67407 44248 67419 44251
rect 67407 44220 68876 44248
rect 67407 44217 67419 44220
rect 67361 44211 67419 44217
rect 68649 44183 68707 44189
rect 68649 44180 68661 44183
rect 66364 44152 68661 44180
rect 66257 44143 66315 44149
rect 68649 44149 68661 44152
rect 68695 44180 68707 44183
rect 68738 44180 68744 44192
rect 68695 44152 68744 44180
rect 68695 44149 68707 44152
rect 68649 44143 68707 44149
rect 68738 44140 68744 44152
rect 68796 44140 68802 44192
rect 68848 44180 68876 44220
rect 71314 44180 71320 44192
rect 68848 44152 71320 44180
rect 71314 44140 71320 44152
rect 71372 44140 71378 44192
rect 71424 44180 71452 44279
rect 72878 44276 72884 44288
rect 72936 44276 72942 44328
rect 73157 44251 73215 44257
rect 73157 44248 73169 44251
rect 72804 44220 73169 44248
rect 72804 44180 72832 44220
rect 73157 44217 73169 44220
rect 73203 44248 73215 44251
rect 77386 44248 77392 44260
rect 73203 44220 77392 44248
rect 73203 44217 73215 44220
rect 73157 44211 73215 44217
rect 77386 44208 77392 44220
rect 77444 44208 77450 44260
rect 72970 44180 72976 44192
rect 71424 44152 72832 44180
rect 72931 44152 72976 44180
rect 72970 44140 72976 44152
rect 73028 44140 73034 44192
rect 1104 44090 108008 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 81046 44090
rect 81098 44038 81110 44090
rect 81162 44038 81174 44090
rect 81226 44038 81238 44090
rect 81290 44038 108008 44090
rect 1104 44016 108008 44038
rect 6914 43976 6920 43988
rect 6875 43948 6920 43976
rect 6914 43936 6920 43948
rect 6972 43936 6978 43988
rect 7745 43979 7803 43985
rect 7745 43945 7757 43979
rect 7791 43976 7803 43979
rect 7834 43976 7840 43988
rect 7791 43948 7840 43976
rect 7791 43945 7803 43948
rect 7745 43939 7803 43945
rect 7009 43843 7067 43849
rect 7009 43809 7021 43843
rect 7055 43840 7067 43843
rect 7098 43840 7104 43852
rect 7055 43812 7104 43840
rect 7055 43809 7067 43812
rect 7009 43803 7067 43809
rect 7098 43800 7104 43812
rect 7156 43800 7162 43852
rect 7377 43843 7435 43849
rect 7377 43809 7389 43843
rect 7423 43840 7435 43843
rect 7760 43840 7788 43939
rect 7834 43936 7840 43948
rect 7892 43936 7898 43988
rect 13814 43936 13820 43988
rect 13872 43976 13878 43988
rect 14001 43979 14059 43985
rect 14001 43976 14013 43979
rect 13872 43948 14013 43976
rect 13872 43936 13878 43948
rect 14001 43945 14013 43948
rect 14047 43945 14059 43979
rect 15654 43976 15660 43988
rect 15615 43948 15660 43976
rect 14001 43939 14059 43945
rect 15654 43936 15660 43948
rect 15712 43936 15718 43988
rect 17218 43936 17224 43988
rect 17276 43976 17282 43988
rect 27341 43979 27399 43985
rect 27341 43976 27353 43979
rect 17276 43948 27353 43976
rect 17276 43936 17282 43948
rect 27341 43945 27353 43948
rect 27387 43945 27399 43979
rect 31938 43976 31944 43988
rect 31899 43948 31944 43976
rect 27341 43939 27399 43945
rect 31938 43936 31944 43948
rect 31996 43936 32002 43988
rect 32950 43976 32956 43988
rect 32416 43948 32956 43976
rect 14274 43908 14280 43920
rect 13740 43880 14280 43908
rect 9674 43840 9680 43852
rect 7423 43812 7788 43840
rect 9635 43812 9680 43840
rect 7423 43809 7435 43812
rect 7377 43803 7435 43809
rect 9674 43800 9680 43812
rect 9732 43800 9738 43852
rect 13740 43849 13768 43880
rect 14274 43868 14280 43880
rect 14332 43908 14338 43920
rect 15381 43911 15439 43917
rect 15381 43908 15393 43911
rect 14332 43880 15393 43908
rect 14332 43868 14338 43880
rect 15381 43877 15393 43880
rect 15427 43877 15439 43911
rect 15381 43871 15439 43877
rect 12989 43843 13047 43849
rect 12989 43809 13001 43843
rect 13035 43840 13047 43843
rect 13541 43843 13599 43849
rect 13541 43840 13553 43843
rect 13035 43812 13553 43840
rect 13035 43809 13047 43812
rect 12989 43803 13047 43809
rect 12805 43775 12863 43781
rect 12805 43741 12817 43775
rect 12851 43741 12863 43775
rect 12805 43735 12863 43741
rect 3694 43664 3700 43716
rect 3752 43704 3758 43716
rect 12710 43704 12716 43716
rect 3752 43676 12716 43704
rect 3752 43664 3758 43676
rect 12710 43664 12716 43676
rect 12768 43704 12774 43716
rect 12820 43704 12848 43735
rect 12768 43676 12848 43704
rect 12768 43664 12774 43676
rect 12894 43664 12900 43716
rect 12952 43704 12958 43716
rect 13188 43704 13216 43812
rect 13541 43809 13553 43812
rect 13587 43809 13599 43843
rect 13541 43803 13599 43809
rect 13725 43843 13783 43849
rect 13725 43809 13737 43843
rect 13771 43809 13783 43843
rect 13725 43803 13783 43809
rect 15289 43843 15347 43849
rect 15289 43809 15301 43843
rect 15335 43840 15347 43843
rect 15672 43840 15700 43936
rect 29178 43908 29184 43920
rect 27724 43880 29184 43908
rect 15335 43812 15700 43840
rect 17221 43843 17279 43849
rect 15335 43809 15347 43812
rect 15289 43803 15347 43809
rect 17221 43809 17233 43843
rect 17267 43809 17279 43843
rect 20898 43840 20904 43852
rect 20859 43812 20904 43840
rect 17221 43803 17279 43809
rect 17126 43732 17132 43784
rect 17184 43772 17190 43784
rect 17236 43772 17264 43803
rect 20898 43800 20904 43812
rect 20956 43800 20962 43852
rect 27724 43840 27752 43880
rect 29178 43868 29184 43880
rect 29236 43868 29242 43920
rect 21008 43812 27752 43840
rect 17681 43775 17739 43781
rect 17681 43772 17693 43775
rect 17184 43744 17693 43772
rect 17184 43732 17190 43744
rect 17681 43741 17693 43744
rect 17727 43772 17739 43775
rect 21008 43772 21036 43812
rect 27798 43800 27804 43852
rect 27856 43840 27862 43852
rect 27893 43843 27951 43849
rect 27893 43840 27905 43843
rect 27856 43812 27905 43840
rect 27856 43800 27862 43812
rect 27893 43809 27905 43812
rect 27939 43809 27951 43843
rect 28258 43840 28264 43852
rect 28219 43812 28264 43840
rect 27893 43803 27951 43809
rect 28258 43800 28264 43812
rect 28316 43800 28322 43852
rect 28445 43843 28503 43849
rect 28445 43809 28457 43843
rect 28491 43840 28503 43843
rect 28626 43840 28632 43852
rect 28491 43812 28632 43840
rect 28491 43809 28503 43812
rect 28445 43803 28503 43809
rect 28626 43800 28632 43812
rect 28684 43800 28690 43852
rect 31956 43840 31984 43936
rect 32030 43868 32036 43920
rect 32088 43908 32094 43920
rect 32416 43908 32444 43948
rect 32950 43936 32956 43948
rect 33008 43936 33014 43988
rect 34238 43936 34244 43988
rect 34296 43976 34302 43988
rect 38565 43979 38623 43985
rect 38565 43976 38577 43979
rect 34296 43948 38577 43976
rect 34296 43936 34302 43948
rect 38565 43945 38577 43948
rect 38611 43976 38623 43979
rect 45554 43976 45560 43988
rect 38611 43948 45560 43976
rect 38611 43945 38623 43948
rect 38565 43939 38623 43945
rect 45554 43936 45560 43948
rect 45612 43936 45618 43988
rect 45830 43936 45836 43988
rect 45888 43976 45894 43988
rect 46566 43976 46572 43988
rect 45888 43948 46572 43976
rect 45888 43936 45894 43948
rect 46566 43936 46572 43948
rect 46624 43936 46630 43988
rect 54110 43936 54116 43988
rect 54168 43976 54174 43988
rect 55217 43979 55275 43985
rect 55217 43976 55229 43979
rect 54168 43948 55229 43976
rect 54168 43936 54174 43948
rect 55217 43945 55229 43948
rect 55263 43945 55275 43979
rect 55217 43939 55275 43945
rect 58989 43979 59047 43985
rect 58989 43945 59001 43979
rect 59035 43976 59047 43979
rect 59446 43976 59452 43988
rect 59035 43948 59452 43976
rect 59035 43945 59047 43948
rect 58989 43939 59047 43945
rect 59446 43936 59452 43948
rect 59504 43976 59510 43988
rect 60366 43976 60372 43988
rect 59504 43948 60372 43976
rect 59504 43936 59510 43948
rect 60366 43936 60372 43948
rect 60424 43936 60430 43988
rect 60458 43936 60464 43988
rect 60516 43976 60522 43988
rect 72878 43976 72884 43988
rect 60516 43948 72648 43976
rect 72839 43948 72884 43976
rect 60516 43936 60522 43948
rect 33505 43911 33563 43917
rect 32088 43880 32444 43908
rect 32088 43868 32094 43880
rect 32416 43849 32444 43880
rect 32600 43880 33180 43908
rect 32217 43843 32275 43849
rect 32217 43840 32229 43843
rect 31956 43812 32229 43840
rect 32217 43809 32229 43812
rect 32263 43809 32275 43843
rect 32217 43803 32275 43809
rect 32401 43843 32459 43849
rect 32401 43809 32413 43843
rect 32447 43809 32459 43843
rect 32401 43803 32459 43809
rect 17727 43744 21036 43772
rect 21913 43775 21971 43781
rect 17727 43741 17739 43744
rect 17681 43735 17739 43741
rect 21913 43741 21925 43775
rect 21959 43741 21971 43775
rect 22186 43772 22192 43784
rect 22147 43744 22192 43772
rect 21913 43735 21971 43741
rect 12952 43676 17448 43704
rect 12952 43664 12958 43676
rect 9766 43636 9772 43648
rect 9727 43608 9772 43636
rect 9766 43596 9772 43608
rect 9824 43596 9830 43648
rect 17420 43645 17448 43676
rect 21928 43648 21956 43735
rect 22186 43732 22192 43744
rect 22244 43732 22250 43784
rect 27985 43775 28043 43781
rect 27985 43741 27997 43775
rect 28031 43741 28043 43775
rect 27985 43735 28043 43741
rect 28000 43704 28028 43735
rect 28994 43732 29000 43784
rect 29052 43772 29058 43784
rect 32600 43772 32628 43880
rect 32950 43840 32956 43852
rect 32911 43812 32956 43840
rect 32950 43800 32956 43812
rect 33008 43800 33014 43852
rect 33152 43849 33180 43880
rect 33505 43877 33517 43911
rect 33551 43908 33563 43911
rect 52365 43911 52423 43917
rect 33551 43880 38700 43908
rect 33551 43877 33563 43880
rect 33505 43871 33563 43877
rect 33137 43843 33195 43849
rect 33137 43809 33149 43843
rect 33183 43840 33195 43843
rect 33183 43812 33824 43840
rect 33183 43809 33195 43812
rect 33137 43803 33195 43809
rect 29052 43744 32628 43772
rect 29052 43732 29058 43744
rect 33796 43713 33824 43812
rect 36354 43800 36360 43852
rect 36412 43840 36418 43852
rect 37001 43843 37059 43849
rect 37001 43840 37013 43843
rect 36412 43812 37013 43840
rect 36412 43800 36418 43812
rect 37001 43809 37013 43812
rect 37047 43809 37059 43843
rect 38470 43840 38476 43852
rect 38431 43812 38476 43840
rect 37001 43803 37059 43809
rect 38470 43800 38476 43812
rect 38528 43800 38534 43852
rect 38672 43840 38700 43880
rect 42168 43880 51120 43908
rect 42168 43849 42196 43880
rect 39945 43843 40003 43849
rect 39945 43840 39957 43843
rect 38672 43812 39957 43840
rect 39945 43809 39957 43812
rect 39991 43809 40003 43843
rect 39945 43803 40003 43809
rect 41325 43843 41383 43849
rect 41325 43809 41337 43843
rect 41371 43840 41383 43843
rect 42153 43843 42211 43849
rect 42153 43840 42165 43843
rect 41371 43812 42165 43840
rect 41371 43809 41383 43812
rect 41325 43803 41383 43809
rect 42153 43809 42165 43812
rect 42199 43809 42211 43843
rect 42153 43803 42211 43809
rect 44542 43800 44548 43852
rect 44600 43840 44606 43852
rect 44729 43843 44787 43849
rect 44729 43840 44741 43843
rect 44600 43812 44741 43840
rect 44600 43800 44606 43812
rect 44729 43809 44741 43812
rect 44775 43809 44787 43843
rect 45278 43840 45284 43852
rect 45239 43812 45284 43840
rect 44729 43803 44787 43809
rect 39482 43732 39488 43784
rect 39540 43772 39546 43784
rect 39669 43775 39727 43781
rect 39669 43772 39681 43775
rect 39540 43744 39681 43772
rect 39540 43732 39546 43744
rect 39669 43741 39681 43744
rect 39715 43741 39727 43775
rect 39669 43735 39727 43741
rect 33781 43707 33839 43713
rect 28000 43676 28856 43704
rect 17405 43639 17463 43645
rect 17405 43605 17417 43639
rect 17451 43636 17463 43639
rect 20346 43636 20352 43648
rect 17451 43608 20352 43636
rect 17451 43605 17463 43608
rect 17405 43599 17463 43605
rect 20346 43596 20352 43608
rect 20404 43596 20410 43648
rect 20990 43636 20996 43648
rect 20951 43608 20996 43636
rect 20990 43596 20996 43608
rect 21048 43596 21054 43648
rect 21821 43639 21879 43645
rect 21821 43605 21833 43639
rect 21867 43636 21879 43639
rect 21910 43636 21916 43648
rect 21867 43608 21916 43636
rect 21867 43605 21879 43608
rect 21821 43599 21879 43605
rect 21910 43596 21916 43608
rect 21968 43636 21974 43648
rect 23382 43636 23388 43648
rect 21968 43608 23388 43636
rect 21968 43596 21974 43608
rect 23382 43596 23388 43608
rect 23440 43596 23446 43648
rect 23477 43639 23535 43645
rect 23477 43605 23489 43639
rect 23523 43636 23535 43639
rect 23658 43636 23664 43648
rect 23523 43608 23664 43636
rect 23523 43605 23535 43608
rect 23477 43599 23535 43605
rect 23658 43596 23664 43608
rect 23716 43596 23722 43648
rect 28626 43636 28632 43648
rect 28587 43608 28632 43636
rect 28626 43596 28632 43608
rect 28684 43596 28690 43648
rect 28828 43645 28856 43676
rect 33781 43673 33793 43707
rect 33827 43704 33839 43707
rect 44744 43704 44772 43803
rect 45278 43800 45284 43812
rect 45336 43800 45342 43852
rect 45830 43840 45836 43852
rect 45791 43812 45836 43840
rect 45830 43800 45836 43812
rect 45888 43800 45894 43852
rect 51092 43849 51120 43880
rect 51828 43880 52132 43908
rect 46017 43843 46075 43849
rect 46017 43809 46029 43843
rect 46063 43840 46075 43843
rect 51077 43843 51135 43849
rect 46063 43812 46244 43840
rect 46063 43809 46075 43812
rect 46017 43803 46075 43809
rect 45094 43772 45100 43784
rect 45055 43744 45100 43772
rect 45094 43732 45100 43744
rect 45152 43732 45158 43784
rect 46216 43704 46244 43812
rect 51077 43809 51089 43843
rect 51123 43809 51135 43843
rect 51258 43840 51264 43852
rect 51219 43812 51264 43840
rect 51077 43803 51135 43809
rect 51258 43800 51264 43812
rect 51316 43800 51322 43852
rect 51828 43849 51856 43880
rect 51813 43843 51871 43849
rect 51813 43809 51825 43843
rect 51859 43809 51871 43843
rect 51813 43803 51871 43809
rect 51902 43800 51908 43852
rect 51960 43840 51966 43852
rect 51997 43843 52055 43849
rect 51997 43840 52009 43843
rect 51960 43812 52009 43840
rect 51960 43800 51966 43812
rect 51997 43809 52009 43812
rect 52043 43809 52055 43843
rect 52104 43840 52132 43880
rect 52365 43877 52377 43911
rect 52411 43908 52423 43911
rect 52454 43908 52460 43920
rect 52411 43880 52460 43908
rect 52411 43877 52423 43880
rect 52365 43871 52423 43877
rect 52454 43868 52460 43880
rect 52512 43868 52518 43920
rect 52822 43868 52828 43920
rect 52880 43908 52886 43920
rect 54573 43911 54631 43917
rect 54573 43908 54585 43911
rect 52880 43880 54585 43908
rect 52880 43868 52886 43880
rect 54573 43877 54585 43880
rect 54619 43877 54631 43911
rect 59078 43908 59084 43920
rect 54573 43871 54631 43877
rect 58912 43880 59084 43908
rect 52104 43812 52684 43840
rect 51997 43803 52055 43809
rect 33827 43676 39620 43704
rect 44744 43676 46244 43704
rect 46293 43707 46351 43713
rect 33827 43673 33839 43676
rect 33781 43667 33839 43673
rect 28813 43639 28871 43645
rect 28813 43605 28825 43639
rect 28859 43636 28871 43639
rect 34238 43636 34244 43648
rect 28859 43608 34244 43636
rect 28859 43605 28871 43608
rect 28813 43599 28871 43605
rect 34238 43596 34244 43608
rect 34296 43596 34302 43648
rect 35434 43596 35440 43648
rect 35492 43636 35498 43648
rect 36817 43639 36875 43645
rect 36817 43636 36829 43639
rect 35492 43608 36829 43636
rect 35492 43596 35498 43608
rect 36817 43605 36829 43608
rect 36863 43636 36875 43639
rect 37182 43636 37188 43648
rect 36863 43608 37188 43636
rect 36863 43605 36875 43608
rect 36817 43599 36875 43605
rect 37182 43596 37188 43608
rect 37240 43636 37246 43648
rect 38746 43636 38752 43648
rect 37240 43608 38752 43636
rect 37240 43596 37246 43608
rect 38746 43596 38752 43608
rect 38804 43636 38810 43648
rect 39482 43636 39488 43648
rect 38804 43608 39488 43636
rect 38804 43596 38810 43608
rect 39482 43596 39488 43608
rect 39540 43596 39546 43648
rect 39592 43636 39620 43676
rect 46293 43673 46305 43707
rect 46339 43704 46351 43707
rect 52454 43704 52460 43716
rect 46339 43676 52460 43704
rect 46339 43673 46351 43676
rect 46293 43667 46351 43673
rect 52454 43664 52460 43676
rect 52512 43664 52518 43716
rect 52656 43713 52684 43812
rect 54662 43800 54668 43852
rect 54720 43849 54726 43852
rect 58912 43849 58940 43880
rect 59078 43868 59084 43880
rect 59136 43908 59142 43920
rect 59173 43911 59231 43917
rect 59173 43908 59185 43911
rect 59136 43880 59185 43908
rect 59136 43868 59142 43880
rect 59173 43877 59185 43880
rect 59219 43877 59231 43911
rect 59173 43871 59231 43877
rect 54720 43843 54778 43849
rect 54720 43809 54732 43843
rect 54766 43809 54778 43843
rect 54720 43803 54778 43809
rect 58897 43843 58955 43849
rect 58897 43809 58909 43843
rect 58943 43809 58955 43843
rect 60182 43840 60188 43852
rect 60143 43812 60188 43840
rect 58897 43803 58955 43809
rect 54720 43800 54726 43803
rect 60182 43800 60188 43812
rect 60240 43800 60246 43852
rect 60384 43849 60412 43936
rect 60734 43868 60740 43920
rect 60792 43908 60798 43920
rect 65978 43908 65984 43920
rect 60792 43880 61792 43908
rect 65939 43880 65984 43908
rect 60792 43868 60798 43880
rect 60369 43843 60427 43849
rect 60369 43809 60381 43843
rect 60415 43809 60427 43843
rect 60369 43803 60427 43809
rect 60550 43800 60556 43852
rect 60608 43840 60614 43852
rect 61764 43849 61792 43880
rect 65978 43868 65984 43880
rect 66036 43868 66042 43920
rect 66165 43911 66223 43917
rect 66165 43877 66177 43911
rect 66211 43908 66223 43911
rect 66898 43908 66904 43920
rect 66211 43880 66904 43908
rect 66211 43877 66223 43880
rect 66165 43871 66223 43877
rect 66898 43868 66904 43880
rect 66956 43868 66962 43920
rect 71409 43911 71467 43917
rect 71409 43877 71421 43911
rect 71455 43908 71467 43911
rect 72510 43908 72516 43920
rect 71455 43880 72516 43908
rect 71455 43877 71467 43880
rect 71409 43871 71467 43877
rect 72510 43868 72516 43880
rect 72568 43868 72574 43920
rect 61565 43843 61623 43849
rect 61565 43840 61577 43843
rect 60608 43812 61577 43840
rect 60608 43800 60614 43812
rect 61565 43809 61577 43812
rect 61611 43809 61623 43843
rect 61565 43803 61623 43809
rect 61749 43843 61807 43849
rect 61749 43809 61761 43843
rect 61795 43809 61807 43843
rect 61749 43803 61807 43809
rect 54938 43772 54944 43784
rect 54899 43744 54944 43772
rect 54938 43732 54944 43744
rect 54996 43732 55002 43784
rect 65996 43772 66024 43868
rect 66254 43800 66260 43852
rect 66312 43840 66318 43852
rect 66717 43843 66775 43849
rect 66717 43840 66729 43843
rect 66312 43812 66729 43840
rect 66312 43800 66318 43812
rect 66717 43809 66729 43812
rect 66763 43809 66775 43843
rect 66990 43840 66996 43852
rect 66951 43812 66996 43840
rect 66717 43803 66775 43809
rect 66990 43800 66996 43812
rect 67048 43800 67054 43852
rect 71590 43840 71596 43852
rect 71551 43812 71596 43840
rect 71590 43800 71596 43812
rect 71648 43800 71654 43852
rect 67177 43775 67235 43781
rect 67177 43772 67189 43775
rect 65996 43744 67189 43772
rect 67177 43741 67189 43744
rect 67223 43741 67235 43775
rect 67177 43735 67235 43741
rect 71774 43732 71780 43784
rect 71832 43772 71838 43784
rect 71869 43775 71927 43781
rect 71869 43772 71881 43775
rect 71832 43744 71881 43772
rect 71832 43732 71838 43744
rect 71869 43741 71881 43744
rect 71915 43741 71927 43775
rect 72620 43772 72648 43948
rect 72878 43936 72884 43948
rect 72936 43936 72942 43988
rect 77386 43976 77392 43988
rect 77347 43948 77392 43976
rect 77386 43936 77392 43948
rect 77444 43936 77450 43988
rect 72786 43840 72792 43852
rect 72747 43812 72792 43840
rect 72786 43800 72792 43812
rect 72844 43800 72850 43852
rect 77404 43840 77432 43936
rect 77573 43843 77631 43849
rect 77573 43840 77585 43843
rect 77404 43812 77585 43840
rect 77573 43809 77585 43812
rect 77619 43809 77631 43843
rect 79594 43840 79600 43852
rect 77573 43803 77631 43809
rect 77680 43812 79600 43840
rect 77680 43772 77708 43812
rect 79594 43800 79600 43812
rect 79652 43800 79658 43852
rect 72620 43744 77708 43772
rect 71869 43735 71927 43741
rect 77754 43732 77760 43784
rect 77812 43772 77818 43784
rect 77849 43775 77907 43781
rect 77849 43772 77861 43775
rect 77812 43744 77861 43772
rect 77812 43732 77818 43744
rect 77849 43741 77861 43744
rect 77895 43741 77907 43775
rect 77849 43735 77907 43741
rect 52641 43707 52699 43713
rect 52641 43673 52653 43707
rect 52687 43704 52699 43707
rect 53282 43704 53288 43716
rect 52687 43676 53288 43704
rect 52687 43673 52699 43676
rect 52641 43667 52699 43673
rect 53282 43664 53288 43676
rect 53340 43704 53346 43716
rect 53340 43676 59308 43704
rect 53340 43664 53346 43676
rect 42242 43636 42248 43648
rect 39592 43608 42248 43636
rect 42242 43596 42248 43608
rect 42300 43596 42306 43648
rect 44542 43596 44548 43648
rect 44600 43636 44606 43648
rect 44913 43639 44971 43645
rect 44913 43636 44925 43639
rect 44600 43608 44925 43636
rect 44600 43596 44606 43608
rect 44913 43605 44925 43608
rect 44959 43636 44971 43639
rect 45094 43636 45100 43648
rect 44959 43608 45100 43636
rect 44959 43605 44971 43608
rect 44913 43599 44971 43605
rect 45094 43596 45100 43608
rect 45152 43596 45158 43648
rect 46750 43636 46756 43648
rect 46711 43608 46756 43636
rect 46750 43596 46756 43608
rect 46808 43596 46814 43648
rect 52914 43596 52920 43648
rect 52972 43636 52978 43648
rect 54849 43639 54907 43645
rect 54849 43636 54861 43639
rect 52972 43608 54861 43636
rect 52972 43596 52978 43608
rect 54849 43605 54861 43608
rect 54895 43605 54907 43639
rect 59280 43636 59308 43676
rect 59998 43664 60004 43716
rect 60056 43704 60062 43716
rect 63218 43704 63224 43716
rect 60056 43676 63224 43704
rect 60056 43664 60062 43676
rect 60274 43636 60280 43648
rect 59280 43608 60280 43636
rect 54849 43599 54907 43605
rect 60274 43596 60280 43608
rect 60332 43596 60338 43648
rect 60458 43636 60464 43648
rect 60419 43608 60464 43636
rect 60458 43596 60464 43608
rect 60516 43596 60522 43648
rect 61856 43645 61884 43676
rect 63218 43664 63224 43676
rect 63276 43664 63282 43716
rect 61841 43639 61899 43645
rect 61841 43605 61853 43639
rect 61887 43605 61899 43639
rect 61841 43599 61899 43605
rect 79137 43639 79195 43645
rect 79137 43605 79149 43639
rect 79183 43636 79195 43639
rect 79686 43636 79692 43648
rect 79183 43608 79692 43636
rect 79183 43605 79195 43608
rect 79137 43599 79195 43605
rect 79686 43596 79692 43608
rect 79744 43596 79750 43648
rect 1104 43546 108008 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 65686 43546
rect 65738 43494 65750 43546
rect 65802 43494 65814 43546
rect 65866 43494 65878 43546
rect 65930 43494 96406 43546
rect 96458 43494 96470 43546
rect 96522 43494 96534 43546
rect 96586 43494 96598 43546
rect 96650 43494 108008 43546
rect 1104 43472 108008 43494
rect 3970 43432 3976 43444
rect 3931 43404 3976 43432
rect 3970 43392 3976 43404
rect 4028 43392 4034 43444
rect 4433 43435 4491 43441
rect 4433 43401 4445 43435
rect 4479 43432 4491 43435
rect 11606 43432 11612 43444
rect 4479 43404 11612 43432
rect 4479 43401 4491 43404
rect 4433 43395 4491 43401
rect 2869 43299 2927 43305
rect 2869 43265 2881 43299
rect 2915 43296 2927 43299
rect 4448 43296 4476 43395
rect 11606 43392 11612 43404
rect 11664 43392 11670 43444
rect 12710 43432 12716 43444
rect 12671 43404 12716 43432
rect 12710 43392 12716 43404
rect 12768 43432 12774 43444
rect 13998 43432 14004 43444
rect 12768 43404 12848 43432
rect 13959 43404 14004 43432
rect 12768 43392 12774 43404
rect 4617 43367 4675 43373
rect 4617 43333 4629 43367
rect 4663 43364 4675 43367
rect 4706 43364 4712 43376
rect 4663 43336 4712 43364
rect 4663 43333 4675 43336
rect 4617 43327 4675 43333
rect 4706 43324 4712 43336
rect 4764 43324 4770 43376
rect 8662 43364 8668 43376
rect 8036 43336 8668 43364
rect 2915 43268 4476 43296
rect 2915 43265 2927 43268
rect 2869 43259 2927 43265
rect 2590 43228 2596 43240
rect 2503 43200 2596 43228
rect 2590 43188 2596 43200
rect 2648 43188 2654 43240
rect 8036 43237 8064 43336
rect 8662 43324 8668 43336
rect 8720 43324 8726 43376
rect 8938 43364 8944 43376
rect 8899 43336 8944 43364
rect 8938 43324 8944 43336
rect 8996 43324 9002 43376
rect 12820 43305 12848 43404
rect 13998 43392 14004 43404
rect 14056 43392 14062 43444
rect 15286 43432 15292 43444
rect 15247 43404 15292 43432
rect 15286 43392 15292 43404
rect 15344 43392 15350 43444
rect 21453 43435 21511 43441
rect 18432 43404 19656 43432
rect 12805 43299 12863 43305
rect 12805 43265 12817 43299
rect 12851 43265 12863 43299
rect 12805 43259 12863 43265
rect 16574 43256 16580 43308
rect 16632 43296 16638 43308
rect 16632 43268 18276 43296
rect 16632 43256 16638 43268
rect 7837 43231 7895 43237
rect 7837 43197 7849 43231
rect 7883 43197 7895 43231
rect 7837 43191 7895 43197
rect 8021 43231 8079 43237
rect 8021 43197 8033 43231
rect 8067 43197 8079 43231
rect 8021 43191 8079 43197
rect 8481 43231 8539 43237
rect 8481 43197 8493 43231
rect 8527 43197 8539 43231
rect 8481 43191 8539 43197
rect 8573 43231 8631 43237
rect 8573 43197 8585 43231
rect 8619 43228 8631 43231
rect 8662 43228 8668 43240
rect 8619 43200 8668 43228
rect 8619 43197 8631 43200
rect 8573 43191 8631 43197
rect 2608 43092 2636 43188
rect 4706 43092 4712 43104
rect 2608 43064 4712 43092
rect 4706 43052 4712 43064
rect 4764 43052 4770 43104
rect 7558 43052 7564 43104
rect 7616 43092 7622 43104
rect 7653 43095 7711 43101
rect 7653 43092 7665 43095
rect 7616 43064 7665 43092
rect 7616 43052 7622 43064
rect 7653 43061 7665 43064
rect 7699 43092 7711 43095
rect 7852 43092 7880 43191
rect 7699 43064 7880 43092
rect 8496 43092 8524 43191
rect 8662 43188 8668 43200
rect 8720 43188 8726 43240
rect 8938 43188 8944 43240
rect 8996 43228 9002 43240
rect 12894 43228 12900 43240
rect 8996 43200 12900 43228
rect 8996 43188 9002 43200
rect 12894 43188 12900 43200
rect 12952 43188 12958 43240
rect 12989 43231 13047 43237
rect 12989 43197 13001 43231
rect 13035 43228 13047 43231
rect 13541 43231 13599 43237
rect 13541 43228 13553 43231
rect 13035 43200 13553 43228
rect 13035 43197 13047 43200
rect 12989 43191 13047 43197
rect 13541 43197 13553 43200
rect 13587 43197 13599 43231
rect 13541 43191 13599 43197
rect 13725 43231 13783 43237
rect 13725 43197 13737 43231
rect 13771 43197 13783 43231
rect 13725 43191 13783 43197
rect 15013 43231 15071 43237
rect 15013 43197 15025 43231
rect 15059 43228 15071 43231
rect 15286 43228 15292 43240
rect 15059 43200 15292 43228
rect 15059 43197 15071 43200
rect 15013 43191 15071 43197
rect 9309 43095 9367 43101
rect 9309 43092 9321 43095
rect 8496 43064 9321 43092
rect 7699 43061 7711 43064
rect 7653 43055 7711 43061
rect 9309 43061 9321 43064
rect 9355 43092 9367 43095
rect 9766 43092 9772 43104
rect 9355 43064 9772 43092
rect 9355 43061 9367 43064
rect 9309 43055 9367 43061
rect 9766 43052 9772 43064
rect 9824 43092 9830 43104
rect 10134 43092 10140 43104
rect 9824 43064 10140 43092
rect 9824 43052 9830 43064
rect 10134 43052 10140 43064
rect 10192 43052 10198 43104
rect 13556 43092 13584 43191
rect 13630 43120 13636 43172
rect 13688 43160 13694 43172
rect 13740 43160 13768 43191
rect 15286 43188 15292 43200
rect 15344 43188 15350 43240
rect 18248 43237 18276 43268
rect 18049 43231 18107 43237
rect 18049 43228 18061 43231
rect 17788 43200 18061 43228
rect 15105 43163 15163 43169
rect 15105 43160 15117 43163
rect 13688 43132 15117 43160
rect 13688 43120 13694 43132
rect 15105 43129 15117 43132
rect 15151 43129 15163 43163
rect 16574 43160 16580 43172
rect 15105 43123 15163 43129
rect 15212 43132 16580 43160
rect 15212 43092 15240 43132
rect 16574 43120 16580 43132
rect 16632 43120 16638 43172
rect 17788 43104 17816 43200
rect 18049 43197 18061 43200
rect 18095 43197 18107 43231
rect 18049 43191 18107 43197
rect 18233 43231 18291 43237
rect 18233 43197 18245 43231
rect 18279 43197 18291 43231
rect 18432 43228 18460 43404
rect 18966 43324 18972 43376
rect 19024 43364 19030 43376
rect 19628 43373 19656 43404
rect 21453 43401 21465 43435
rect 21499 43432 21511 43435
rect 22186 43432 22192 43444
rect 21499 43404 22192 43432
rect 21499 43401 21511 43404
rect 21453 43395 21511 43401
rect 22186 43392 22192 43404
rect 22244 43392 22250 43444
rect 22646 43432 22652 43444
rect 22607 43404 22652 43432
rect 22646 43392 22652 43404
rect 22704 43392 22710 43444
rect 23382 43392 23388 43444
rect 23440 43432 23446 43444
rect 25777 43435 25835 43441
rect 25777 43432 25789 43435
rect 23440 43404 25789 43432
rect 23440 43392 23446 43404
rect 25777 43401 25789 43404
rect 25823 43401 25835 43435
rect 25777 43395 25835 43401
rect 19153 43367 19211 43373
rect 19153 43364 19165 43367
rect 19024 43336 19165 43364
rect 19024 43324 19030 43336
rect 19153 43333 19165 43336
rect 19199 43333 19211 43367
rect 19153 43327 19211 43333
rect 19613 43367 19671 43373
rect 19613 43333 19625 43367
rect 19659 43364 19671 43367
rect 19886 43364 19892 43376
rect 19659 43336 19892 43364
rect 19659 43333 19671 43336
rect 19613 43327 19671 43333
rect 19886 43324 19892 43336
rect 19944 43364 19950 43376
rect 20990 43364 20996 43376
rect 19944 43336 20996 43364
rect 19944 43324 19950 43336
rect 20990 43324 20996 43336
rect 21048 43364 21054 43376
rect 24762 43364 24768 43376
rect 21048 43336 24256 43364
rect 24723 43336 24768 43364
rect 21048 43324 21054 43336
rect 24118 43296 24124 43308
rect 22296 43268 24124 43296
rect 18693 43231 18751 43237
rect 18693 43228 18705 43231
rect 18432 43200 18705 43228
rect 18233 43191 18291 43197
rect 18693 43197 18705 43200
rect 18739 43197 18751 43231
rect 18693 43191 18751 43197
rect 18785 43231 18843 43237
rect 18785 43197 18797 43231
rect 18831 43228 18843 43231
rect 20254 43228 20260 43240
rect 18831 43200 20260 43228
rect 18831 43197 18843 43200
rect 18785 43191 18843 43197
rect 18064 43160 18092 43191
rect 20254 43188 20260 43200
rect 20312 43188 20318 43240
rect 20346 43188 20352 43240
rect 20404 43228 20410 43240
rect 20441 43231 20499 43237
rect 20441 43228 20453 43231
rect 20404 43200 20453 43228
rect 20404 43188 20410 43200
rect 20441 43197 20453 43200
rect 20487 43197 20499 43231
rect 20441 43191 20499 43197
rect 20533 43231 20591 43237
rect 20533 43197 20545 43231
rect 20579 43197 20591 43231
rect 20907 43231 20965 43237
rect 20907 43228 20919 43231
rect 20533 43191 20591 43197
rect 20824 43200 20919 43228
rect 20073 43163 20131 43169
rect 20073 43160 20085 43163
rect 18064 43132 20085 43160
rect 20073 43129 20085 43132
rect 20119 43160 20131 43163
rect 20548 43160 20576 43191
rect 20824 43172 20852 43200
rect 20907 43197 20919 43200
rect 20953 43197 20965 43231
rect 20907 43191 20965 43197
rect 20993 43231 21051 43237
rect 20993 43197 21005 43231
rect 21039 43228 21051 43231
rect 22296 43228 22324 43268
rect 24118 43256 24124 43268
rect 24176 43256 24182 43308
rect 22462 43228 22468 43240
rect 21039 43200 22324 43228
rect 22423 43200 22468 43228
rect 21039 43197 21051 43200
rect 20993 43191 21051 43197
rect 22462 43188 22468 43200
rect 22520 43188 22526 43240
rect 23658 43228 23664 43240
rect 23619 43200 23664 43228
rect 23658 43188 23664 43200
rect 23716 43188 23722 43240
rect 20806 43160 20812 43172
rect 20119 43132 20576 43160
rect 20719 43132 20812 43160
rect 20119 43129 20131 43132
rect 20073 43123 20131 43129
rect 20806 43120 20812 43132
rect 20864 43160 20870 43172
rect 21821 43163 21879 43169
rect 21821 43160 21833 43163
rect 20864 43132 21833 43160
rect 20864 43120 20870 43132
rect 21821 43129 21833 43132
rect 21867 43160 21879 43163
rect 24228 43160 24256 43336
rect 24762 43324 24768 43336
rect 24820 43324 24826 43376
rect 25792 43364 25820 43395
rect 28626 43392 28632 43444
rect 28684 43432 28690 43444
rect 33318 43432 33324 43444
rect 28684 43404 33324 43432
rect 28684 43392 28690 43404
rect 33318 43392 33324 43404
rect 33376 43392 33382 43444
rect 37001 43435 37059 43441
rect 37001 43401 37013 43435
rect 37047 43432 37059 43435
rect 38378 43432 38384 43444
rect 37047 43404 38384 43432
rect 37047 43401 37059 43404
rect 37001 43395 37059 43401
rect 38378 43392 38384 43404
rect 38436 43392 38442 43444
rect 52914 43432 52920 43444
rect 52875 43404 52920 43432
rect 52914 43392 52920 43404
rect 52972 43392 52978 43444
rect 53190 43392 53196 43444
rect 53248 43432 53254 43444
rect 53469 43435 53527 43441
rect 53469 43432 53481 43435
rect 53248 43404 53481 43432
rect 53248 43392 53254 43404
rect 53469 43401 53481 43404
rect 53515 43432 53527 43435
rect 59078 43432 59084 43444
rect 53515 43404 59084 43432
rect 53515 43401 53527 43404
rect 53469 43395 53527 43401
rect 59078 43392 59084 43404
rect 59136 43392 59142 43444
rect 59538 43392 59544 43444
rect 59596 43432 59602 43444
rect 60277 43435 60335 43441
rect 60277 43432 60289 43435
rect 59596 43404 60289 43432
rect 59596 43392 59602 43404
rect 60277 43401 60289 43404
rect 60323 43401 60335 43435
rect 60277 43395 60335 43401
rect 37182 43364 37188 43376
rect 25792 43336 26004 43364
rect 37143 43336 37188 43364
rect 24780 43228 24808 43324
rect 25976 43237 26004 43336
rect 37182 43324 37188 43336
rect 37240 43364 37246 43376
rect 37737 43367 37795 43373
rect 37737 43364 37749 43367
rect 37240 43336 37749 43364
rect 37240 43324 37246 43336
rect 32766 43296 32772 43308
rect 26068 43268 32772 43296
rect 24949 43231 25007 43237
rect 24949 43228 24961 43231
rect 24780 43200 24961 43228
rect 24949 43197 24961 43200
rect 24995 43197 25007 43231
rect 24949 43191 25007 43197
rect 25961 43231 26019 43237
rect 25961 43197 25973 43231
rect 26007 43197 26019 43231
rect 25961 43191 26019 43197
rect 26068 43160 26096 43268
rect 32766 43256 32772 43268
rect 32824 43256 32830 43308
rect 35434 43296 35440 43308
rect 35395 43268 35440 43296
rect 35434 43256 35440 43268
rect 35492 43256 35498 43308
rect 26234 43228 26240 43240
rect 26195 43200 26240 43228
rect 26234 43188 26240 43200
rect 26292 43188 26298 43240
rect 32401 43231 32459 43237
rect 32401 43228 32413 43231
rect 32324 43200 32413 43228
rect 21867 43132 23796 43160
rect 24228 43132 26096 43160
rect 21867 43129 21879 43132
rect 21821 43123 21879 43129
rect 23768 43104 23796 43132
rect 32324 43104 32352 43200
rect 32401 43197 32413 43200
rect 32447 43197 32459 43231
rect 32401 43191 32459 43197
rect 32585 43231 32643 43237
rect 32585 43197 32597 43231
rect 32631 43228 32643 43231
rect 32950 43228 32956 43240
rect 32631 43200 32956 43228
rect 32631 43197 32643 43200
rect 32585 43191 32643 43197
rect 32950 43188 32956 43200
rect 33008 43188 33014 43240
rect 33137 43231 33195 43237
rect 33137 43197 33149 43231
rect 33183 43197 33195 43231
rect 33318 43228 33324 43240
rect 33231 43200 33324 43228
rect 33137 43191 33195 43197
rect 32968 43160 32996 43188
rect 33152 43160 33180 43191
rect 33318 43188 33324 43200
rect 33376 43188 33382 43240
rect 35710 43228 35716 43240
rect 35671 43200 35716 43228
rect 35710 43188 35716 43200
rect 35768 43188 35774 43240
rect 37660 43228 37688 43336
rect 37737 43333 37749 43336
rect 37783 43333 37795 43367
rect 37737 43327 37795 43333
rect 42242 43324 42248 43376
rect 42300 43364 42306 43376
rect 56594 43364 56600 43376
rect 42300 43336 56600 43364
rect 42300 43324 42306 43336
rect 56594 43324 56600 43336
rect 56652 43324 56658 43376
rect 60182 43324 60188 43376
rect 60240 43364 60246 43376
rect 60240 43336 60794 43364
rect 60240 43324 60246 43336
rect 37826 43256 37832 43308
rect 37884 43296 37890 43308
rect 44818 43296 44824 43308
rect 37884 43268 44824 43296
rect 37884 43256 37890 43268
rect 44818 43256 44824 43268
rect 44876 43256 44882 43308
rect 53006 43256 53012 43308
rect 53064 43296 53070 43308
rect 53285 43299 53343 43305
rect 53285 43296 53297 43299
rect 53064 43268 53297 43296
rect 53064 43256 53070 43268
rect 53285 43265 53297 43268
rect 53331 43296 53343 43299
rect 58710 43296 58716 43308
rect 53331 43268 58716 43296
rect 53331 43265 53343 43268
rect 53285 43259 53343 43265
rect 58710 43256 58716 43268
rect 58768 43256 58774 43308
rect 60458 43296 60464 43308
rect 58820 43268 60464 43296
rect 37921 43231 37979 43237
rect 37921 43228 37933 43231
rect 37660 43200 37933 43228
rect 37921 43197 37933 43200
rect 37967 43197 37979 43231
rect 38197 43231 38255 43237
rect 38197 43228 38209 43231
rect 37921 43191 37979 43197
rect 38028 43200 38209 43228
rect 32968 43132 33180 43160
rect 17770 43092 17776 43104
rect 13556 43064 15240 43092
rect 17731 43064 17776 43092
rect 17770 43052 17776 43064
rect 17828 43052 17834 43104
rect 17862 43052 17868 43104
rect 17920 43092 17926 43104
rect 22281 43095 22339 43101
rect 22281 43092 22293 43095
rect 17920 43064 22293 43092
rect 17920 43052 17926 43064
rect 22281 43061 22293 43064
rect 22327 43092 22339 43095
rect 22462 43092 22468 43104
rect 22327 43064 22468 43092
rect 22327 43061 22339 43064
rect 22281 43055 22339 43061
rect 22462 43052 22468 43064
rect 22520 43052 22526 43104
rect 23750 43092 23756 43104
rect 23711 43064 23756 43092
rect 23750 43052 23756 43064
rect 23808 43052 23814 43104
rect 25038 43092 25044 43104
rect 24999 43064 25044 43092
rect 25038 43052 25044 43064
rect 25096 43052 25102 43104
rect 27522 43092 27528 43104
rect 27483 43064 27528 43092
rect 27522 43052 27528 43064
rect 27580 43052 27586 43104
rect 32306 43092 32312 43104
rect 32267 43064 32312 43092
rect 32306 43052 32312 43064
rect 32364 43052 32370 43104
rect 33336 43092 33364 43188
rect 33689 43163 33747 43169
rect 33689 43129 33701 43163
rect 33735 43160 33747 43163
rect 38028 43160 38056 43200
rect 38197 43197 38209 43200
rect 38243 43197 38255 43231
rect 38197 43191 38255 43197
rect 51442 43188 51448 43240
rect 51500 43228 51506 43240
rect 51721 43231 51779 43237
rect 51721 43228 51733 43231
rect 51500 43200 51733 43228
rect 51500 43188 51506 43200
rect 51721 43197 51733 43200
rect 51767 43197 51779 43231
rect 51721 43191 51779 43197
rect 51905 43231 51963 43237
rect 51905 43197 51917 43231
rect 51951 43228 51963 43231
rect 51994 43228 52000 43240
rect 51951 43200 52000 43228
rect 51951 43197 51963 43200
rect 51905 43191 51963 43197
rect 51994 43188 52000 43200
rect 52052 43188 52058 43240
rect 52365 43231 52423 43237
rect 52365 43197 52377 43231
rect 52411 43197 52423 43231
rect 52365 43191 52423 43197
rect 52457 43231 52515 43237
rect 52457 43197 52469 43231
rect 52503 43228 52515 43231
rect 53190 43228 53196 43240
rect 52503 43200 53196 43228
rect 52503 43197 52515 43200
rect 52457 43191 52515 43197
rect 33735 43132 35572 43160
rect 33735 43129 33747 43132
rect 33689 43123 33747 43129
rect 33962 43092 33968 43104
rect 33336 43064 33968 43092
rect 33962 43052 33968 43064
rect 34020 43052 34026 43104
rect 35544 43092 35572 43132
rect 36740 43132 38056 43160
rect 36740 43092 36768 43132
rect 44818 43120 44824 43172
rect 44876 43160 44882 43172
rect 51261 43163 51319 43169
rect 51261 43160 51273 43163
rect 44876 43132 51273 43160
rect 44876 43120 44882 43132
rect 51261 43129 51273 43132
rect 51307 43160 51319 43163
rect 52380 43160 52408 43191
rect 53190 43188 53196 43200
rect 53248 43188 53254 43240
rect 58820 43237 58848 43268
rect 60458 43256 60464 43268
rect 60516 43296 60522 43308
rect 60766 43296 60794 43336
rect 71038 43324 71044 43376
rect 71096 43364 71102 43376
rect 72970 43364 72976 43376
rect 71096 43336 72976 43364
rect 71096 43324 71102 43336
rect 71593 43299 71651 43305
rect 71593 43296 71605 43299
rect 60516 43268 60596 43296
rect 60766 43268 71605 43296
rect 60516 43256 60522 43268
rect 58805 43231 58863 43237
rect 58805 43197 58817 43231
rect 58851 43197 58863 43231
rect 58805 43191 58863 43197
rect 59446 43188 59452 43240
rect 59504 43228 59510 43240
rect 59817 43231 59875 43237
rect 59817 43228 59829 43231
rect 59504 43200 59829 43228
rect 59504 43188 59510 43200
rect 59817 43197 59829 43200
rect 59863 43197 59875 43231
rect 60090 43228 60096 43240
rect 60051 43200 60096 43228
rect 59817 43191 59875 43197
rect 51307 43132 52408 43160
rect 51307 43129 51319 43132
rect 51261 43123 51319 43129
rect 39482 43092 39488 43104
rect 35544 43064 36768 43092
rect 39443 43064 39488 43092
rect 39482 43052 39488 43064
rect 39540 43052 39546 43104
rect 51442 43092 51448 43104
rect 51403 43064 51448 43092
rect 51442 43052 51448 43064
rect 51500 43052 51506 43104
rect 58897 43095 58955 43101
rect 58897 43061 58909 43095
rect 58943 43092 58955 43095
rect 59170 43092 59176 43104
rect 58943 43064 59176 43092
rect 58943 43061 58955 43064
rect 58897 43055 58955 43061
rect 59170 43052 59176 43064
rect 59228 43092 59234 43104
rect 59630 43092 59636 43104
rect 59228 43064 59636 43092
rect 59228 43052 59234 43064
rect 59630 43052 59636 43064
rect 59688 43052 59694 43104
rect 59832 43092 59860 43191
rect 60090 43188 60096 43200
rect 60148 43188 60154 43240
rect 60568 43228 60596 43268
rect 71593 43265 71605 43268
rect 71639 43265 71651 43299
rect 71593 43259 71651 43265
rect 61381 43231 61439 43237
rect 61381 43228 61393 43231
rect 60568 43200 61393 43228
rect 61381 43197 61393 43200
rect 61427 43197 61439 43231
rect 61562 43228 61568 43240
rect 61523 43200 61568 43228
rect 61381 43191 61439 43197
rect 61562 43188 61568 43200
rect 61620 43188 61626 43240
rect 66898 43228 66904 43240
rect 66859 43200 66904 43228
rect 66898 43188 66904 43200
rect 66956 43188 66962 43240
rect 67082 43188 67088 43240
rect 67140 43228 67146 43240
rect 71038 43228 71044 43240
rect 67140 43200 71044 43228
rect 67140 43188 67146 43200
rect 71038 43188 71044 43200
rect 71096 43188 71102 43240
rect 71133 43231 71191 43237
rect 71133 43197 71145 43231
rect 71179 43197 71191 43231
rect 71133 43191 71191 43197
rect 59998 43160 60004 43172
rect 59959 43132 60004 43160
rect 59998 43120 60004 43132
rect 60056 43120 60062 43172
rect 60182 43120 60188 43172
rect 60240 43160 60246 43172
rect 60550 43160 60556 43172
rect 60240 43132 60556 43160
rect 60240 43120 60246 43132
rect 60550 43120 60556 43132
rect 60608 43160 60614 43172
rect 66714 43160 66720 43172
rect 60608 43132 61700 43160
rect 66675 43132 66720 43160
rect 60608 43120 60614 43132
rect 60642 43092 60648 43104
rect 59832 43064 60648 43092
rect 60642 43052 60648 43064
rect 60700 43052 60706 43104
rect 61672 43101 61700 43132
rect 66714 43120 66720 43132
rect 66772 43120 66778 43172
rect 71148 43160 71176 43191
rect 71222 43188 71228 43240
rect 71280 43228 71286 43240
rect 71409 43231 71467 43237
rect 71280 43200 71325 43228
rect 71280 43188 71286 43200
rect 71409 43197 71421 43231
rect 71455 43228 71467 43231
rect 71866 43228 71872 43240
rect 71455 43200 71872 43228
rect 71455 43197 71467 43200
rect 71409 43191 71467 43197
rect 71866 43188 71872 43200
rect 71924 43188 71930 43240
rect 72712 43237 72740 43336
rect 72970 43324 72976 43336
rect 73028 43324 73034 43376
rect 77573 43299 77631 43305
rect 77573 43265 77585 43299
rect 77619 43296 77631 43299
rect 77754 43296 77760 43308
rect 77619 43268 77760 43296
rect 77619 43265 77631 43268
rect 77573 43259 77631 43265
rect 77754 43256 77760 43268
rect 77812 43256 77818 43308
rect 72697 43231 72755 43237
rect 72697 43197 72709 43231
rect 72743 43197 72755 43231
rect 72697 43191 72755 43197
rect 77846 43188 77852 43240
rect 77904 43228 77910 43240
rect 78125 43231 78183 43237
rect 78125 43228 78137 43231
rect 77904 43200 78137 43228
rect 77904 43188 77910 43200
rect 78125 43197 78137 43200
rect 78171 43197 78183 43231
rect 78398 43228 78404 43240
rect 78359 43200 78404 43228
rect 78125 43191 78183 43197
rect 78398 43188 78404 43200
rect 78456 43188 78462 43240
rect 78582 43228 78588 43240
rect 78543 43200 78588 43228
rect 78582 43188 78588 43200
rect 78640 43188 78646 43240
rect 71958 43160 71964 43172
rect 71148 43132 71964 43160
rect 71958 43120 71964 43132
rect 72016 43120 72022 43172
rect 61657 43095 61715 43101
rect 61657 43061 61669 43095
rect 61703 43061 61715 43095
rect 61657 43055 61715 43061
rect 66346 43052 66352 43104
rect 66404 43092 66410 43104
rect 66990 43092 66996 43104
rect 66404 43064 66996 43092
rect 66404 43052 66410 43064
rect 66990 43052 66996 43064
rect 67048 43052 67054 43104
rect 72418 43052 72424 43104
rect 72476 43092 72482 43104
rect 72789 43095 72847 43101
rect 72789 43092 72801 43095
rect 72476 43064 72801 43092
rect 72476 43052 72482 43064
rect 72789 43061 72801 43064
rect 72835 43061 72847 43095
rect 77478 43092 77484 43104
rect 77439 43064 77484 43092
rect 72789 43055 72847 43061
rect 77478 43052 77484 43064
rect 77536 43052 77542 43104
rect 1104 43002 108008 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 81046 43002
rect 81098 42950 81110 43002
rect 81162 42950 81174 43002
rect 81226 42950 81238 43002
rect 81290 42950 108008 43002
rect 1104 42928 108008 42950
rect 4062 42848 4068 42900
rect 4120 42888 4126 42900
rect 32306 42888 32312 42900
rect 4120 42860 32312 42888
rect 4120 42848 4126 42860
rect 32306 42848 32312 42860
rect 32364 42888 32370 42900
rect 32493 42891 32551 42897
rect 32493 42888 32505 42891
rect 32364 42860 32505 42888
rect 32364 42848 32370 42860
rect 32493 42857 32505 42860
rect 32539 42857 32551 42891
rect 32493 42851 32551 42857
rect 33962 42848 33968 42900
rect 34020 42888 34026 42900
rect 39025 42891 39083 42897
rect 39025 42888 39037 42891
rect 34020 42860 39037 42888
rect 34020 42848 34026 42860
rect 39025 42857 39037 42860
rect 39071 42888 39083 42891
rect 44726 42888 44732 42900
rect 39071 42860 44732 42888
rect 39071 42857 39083 42860
rect 39025 42851 39083 42857
rect 44726 42848 44732 42860
rect 44784 42848 44790 42900
rect 44818 42848 44824 42900
rect 44876 42888 44882 42900
rect 46566 42888 46572 42900
rect 44876 42860 44921 42888
rect 46527 42860 46572 42888
rect 44876 42848 44882 42860
rect 46566 42848 46572 42860
rect 46624 42848 46630 42900
rect 51169 42891 51227 42897
rect 51169 42857 51181 42891
rect 51215 42888 51227 42891
rect 51258 42888 51264 42900
rect 51215 42860 51264 42888
rect 51215 42857 51227 42860
rect 51169 42851 51227 42857
rect 51258 42848 51264 42860
rect 51316 42888 51322 42900
rect 51810 42888 51816 42900
rect 51316 42860 51816 42888
rect 51316 42848 51322 42860
rect 51810 42848 51816 42860
rect 51868 42848 51874 42900
rect 51994 42848 52000 42900
rect 52052 42888 52058 42900
rect 53006 42888 53012 42900
rect 52052 42860 53012 42888
rect 52052 42848 52058 42860
rect 53006 42848 53012 42860
rect 53064 42848 53070 42900
rect 53190 42888 53196 42900
rect 53151 42860 53196 42888
rect 53190 42848 53196 42860
rect 53248 42848 53254 42900
rect 77846 42888 77852 42900
rect 77807 42860 77852 42888
rect 77846 42848 77852 42860
rect 77904 42848 77910 42900
rect 6730 42780 6736 42832
rect 6788 42820 6794 42832
rect 7561 42823 7619 42829
rect 7561 42820 7573 42823
rect 6788 42792 7573 42820
rect 6788 42780 6794 42792
rect 7561 42789 7573 42792
rect 7607 42789 7619 42823
rect 17218 42820 17224 42832
rect 7561 42783 7619 42789
rect 7760 42792 17224 42820
rect 7098 42752 7104 42764
rect 7059 42724 7104 42752
rect 7098 42712 7104 42724
rect 7156 42712 7162 42764
rect 7760 42761 7788 42792
rect 17218 42780 17224 42792
rect 17276 42780 17282 42832
rect 23750 42780 23756 42832
rect 23808 42820 23814 42832
rect 44542 42820 44548 42832
rect 23808 42792 44548 42820
rect 23808 42780 23814 42792
rect 44542 42780 44548 42792
rect 44600 42780 44606 42832
rect 7377 42755 7435 42761
rect 7377 42721 7389 42755
rect 7423 42752 7435 42755
rect 7745 42755 7803 42761
rect 7745 42752 7757 42755
rect 7423 42724 7757 42752
rect 7423 42721 7435 42724
rect 7377 42715 7435 42721
rect 7745 42721 7757 42724
rect 7791 42721 7803 42755
rect 13722 42752 13728 42764
rect 13683 42724 13728 42752
rect 7745 42715 7803 42721
rect 13722 42712 13728 42724
rect 13780 42712 13786 42764
rect 13998 42712 14004 42764
rect 14056 42752 14062 42764
rect 14093 42755 14151 42761
rect 14093 42752 14105 42755
rect 14056 42724 14105 42752
rect 14056 42712 14062 42724
rect 14093 42721 14105 42724
rect 14139 42721 14151 42755
rect 14274 42752 14280 42764
rect 14235 42724 14280 42752
rect 14093 42715 14151 42721
rect 14274 42712 14280 42724
rect 14332 42712 14338 42764
rect 16390 42712 16396 42764
rect 16448 42752 16454 42764
rect 20901 42755 20959 42761
rect 20901 42752 20913 42755
rect 16448 42724 20913 42752
rect 16448 42712 16454 42724
rect 20901 42721 20913 42724
rect 20947 42752 20959 42755
rect 21269 42755 21327 42761
rect 21269 42752 21281 42755
rect 20947 42724 21281 42752
rect 20947 42721 20959 42724
rect 20901 42715 20959 42721
rect 21269 42721 21281 42724
rect 21315 42721 21327 42755
rect 21269 42715 21327 42721
rect 29914 42712 29920 42764
rect 29972 42752 29978 42764
rect 30837 42755 30895 42761
rect 30837 42752 30849 42755
rect 29972 42724 30849 42752
rect 29972 42712 29978 42724
rect 30837 42721 30849 42724
rect 30883 42752 30895 42755
rect 30929 42755 30987 42761
rect 30929 42752 30941 42755
rect 30883 42724 30941 42752
rect 30883 42721 30895 42724
rect 30837 42715 30895 42721
rect 30929 42721 30941 42724
rect 30975 42721 30987 42755
rect 30929 42715 30987 42721
rect 32306 42712 32312 42764
rect 32364 42752 32370 42764
rect 32677 42755 32735 42761
rect 32677 42752 32689 42755
rect 32364 42724 32689 42752
rect 32364 42712 32370 42724
rect 32677 42721 32689 42724
rect 32723 42721 32735 42755
rect 32858 42752 32864 42764
rect 32819 42724 32864 42752
rect 32677 42715 32735 42721
rect 32858 42712 32864 42724
rect 32916 42752 32922 42764
rect 33413 42755 33471 42761
rect 33413 42752 33425 42755
rect 32916 42724 33425 42752
rect 32916 42712 32922 42724
rect 33413 42721 33425 42724
rect 33459 42721 33471 42755
rect 33413 42715 33471 42721
rect 33597 42755 33655 42761
rect 33597 42721 33609 42755
rect 33643 42752 33655 42755
rect 34238 42752 34244 42764
rect 33643 42724 34244 42752
rect 33643 42721 33655 42724
rect 33597 42715 33655 42721
rect 34238 42712 34244 42724
rect 34296 42712 34302 42764
rect 38933 42755 38991 42761
rect 38933 42721 38945 42755
rect 38979 42752 38991 42755
rect 39482 42752 39488 42764
rect 38979 42724 39488 42752
rect 38979 42721 38991 42724
rect 38933 42715 38991 42721
rect 39482 42712 39488 42724
rect 39540 42712 39546 42764
rect 44358 42712 44364 42764
rect 44416 42752 44422 42764
rect 44637 42755 44695 42761
rect 44637 42752 44649 42755
rect 44416 42724 44649 42752
rect 44416 42712 44422 42724
rect 44637 42721 44649 42724
rect 44683 42721 44695 42755
rect 44836 42752 44864 42848
rect 45278 42820 45284 42832
rect 45191 42792 45284 42820
rect 45204 42761 45232 42792
rect 45278 42780 45284 42792
rect 45336 42820 45342 42832
rect 52012 42820 52040 42848
rect 45336 42792 46796 42820
rect 45336 42780 45342 42792
rect 46768 42764 46796 42792
rect 51644 42792 52040 42820
rect 45005 42755 45063 42761
rect 45005 42752 45017 42755
rect 44836 42724 45017 42752
rect 44637 42715 44695 42721
rect 45005 42721 45017 42724
rect 45051 42721 45063 42755
rect 45005 42715 45063 42721
rect 45189 42755 45247 42761
rect 45189 42721 45201 42755
rect 45235 42721 45247 42755
rect 45189 42715 45247 42721
rect 45554 42712 45560 42764
rect 45612 42752 45618 42764
rect 45649 42755 45707 42761
rect 45649 42752 45661 42755
rect 45612 42724 45661 42752
rect 45612 42712 45618 42724
rect 45649 42721 45661 42724
rect 45695 42721 45707 42755
rect 45649 42715 45707 42721
rect 45741 42755 45799 42761
rect 45741 42721 45753 42755
rect 45787 42752 45799 42755
rect 46566 42752 46572 42764
rect 45787 42724 46572 42752
rect 45787 42721 45799 42724
rect 45741 42715 45799 42721
rect 46566 42712 46572 42724
rect 46624 42712 46630 42764
rect 46750 42712 46756 42764
rect 46808 42752 46814 42764
rect 51644 42761 51672 42792
rect 51629 42755 51687 42761
rect 46808 42724 51580 42752
rect 46808 42712 46814 42724
rect 11054 42644 11060 42696
rect 11112 42684 11118 42696
rect 13081 42687 13139 42693
rect 13081 42684 13093 42687
rect 11112 42656 13093 42684
rect 11112 42644 11118 42656
rect 13081 42653 13093 42656
rect 13127 42653 13139 42687
rect 13630 42684 13636 42696
rect 13591 42656 13636 42684
rect 13081 42647 13139 42653
rect 13630 42644 13636 42656
rect 13688 42644 13694 42696
rect 33965 42687 34023 42693
rect 33965 42653 33977 42687
rect 34011 42684 34023 42687
rect 35710 42684 35716 42696
rect 34011 42656 35716 42684
rect 34011 42653 34023 42656
rect 33965 42647 34023 42653
rect 35710 42644 35716 42656
rect 35768 42644 35774 42696
rect 46124 42656 50660 42684
rect 4062 42576 4068 42628
rect 4120 42616 4126 42628
rect 30834 42616 30840 42628
rect 4120 42588 30840 42616
rect 4120 42576 4126 42588
rect 30834 42576 30840 42588
rect 30892 42576 30898 42628
rect 44542 42576 44548 42628
rect 44600 42616 44606 42628
rect 46124 42616 46152 42656
rect 44600 42588 46152 42616
rect 46201 42619 46259 42625
rect 44600 42576 44606 42588
rect 46201 42585 46213 42619
rect 46247 42616 46259 42619
rect 50632 42616 50660 42656
rect 51258 42644 51264 42696
rect 51316 42684 51322 42696
rect 51445 42687 51503 42693
rect 51445 42684 51457 42687
rect 51316 42656 51457 42684
rect 51316 42644 51322 42656
rect 51445 42653 51457 42656
rect 51491 42653 51503 42687
rect 51552 42684 51580 42724
rect 51629 42721 51641 42755
rect 51675 42721 51687 42755
rect 51629 42715 51687 42721
rect 51718 42712 51724 42764
rect 51776 42752 51782 42764
rect 52089 42755 52147 42761
rect 52089 42752 52101 42755
rect 51776 42724 52101 42752
rect 51776 42712 51782 42724
rect 52089 42721 52101 42724
rect 52135 42721 52147 42755
rect 52089 42715 52147 42721
rect 52178 42712 52184 42764
rect 52236 42752 52242 42764
rect 53208 42752 53236 42848
rect 66346 42820 66352 42832
rect 58636 42792 59032 42820
rect 66307 42792 66352 42820
rect 58636 42761 58664 42792
rect 52236 42724 53236 42752
rect 58621 42755 58679 42761
rect 52236 42712 52242 42724
rect 58621 42721 58633 42755
rect 58667 42721 58679 42755
rect 58621 42715 58679 42721
rect 58713 42755 58771 42761
rect 58713 42721 58725 42755
rect 58759 42721 58771 42755
rect 58713 42715 58771 42721
rect 58805 42755 58863 42761
rect 58805 42721 58817 42755
rect 58851 42752 58863 42755
rect 58894 42752 58900 42764
rect 58851 42724 58900 42752
rect 58851 42721 58863 42724
rect 58805 42715 58863 42721
rect 58728 42684 58756 42715
rect 58894 42712 58900 42724
rect 58952 42712 58958 42764
rect 59004 42752 59032 42792
rect 66346 42780 66352 42792
rect 66404 42780 66410 42832
rect 71590 42820 71596 42832
rect 69308 42792 71596 42820
rect 59446 42752 59452 42764
rect 59004 42724 59452 42752
rect 59446 42712 59452 42724
rect 59504 42712 59510 42764
rect 60182 42752 60188 42764
rect 60095 42724 60188 42752
rect 60182 42712 60188 42724
rect 60240 42712 60246 42764
rect 60737 42755 60795 42761
rect 60737 42752 60749 42755
rect 60660 42724 60749 42752
rect 60200 42684 60228 42712
rect 51552 42656 51856 42684
rect 58728 42656 60228 42684
rect 51445 42647 51503 42653
rect 51353 42619 51411 42625
rect 51353 42616 51365 42619
rect 46247 42588 48636 42616
rect 50632 42588 51365 42616
rect 46247 42585 46259 42588
rect 46201 42579 46259 42585
rect 21082 42548 21088 42560
rect 21043 42520 21088 42548
rect 21082 42508 21088 42520
rect 21140 42508 21146 42560
rect 31113 42551 31171 42557
rect 31113 42517 31125 42551
rect 31159 42548 31171 42551
rect 32858 42548 32864 42560
rect 31159 42520 32864 42548
rect 31159 42517 31171 42520
rect 31113 42511 31171 42517
rect 32858 42508 32864 42520
rect 32916 42508 32922 42560
rect 48608 42548 48636 42588
rect 51353 42585 51365 42588
rect 51399 42616 51411 42619
rect 51718 42616 51724 42628
rect 51399 42588 51724 42616
rect 51399 42585 51411 42588
rect 51353 42579 51411 42585
rect 51718 42576 51724 42588
rect 51776 42576 51782 42628
rect 51828 42616 51856 42656
rect 52178 42616 52184 42628
rect 51828 42588 52184 42616
rect 52178 42576 52184 42588
rect 52236 42576 52242 42628
rect 52546 42616 52552 42628
rect 52507 42588 52552 42616
rect 52546 42576 52552 42588
rect 52604 42576 52610 42628
rect 58728 42588 59124 42616
rect 51166 42548 51172 42560
rect 48608 42520 51172 42548
rect 51166 42508 51172 42520
rect 51224 42508 51230 42560
rect 52270 42508 52276 42560
rect 52328 42548 52334 42560
rect 58728 42548 58756 42588
rect 52328 42520 58756 42548
rect 52328 42508 52334 42520
rect 58802 42508 58808 42560
rect 58860 42548 58866 42560
rect 58989 42551 59047 42557
rect 58989 42548 59001 42551
rect 58860 42520 59001 42548
rect 58860 42508 58866 42520
rect 58989 42517 59001 42520
rect 59035 42517 59047 42551
rect 59096 42548 59124 42588
rect 60090 42576 60096 42628
rect 60148 42616 60154 42628
rect 60277 42619 60335 42625
rect 60277 42616 60289 42619
rect 60148 42588 60289 42616
rect 60148 42576 60154 42588
rect 60277 42585 60289 42588
rect 60323 42585 60335 42619
rect 60277 42579 60335 42585
rect 60660 42548 60688 42724
rect 60737 42721 60749 42724
rect 60783 42721 60795 42755
rect 60737 42715 60795 42721
rect 66441 42755 66499 42761
rect 66441 42721 66453 42755
rect 66487 42752 66499 42755
rect 66990 42752 66996 42764
rect 66487 42724 66996 42752
rect 66487 42721 66499 42724
rect 66441 42715 66499 42721
rect 66990 42712 66996 42724
rect 67048 42712 67054 42764
rect 68738 42752 68744 42764
rect 68699 42724 68744 42752
rect 68738 42712 68744 42724
rect 68796 42752 68802 42764
rect 68925 42755 68983 42761
rect 68925 42752 68937 42755
rect 68796 42724 68937 42752
rect 68796 42712 68802 42724
rect 68925 42721 68937 42724
rect 68971 42721 68983 42755
rect 68925 42715 68983 42721
rect 69308 42693 69336 42792
rect 71590 42780 71596 42792
rect 71648 42820 71654 42832
rect 71648 42792 72188 42820
rect 71648 42780 71654 42792
rect 69661 42755 69719 42761
rect 69661 42721 69673 42755
rect 69707 42752 69719 42755
rect 71222 42752 71228 42764
rect 69707 42724 71228 42752
rect 69707 42721 69719 42724
rect 69661 42715 69719 42721
rect 71222 42712 71228 42724
rect 71280 42712 71286 42764
rect 72050 42752 72056 42764
rect 72011 42724 72056 42752
rect 72050 42712 72056 42724
rect 72108 42712 72114 42764
rect 72160 42752 72188 42792
rect 77478 42780 77484 42832
rect 77536 42820 77542 42832
rect 78582 42820 78588 42832
rect 77536 42792 78588 42820
rect 77536 42780 77542 42792
rect 72418 42752 72424 42764
rect 72160 42724 72424 42752
rect 72418 42712 72424 42724
rect 72476 42712 72482 42764
rect 72510 42712 72516 42764
rect 72568 42752 72574 42764
rect 78324 42761 78352 42792
rect 78582 42780 78588 42792
rect 78640 42780 78646 42832
rect 77757 42755 77815 42761
rect 77757 42752 77769 42755
rect 72568 42724 72613 42752
rect 77404 42724 77769 42752
rect 72568 42712 72574 42724
rect 69293 42687 69351 42693
rect 69293 42653 69305 42687
rect 69339 42653 69351 42687
rect 69293 42647 69351 42653
rect 71406 42644 71412 42696
rect 71464 42684 71470 42696
rect 71961 42687 72019 42693
rect 71961 42684 71973 42687
rect 71464 42656 71973 42684
rect 71464 42644 71470 42656
rect 71961 42653 71973 42656
rect 72007 42684 72019 42687
rect 72697 42687 72755 42693
rect 72697 42684 72709 42687
rect 72007 42656 72709 42684
rect 72007 42653 72019 42656
rect 71961 42647 72019 42653
rect 72697 42653 72709 42656
rect 72743 42684 72755 42687
rect 73338 42684 73344 42696
rect 72743 42656 73344 42684
rect 72743 42653 72755 42656
rect 72697 42647 72755 42653
rect 73338 42644 73344 42656
rect 73396 42644 73402 42696
rect 73614 42644 73620 42696
rect 73672 42684 73678 42696
rect 77404 42693 77432 42724
rect 77389 42687 77447 42693
rect 77389 42684 77401 42687
rect 73672 42656 77401 42684
rect 73672 42644 73678 42656
rect 77389 42653 77401 42656
rect 77435 42653 77447 42687
rect 77389 42647 77447 42653
rect 66165 42619 66223 42625
rect 66165 42585 66177 42619
rect 66211 42616 66223 42619
rect 66211 42588 66852 42616
rect 66211 42585 66223 42588
rect 66165 42579 66223 42585
rect 66824 42560 66852 42588
rect 67450 42576 67456 42628
rect 67508 42616 67514 42628
rect 69063 42619 69121 42625
rect 69063 42616 69075 42619
rect 67508 42588 69075 42616
rect 67508 42576 67514 42588
rect 69063 42585 69075 42588
rect 69109 42585 69121 42619
rect 69063 42579 69121 42585
rect 71501 42619 71559 42625
rect 71501 42585 71513 42619
rect 71547 42616 71559 42619
rect 72786 42616 72792 42628
rect 71547 42588 72792 42616
rect 71547 42585 71559 42588
rect 71501 42579 71559 42585
rect 72786 42576 72792 42588
rect 72844 42576 72850 42628
rect 60734 42548 60740 42560
rect 59096 42520 60740 42548
rect 58989 42511 59047 42517
rect 60734 42508 60740 42520
rect 60792 42508 60798 42560
rect 66622 42548 66628 42560
rect 66583 42520 66628 42548
rect 66622 42508 66628 42520
rect 66680 42508 66686 42560
rect 66806 42508 66812 42560
rect 66864 42548 66870 42560
rect 66993 42551 67051 42557
rect 66993 42548 67005 42551
rect 66864 42520 67005 42548
rect 66864 42508 66870 42520
rect 66993 42517 67005 42520
rect 67039 42517 67051 42551
rect 69198 42548 69204 42560
rect 69159 42520 69204 42548
rect 66993 42511 67051 42517
rect 69198 42508 69204 42520
rect 69256 42508 69262 42560
rect 77478 42508 77484 42560
rect 77536 42548 77542 42560
rect 77573 42551 77631 42557
rect 77573 42548 77585 42551
rect 77536 42520 77585 42548
rect 77536 42508 77542 42520
rect 77573 42517 77585 42520
rect 77619 42517 77631 42551
rect 77680 42548 77708 42724
rect 77757 42721 77769 42724
rect 77803 42721 77815 42755
rect 77757 42715 77815 42721
rect 78309 42755 78367 42761
rect 78309 42721 78321 42755
rect 78355 42721 78367 42755
rect 79686 42752 79692 42764
rect 79647 42724 79692 42752
rect 78309 42715 78367 42721
rect 79686 42712 79692 42724
rect 79744 42712 79750 42764
rect 78398 42684 78404 42696
rect 77772 42656 78404 42684
rect 77772 42628 77800 42656
rect 78398 42644 78404 42656
rect 78456 42684 78462 42696
rect 78585 42687 78643 42693
rect 78585 42684 78597 42687
rect 78456 42656 78597 42684
rect 78456 42644 78462 42656
rect 78585 42653 78597 42656
rect 78631 42653 78643 42687
rect 82170 42684 82176 42696
rect 78585 42647 78643 42653
rect 78692 42656 82176 42684
rect 77754 42576 77760 42628
rect 77812 42576 77818 42628
rect 78692 42548 78720 42656
rect 82170 42644 82176 42656
rect 82228 42644 82234 42696
rect 79778 42548 79784 42560
rect 77680 42520 78720 42548
rect 79739 42520 79784 42548
rect 77573 42511 77631 42517
rect 79778 42508 79784 42520
rect 79836 42508 79842 42560
rect 1104 42458 108008 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 65686 42458
rect 65738 42406 65750 42458
rect 65802 42406 65814 42458
rect 65866 42406 65878 42458
rect 65930 42406 96406 42458
rect 96458 42406 96470 42458
rect 96522 42406 96534 42458
rect 96586 42406 96598 42458
rect 96650 42406 108008 42458
rect 1104 42384 108008 42406
rect 3970 42344 3976 42356
rect 3931 42316 3976 42344
rect 3970 42304 3976 42316
rect 4028 42304 4034 42356
rect 4614 42344 4620 42356
rect 4575 42316 4620 42344
rect 4614 42304 4620 42316
rect 4672 42304 4678 42356
rect 7098 42304 7104 42356
rect 7156 42344 7162 42356
rect 7653 42347 7711 42353
rect 7653 42344 7665 42347
rect 7156 42316 7665 42344
rect 7156 42304 7162 42316
rect 7653 42313 7665 42316
rect 7699 42313 7711 42347
rect 7653 42307 7711 42313
rect 16209 42347 16267 42353
rect 16209 42313 16221 42347
rect 16255 42344 16267 42347
rect 16666 42344 16672 42356
rect 16255 42316 16672 42344
rect 16255 42313 16267 42316
rect 16209 42307 16267 42313
rect 16666 42304 16672 42316
rect 16724 42344 16730 42356
rect 17862 42344 17868 42356
rect 16724 42316 17868 42344
rect 16724 42304 16730 42316
rect 17862 42304 17868 42316
rect 17920 42304 17926 42356
rect 19613 42347 19671 42353
rect 19613 42313 19625 42347
rect 19659 42344 19671 42347
rect 20806 42344 20812 42356
rect 19659 42316 20812 42344
rect 19659 42313 19671 42316
rect 19613 42307 19671 42313
rect 2590 42208 2596 42220
rect 2503 42180 2596 42208
rect 2590 42168 2596 42180
rect 2648 42208 2654 42220
rect 4632 42208 4660 42304
rect 13722 42236 13728 42288
rect 13780 42276 13786 42288
rect 15933 42279 15991 42285
rect 15933 42276 15945 42279
rect 13780 42248 15945 42276
rect 13780 42236 13786 42248
rect 15933 42245 15945 42248
rect 15979 42276 15991 42279
rect 15979 42248 18920 42276
rect 15979 42245 15991 42248
rect 15933 42239 15991 42245
rect 2648 42180 4660 42208
rect 2648 42168 2654 42180
rect 2869 42143 2927 42149
rect 2869 42109 2881 42143
rect 2915 42140 2927 42143
rect 4341 42143 4399 42149
rect 4341 42140 4353 42143
rect 2915 42112 4353 42140
rect 2915 42109 2927 42112
rect 2869 42103 2927 42109
rect 4341 42109 4353 42112
rect 4387 42140 4399 42143
rect 4798 42140 4804 42152
rect 4387 42112 4804 42140
rect 4387 42109 4399 42112
rect 4341 42103 4399 42109
rect 4798 42100 4804 42112
rect 4856 42100 4862 42152
rect 7282 42100 7288 42152
rect 7340 42140 7346 42152
rect 7469 42143 7527 42149
rect 7469 42140 7481 42143
rect 7340 42112 7481 42140
rect 7340 42100 7346 42112
rect 7469 42109 7481 42112
rect 7515 42109 7527 42143
rect 7469 42103 7527 42109
rect 15749 42143 15807 42149
rect 15749 42109 15761 42143
rect 15795 42140 15807 42143
rect 16666 42140 16672 42152
rect 15795 42112 16672 42140
rect 15795 42109 15807 42112
rect 15749 42103 15807 42109
rect 16666 42100 16672 42112
rect 16724 42100 16730 42152
rect 18892 42149 18920 42248
rect 18969 42211 19027 42217
rect 18969 42177 18981 42211
rect 19015 42208 19027 42211
rect 19015 42180 19380 42208
rect 19015 42177 19027 42180
rect 18969 42171 19027 42177
rect 18877 42143 18935 42149
rect 18877 42109 18889 42143
rect 18923 42140 18935 42143
rect 19150 42140 19156 42152
rect 18923 42112 19156 42140
rect 18923 42109 18935 42112
rect 18877 42103 18935 42109
rect 19150 42100 19156 42112
rect 19208 42100 19214 42152
rect 19245 42143 19303 42149
rect 19245 42109 19257 42143
rect 19291 42109 19303 42143
rect 19245 42103 19303 42109
rect 17402 42032 17408 42084
rect 17460 42072 17466 42084
rect 18233 42075 18291 42081
rect 18233 42072 18245 42075
rect 17460 42044 18245 42072
rect 17460 42032 17466 42044
rect 18233 42041 18245 42044
rect 18279 42041 18291 42075
rect 18233 42035 18291 42041
rect 16206 41964 16212 42016
rect 16264 42004 16270 42016
rect 19260 42004 19288 42103
rect 19352 42072 19380 42180
rect 19429 42143 19487 42149
rect 19429 42109 19441 42143
rect 19475 42140 19487 42143
rect 19628 42140 19656 42307
rect 20806 42304 20812 42316
rect 20864 42304 20870 42356
rect 25409 42347 25467 42353
rect 25409 42313 25421 42347
rect 25455 42344 25467 42347
rect 26234 42344 26240 42356
rect 25455 42316 26240 42344
rect 25455 42313 25467 42316
rect 25409 42307 25467 42313
rect 26234 42304 26240 42316
rect 26292 42304 26298 42356
rect 27249 42347 27307 42353
rect 27249 42313 27261 42347
rect 27295 42344 27307 42347
rect 27522 42344 27528 42356
rect 27295 42316 27528 42344
rect 27295 42313 27307 42316
rect 27249 42307 27307 42313
rect 19797 42279 19855 42285
rect 19797 42245 19809 42279
rect 19843 42276 19855 42279
rect 19886 42276 19892 42288
rect 19843 42248 19892 42276
rect 19843 42245 19855 42248
rect 19797 42239 19855 42245
rect 19475 42112 19656 42140
rect 19475 42109 19487 42112
rect 19429 42103 19487 42109
rect 19812 42072 19840 42239
rect 19886 42236 19892 42248
rect 19944 42236 19950 42288
rect 20254 42168 20260 42220
rect 20312 42208 20318 42220
rect 20312 42180 20760 42208
rect 20312 42168 20318 42180
rect 20732 42140 20760 42180
rect 23952 42180 24440 42208
rect 23952 42140 23980 42180
rect 24412 42149 24440 42180
rect 24213 42143 24271 42149
rect 24213 42140 24225 42143
rect 20732 42112 23980 42140
rect 24044 42112 24225 42140
rect 19352 42044 19840 42072
rect 19334 42004 19340 42016
rect 16264 41976 19340 42004
rect 16264 41964 16270 41976
rect 19334 41964 19340 41976
rect 19392 41964 19398 42016
rect 23750 41964 23756 42016
rect 23808 42004 23814 42016
rect 24044 42013 24072 42112
rect 24213 42109 24225 42112
rect 24259 42109 24271 42143
rect 24213 42103 24271 42109
rect 24397 42143 24455 42149
rect 24397 42109 24409 42143
rect 24443 42140 24455 42143
rect 24949 42143 25007 42149
rect 24949 42140 24961 42143
rect 24443 42112 24961 42140
rect 24443 42109 24455 42112
rect 24397 42103 24455 42109
rect 24949 42109 24961 42112
rect 24995 42109 25007 42143
rect 25130 42140 25136 42152
rect 25091 42112 25136 42140
rect 24949 42103 25007 42109
rect 24964 42072 24992 42103
rect 25130 42100 25136 42112
rect 25188 42100 25194 42152
rect 26881 42143 26939 42149
rect 26881 42109 26893 42143
rect 26927 42140 26939 42143
rect 27264 42140 27292 42307
rect 27522 42304 27528 42316
rect 27580 42344 27586 42356
rect 51353 42347 51411 42353
rect 51353 42344 51365 42347
rect 27580 42316 51365 42344
rect 27580 42304 27586 42316
rect 51353 42313 51365 42316
rect 51399 42344 51411 42347
rect 51537 42347 51595 42353
rect 51537 42344 51549 42347
rect 51399 42316 51549 42344
rect 51399 42313 51411 42316
rect 51353 42307 51411 42313
rect 51537 42313 51549 42316
rect 51583 42313 51595 42347
rect 51537 42307 51595 42313
rect 53006 42304 53012 42356
rect 53064 42344 53070 42356
rect 53193 42347 53251 42353
rect 53193 42344 53205 42347
rect 53064 42316 53205 42344
rect 53064 42304 53070 42316
rect 53193 42313 53205 42316
rect 53239 42344 53251 42347
rect 53466 42344 53472 42356
rect 53239 42316 53472 42344
rect 53239 42313 53251 42316
rect 53193 42307 53251 42313
rect 53466 42304 53472 42316
rect 53524 42304 53530 42356
rect 58894 42304 58900 42356
rect 58952 42344 58958 42356
rect 60921 42347 60979 42353
rect 60921 42344 60933 42347
rect 58952 42316 60933 42344
rect 58952 42304 58958 42316
rect 60921 42313 60933 42316
rect 60967 42313 60979 42347
rect 64322 42344 64328 42356
rect 64283 42316 64328 42344
rect 60921 42307 60979 42313
rect 64322 42304 64328 42316
rect 64380 42304 64386 42356
rect 66990 42344 66996 42356
rect 66951 42316 66996 42344
rect 66990 42304 66996 42316
rect 67048 42304 67054 42356
rect 70486 42304 70492 42356
rect 70544 42344 70550 42356
rect 70765 42347 70823 42353
rect 70765 42344 70777 42347
rect 70544 42316 70777 42344
rect 70544 42304 70550 42316
rect 70765 42313 70777 42316
rect 70811 42344 70823 42347
rect 72050 42344 72056 42356
rect 70811 42316 72056 42344
rect 70811 42313 70823 42316
rect 70765 42307 70823 42313
rect 72050 42304 72056 42316
rect 72108 42304 72114 42356
rect 77846 42304 77852 42356
rect 77904 42344 77910 42356
rect 78033 42347 78091 42353
rect 78033 42344 78045 42347
rect 77904 42316 78045 42344
rect 77904 42304 77910 42316
rect 78033 42313 78045 42316
rect 78079 42313 78091 42347
rect 78033 42307 78091 42313
rect 29178 42236 29184 42288
rect 29236 42276 29242 42288
rect 31202 42276 31208 42288
rect 29236 42248 31208 42276
rect 29236 42236 29242 42248
rect 31202 42236 31208 42248
rect 31260 42236 31266 42288
rect 31297 42279 31355 42285
rect 31297 42245 31309 42279
rect 31343 42276 31355 42279
rect 32030 42276 32036 42288
rect 31343 42248 32036 42276
rect 31343 42245 31355 42248
rect 31297 42239 31355 42245
rect 32030 42236 32036 42248
rect 32088 42236 32094 42288
rect 32122 42236 32128 42288
rect 32180 42276 32186 42288
rect 58158 42276 58164 42288
rect 32180 42248 58164 42276
rect 32180 42236 32186 42248
rect 58158 42236 58164 42248
rect 58216 42236 58222 42288
rect 59262 42236 59268 42288
rect 59320 42276 59326 42288
rect 60001 42279 60059 42285
rect 60001 42276 60013 42279
rect 59320 42248 60013 42276
rect 59320 42236 59326 42248
rect 60001 42245 60013 42248
rect 60047 42276 60059 42279
rect 61102 42276 61108 42288
rect 60047 42248 61108 42276
rect 60047 42245 60059 42248
rect 60001 42239 60059 42245
rect 61102 42236 61108 42248
rect 61160 42236 61166 42288
rect 27338 42168 27344 42220
rect 27396 42208 27402 42220
rect 28994 42208 29000 42220
rect 27396 42180 29000 42208
rect 27396 42168 27402 42180
rect 28994 42168 29000 42180
rect 29052 42168 29058 42220
rect 40126 42168 40132 42220
rect 40184 42208 40190 42220
rect 45557 42211 45615 42217
rect 45557 42208 45569 42211
rect 40184 42180 45569 42208
rect 40184 42168 40190 42180
rect 45557 42177 45569 42180
rect 45603 42208 45615 42211
rect 46109 42211 46167 42217
rect 46109 42208 46121 42211
rect 45603 42180 46121 42208
rect 45603 42177 45615 42180
rect 45557 42171 45615 42177
rect 46109 42177 46121 42180
rect 46155 42177 46167 42211
rect 46109 42171 46167 42177
rect 51537 42211 51595 42217
rect 51537 42177 51549 42211
rect 51583 42208 51595 42211
rect 51721 42211 51779 42217
rect 51721 42208 51733 42211
rect 51583 42180 51733 42208
rect 51583 42177 51595 42180
rect 51537 42171 51595 42177
rect 51721 42177 51733 42180
rect 51767 42177 51779 42211
rect 51721 42171 51779 42177
rect 53006 42168 53012 42220
rect 53064 42168 53070 42220
rect 58437 42211 58495 42217
rect 58437 42177 58449 42211
rect 58483 42208 58495 42211
rect 58802 42208 58808 42220
rect 58483 42180 58808 42208
rect 58483 42177 58495 42180
rect 58437 42171 58495 42177
rect 58802 42168 58808 42180
rect 58860 42168 58866 42220
rect 64340 42208 64368 42304
rect 64417 42211 64475 42217
rect 64417 42208 64429 42211
rect 64340 42180 64429 42208
rect 64417 42177 64429 42180
rect 64463 42177 64475 42211
rect 64417 42171 64475 42177
rect 64693 42211 64751 42217
rect 64693 42177 64705 42211
rect 64739 42208 64751 42211
rect 66622 42208 66628 42220
rect 64739 42180 66628 42208
rect 64739 42177 64751 42180
rect 64693 42171 64751 42177
rect 66622 42168 66628 42180
rect 66680 42168 66686 42220
rect 66714 42168 66720 42220
rect 66772 42208 66778 42220
rect 69109 42211 69167 42217
rect 69109 42208 69121 42211
rect 66772 42180 69121 42208
rect 66772 42168 66778 42180
rect 31113 42143 31171 42149
rect 31113 42140 31125 42143
rect 26927 42112 27292 42140
rect 30944 42112 31125 42140
rect 26927 42109 26939 42112
rect 26881 42103 26939 42109
rect 29638 42072 29644 42084
rect 24964 42044 29644 42072
rect 29638 42032 29644 42044
rect 29696 42032 29702 42084
rect 24029 42007 24087 42013
rect 24029 42004 24041 42007
rect 23808 41976 24041 42004
rect 23808 41964 23814 41976
rect 24029 41973 24041 41976
rect 24075 41973 24087 42007
rect 24029 41967 24087 41973
rect 26510 41964 26516 42016
rect 26568 42004 26574 42016
rect 26973 42007 27031 42013
rect 26973 42004 26985 42007
rect 26568 41976 26985 42004
rect 26568 41964 26574 41976
rect 26973 41973 26985 41976
rect 27019 41973 27031 42007
rect 26973 41967 27031 41973
rect 29270 41964 29276 42016
rect 29328 42004 29334 42016
rect 30944 42013 30972 42112
rect 31113 42109 31125 42112
rect 31159 42109 31171 42143
rect 31113 42103 31171 42109
rect 31202 42100 31208 42152
rect 31260 42140 31266 42152
rect 36262 42140 36268 42152
rect 31260 42112 36268 42140
rect 31260 42100 31266 42112
rect 36262 42100 36268 42112
rect 36320 42100 36326 42152
rect 46290 42100 46296 42152
rect 46348 42140 46354 42152
rect 46753 42143 46811 42149
rect 46348 42112 46393 42140
rect 46348 42100 46354 42112
rect 46753 42109 46765 42143
rect 46799 42109 46811 42143
rect 46753 42103 46811 42109
rect 46845 42143 46903 42149
rect 46845 42109 46857 42143
rect 46891 42109 46903 42143
rect 46845 42103 46903 42109
rect 51905 42143 51963 42149
rect 51905 42109 51917 42143
rect 51951 42140 51963 42143
rect 52270 42140 52276 42152
rect 51951 42112 52276 42140
rect 51951 42109 51963 42112
rect 51905 42103 51963 42109
rect 46768 42016 46796 42103
rect 30929 42007 30987 42013
rect 30929 42004 30941 42007
rect 29328 41976 30941 42004
rect 29328 41964 29334 41976
rect 30929 41973 30941 41976
rect 30975 41973 30987 42007
rect 30929 41967 30987 41973
rect 40034 41964 40040 42016
rect 40092 42004 40098 42016
rect 41230 42004 41236 42016
rect 40092 41976 41236 42004
rect 40092 41964 40098 41976
rect 41230 41964 41236 41976
rect 41288 41964 41294 42016
rect 45833 42007 45891 42013
rect 45833 41973 45845 42007
rect 45879 42004 45891 42007
rect 46750 42004 46756 42016
rect 45879 41976 46756 42004
rect 45879 41973 45891 41976
rect 45833 41967 45891 41973
rect 46750 41964 46756 41976
rect 46808 41964 46814 42016
rect 46860 42004 46888 42103
rect 52270 42100 52276 42112
rect 52328 42100 52334 42152
rect 52365 42143 52423 42149
rect 52365 42109 52377 42143
rect 52411 42109 52423 42143
rect 52365 42103 52423 42109
rect 52457 42143 52515 42149
rect 52457 42109 52469 42143
rect 52503 42140 52515 42143
rect 53024 42140 53052 42168
rect 52503 42112 53052 42140
rect 58161 42143 58219 42149
rect 52503 42109 52515 42112
rect 52457 42103 52515 42109
rect 58161 42109 58173 42143
rect 58207 42140 58219 42143
rect 59262 42140 59268 42152
rect 58207 42112 59268 42140
rect 58207 42109 58219 42112
rect 58161 42103 58219 42109
rect 47397 42075 47455 42081
rect 47397 42041 47409 42075
rect 47443 42072 47455 42075
rect 49510 42072 49516 42084
rect 47443 42044 49516 42072
rect 47443 42041 47455 42044
rect 47397 42035 47455 42041
rect 49510 42032 49516 42044
rect 49568 42032 49574 42084
rect 51442 42072 51448 42084
rect 51184 42044 51448 42072
rect 51184 42016 51212 42044
rect 51442 42032 51448 42044
rect 51500 42072 51506 42084
rect 52380 42072 52408 42103
rect 59262 42100 59268 42112
rect 59320 42100 59326 42152
rect 67192 42149 67220 42180
rect 69109 42177 69121 42180
rect 69155 42177 69167 42211
rect 69109 42171 69167 42177
rect 72421 42211 72479 42217
rect 72421 42177 72433 42211
rect 72467 42208 72479 42211
rect 72510 42208 72516 42220
rect 72467 42180 72516 42208
rect 72467 42177 72479 42180
rect 72421 42171 72479 42177
rect 72510 42168 72516 42180
rect 72568 42168 72574 42220
rect 77570 42208 77576 42220
rect 77483 42180 77576 42208
rect 77570 42168 77576 42180
rect 77628 42208 77634 42220
rect 78401 42211 78459 42217
rect 78401 42208 78413 42211
rect 77628 42180 78413 42208
rect 77628 42168 77634 42180
rect 78401 42177 78413 42180
rect 78447 42177 78459 42211
rect 78401 42171 78459 42177
rect 60829 42143 60887 42149
rect 60829 42109 60841 42143
rect 60875 42109 60887 42143
rect 60829 42103 60887 42109
rect 67177 42143 67235 42149
rect 67177 42109 67189 42143
rect 67223 42109 67235 42143
rect 67450 42140 67456 42152
rect 67411 42112 67456 42140
rect 67177 42103 67235 42109
rect 53006 42072 53012 42084
rect 51500 42044 52408 42072
rect 52967 42044 53012 42072
rect 51500 42032 51506 42044
rect 53006 42032 53012 42044
rect 53064 42032 53070 42084
rect 53116 42044 53328 42072
rect 47670 42004 47676 42016
rect 46860 41976 47676 42004
rect 47670 41964 47676 41976
rect 47728 41964 47734 42016
rect 51166 42004 51172 42016
rect 51127 41976 51172 42004
rect 51166 41964 51172 41976
rect 51224 41964 51230 42016
rect 51258 41964 51264 42016
rect 51316 42004 51322 42016
rect 53116 42004 53144 42044
rect 51316 41976 53144 42004
rect 53300 42004 53328 42044
rect 59630 42032 59636 42084
rect 59688 42072 59694 42084
rect 60645 42075 60703 42081
rect 60645 42072 60657 42075
rect 59688 42044 60657 42072
rect 59688 42032 59694 42044
rect 60645 42041 60657 42044
rect 60691 42041 60703 42075
rect 60645 42035 60703 42041
rect 58434 42004 58440 42016
rect 53300 41976 58440 42004
rect 51316 41964 51322 41976
rect 58434 41964 58440 41976
rect 58492 41964 58498 42016
rect 59722 42004 59728 42016
rect 59683 41976 59728 42004
rect 59722 41964 59728 41976
rect 59780 42004 59786 42016
rect 60844 42004 60872 42103
rect 67450 42100 67456 42112
rect 67508 42100 67514 42152
rect 68833 42143 68891 42149
rect 68833 42140 68845 42143
rect 68480 42112 68845 42140
rect 66070 42032 66076 42084
rect 66128 42072 66134 42084
rect 68480 42072 68508 42112
rect 68833 42109 68845 42112
rect 68879 42140 68891 42143
rect 69198 42140 69204 42152
rect 68879 42112 69204 42140
rect 68879 42109 68891 42112
rect 68833 42103 68891 42109
rect 69198 42100 69204 42112
rect 69256 42100 69262 42152
rect 70681 42143 70739 42149
rect 70681 42109 70693 42143
rect 70727 42109 70739 42143
rect 70681 42103 70739 42109
rect 66128 42044 68508 42072
rect 68649 42075 68707 42081
rect 66128 42032 66134 42044
rect 68649 42041 68661 42075
rect 68695 42072 68707 42075
rect 68695 42044 70440 42072
rect 68695 42041 68707 42044
rect 68649 42035 68707 42041
rect 65978 42004 65984 42016
rect 59780 41976 60872 42004
rect 65939 41976 65984 42004
rect 59780 41964 59786 41976
rect 65978 41964 65984 41976
rect 66036 41964 66042 42016
rect 66438 41964 66444 42016
rect 66496 42004 66502 42016
rect 66898 42004 66904 42016
rect 66496 41976 66904 42004
rect 66496 41964 66502 41976
rect 66898 41964 66904 41976
rect 66956 42004 66962 42016
rect 67450 42004 67456 42016
rect 66956 41976 67456 42004
rect 66956 41964 66962 41976
rect 67450 41964 67456 41976
rect 67508 41964 67514 42016
rect 70412 42004 70440 42044
rect 70688 42004 70716 42103
rect 71958 42100 71964 42152
rect 72016 42140 72022 42152
rect 72053 42143 72111 42149
rect 72053 42140 72065 42143
rect 72016 42112 72065 42140
rect 72016 42100 72022 42112
rect 72053 42109 72065 42112
rect 72099 42140 72111 42143
rect 72605 42143 72663 42149
rect 72605 42140 72617 42143
rect 72099 42112 72617 42140
rect 72099 42109 72111 42112
rect 72053 42103 72111 42109
rect 72605 42109 72617 42112
rect 72651 42109 72663 42143
rect 72605 42103 72663 42109
rect 77662 42100 77668 42152
rect 77720 42140 77726 42152
rect 77849 42143 77907 42149
rect 77849 42140 77861 42143
rect 77720 42112 77861 42140
rect 77720 42100 77726 42112
rect 77849 42109 77861 42112
rect 77895 42109 77907 42143
rect 77849 42103 77907 42109
rect 71866 42072 71872 42084
rect 71779 42044 71872 42072
rect 71866 42032 71872 42044
rect 71924 42072 71930 42084
rect 72694 42072 72700 42084
rect 71924 42044 72700 42072
rect 71924 42032 71930 42044
rect 72694 42032 72700 42044
rect 72752 42032 72758 42084
rect 77754 42072 77760 42084
rect 77715 42044 77760 42072
rect 77754 42032 77760 42044
rect 77812 42032 77818 42084
rect 71774 42004 71780 42016
rect 70412 41976 71780 42004
rect 71774 41964 71780 41976
rect 71832 41964 71838 42016
rect 1104 41914 108008 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 81046 41914
rect 81098 41862 81110 41914
rect 81162 41862 81174 41914
rect 81226 41862 81238 41914
rect 81290 41862 108008 41914
rect 1104 41840 108008 41862
rect 4614 41760 4620 41812
rect 4672 41800 4678 41812
rect 5997 41803 6055 41809
rect 5997 41800 6009 41803
rect 4672 41772 6009 41800
rect 4672 41760 4678 41772
rect 5997 41769 6009 41772
rect 6043 41769 6055 41803
rect 5997 41763 6055 41769
rect 12897 41803 12955 41809
rect 12897 41769 12909 41803
rect 12943 41800 12955 41803
rect 13446 41800 13452 41812
rect 12943 41772 13452 41800
rect 12943 41769 12955 41772
rect 12897 41763 12955 41769
rect 11146 41732 11152 41744
rect 7208 41704 11152 41732
rect 6181 41667 6239 41673
rect 6181 41633 6193 41667
rect 6227 41633 6239 41667
rect 6181 41627 6239 41633
rect 6457 41667 6515 41673
rect 6457 41633 6469 41667
rect 6503 41664 6515 41667
rect 7208 41664 7236 41704
rect 11146 41692 11152 41704
rect 11204 41692 11210 41744
rect 6503 41636 7236 41664
rect 6503 41633 6515 41636
rect 6457 41627 6515 41633
rect 6196 41596 6224 41627
rect 7282 41624 7288 41676
rect 7340 41664 7346 41676
rect 7469 41667 7527 41673
rect 7469 41664 7481 41667
rect 7340 41636 7481 41664
rect 7340 41624 7346 41636
rect 7469 41633 7481 41636
rect 7515 41633 7527 41667
rect 7469 41627 7527 41633
rect 11057 41667 11115 41673
rect 11057 41633 11069 41667
rect 11103 41664 11115 41667
rect 12912 41664 12940 41763
rect 13446 41760 13452 41772
rect 13504 41760 13510 41812
rect 13998 41760 14004 41812
rect 14056 41800 14062 41812
rect 16117 41803 16175 41809
rect 16117 41800 16129 41803
rect 14056 41772 16129 41800
rect 14056 41760 14062 41772
rect 16117 41769 16129 41772
rect 16163 41800 16175 41803
rect 16206 41800 16212 41812
rect 16163 41772 16212 41800
rect 16163 41769 16175 41772
rect 16117 41763 16175 41769
rect 16206 41760 16212 41772
rect 16264 41760 16270 41812
rect 16390 41800 16396 41812
rect 16351 41772 16396 41800
rect 16390 41760 16396 41772
rect 16448 41760 16454 41812
rect 19426 41760 19432 41812
rect 19484 41800 19490 41812
rect 25130 41800 25136 41812
rect 19484 41772 25136 41800
rect 19484 41760 19490 41772
rect 25130 41760 25136 41772
rect 25188 41760 25194 41812
rect 27249 41803 27307 41809
rect 27249 41769 27261 41803
rect 27295 41800 27307 41803
rect 27338 41800 27344 41812
rect 27295 41772 27344 41800
rect 27295 41769 27307 41772
rect 27249 41763 27307 41769
rect 11103 41636 12940 41664
rect 15933 41667 15991 41673
rect 11103 41633 11115 41636
rect 11057 41627 11115 41633
rect 15933 41633 15945 41667
rect 15979 41664 15991 41667
rect 16114 41664 16120 41676
rect 15979 41636 16120 41664
rect 15979 41633 15991 41636
rect 15933 41627 15991 41633
rect 16114 41624 16120 41636
rect 16172 41664 16178 41676
rect 16390 41664 16396 41676
rect 16172 41636 16396 41664
rect 16172 41624 16178 41636
rect 16390 41624 16396 41636
rect 16448 41624 16454 41676
rect 25148 41664 25176 41760
rect 26510 41664 26516 41676
rect 25148 41636 26516 41664
rect 26510 41624 26516 41636
rect 26568 41624 26574 41676
rect 26605 41667 26663 41673
rect 26605 41633 26617 41667
rect 26651 41664 26663 41667
rect 27264 41664 27292 41763
rect 27338 41760 27344 41772
rect 27396 41760 27402 41812
rect 29638 41800 29644 41812
rect 29599 41772 29644 41800
rect 29638 41760 29644 41772
rect 29696 41760 29702 41812
rect 29914 41800 29920 41812
rect 29875 41772 29920 41800
rect 29914 41760 29920 41772
rect 29972 41760 29978 41812
rect 34701 41803 34759 41809
rect 34701 41769 34713 41803
rect 34747 41800 34759 41803
rect 51258 41800 51264 41812
rect 34747 41772 51264 41800
rect 34747 41769 34759 41772
rect 34701 41763 34759 41769
rect 51258 41760 51264 41772
rect 51316 41760 51322 41812
rect 53466 41800 53472 41812
rect 53427 41772 53472 41800
rect 53466 41760 53472 41772
rect 53524 41760 53530 41812
rect 60277 41803 60335 41809
rect 60277 41769 60289 41803
rect 60323 41800 60335 41803
rect 60734 41800 60740 41812
rect 60323 41772 60740 41800
rect 60323 41769 60335 41772
rect 60277 41763 60335 41769
rect 60734 41760 60740 41772
rect 60792 41760 60798 41812
rect 79778 41800 79784 41812
rect 76208 41772 79784 41800
rect 27893 41667 27951 41673
rect 27893 41664 27905 41667
rect 26651 41636 27292 41664
rect 27632 41636 27905 41664
rect 26651 41633 26663 41636
rect 26605 41627 26663 41633
rect 6822 41596 6828 41608
rect 6196 41568 6828 41596
rect 6822 41556 6828 41568
rect 6880 41596 6886 41608
rect 11330 41596 11336 41608
rect 6880 41568 7696 41596
rect 11291 41568 11336 41596
rect 6880 41556 6886 41568
rect 7668 41537 7696 41568
rect 11330 41556 11336 41568
rect 11388 41556 11394 41608
rect 7653 41531 7711 41537
rect 7653 41497 7665 41531
rect 7699 41497 7711 41531
rect 27632 41528 27660 41636
rect 27893 41633 27905 41636
rect 27939 41633 27951 41667
rect 27893 41627 27951 41633
rect 29362 41624 29368 41676
rect 29420 41664 29426 41676
rect 29457 41667 29515 41673
rect 29457 41664 29469 41667
rect 29420 41636 29469 41664
rect 29420 41624 29426 41636
rect 29457 41633 29469 41636
rect 29503 41664 29515 41667
rect 29932 41664 29960 41760
rect 34977 41735 35035 41741
rect 34977 41701 34989 41735
rect 35023 41732 35035 41735
rect 35434 41732 35440 41744
rect 35023 41704 35440 41732
rect 35023 41701 35035 41704
rect 34977 41695 35035 41701
rect 29503 41636 29960 41664
rect 29503 41633 29515 41636
rect 29457 41627 29515 41633
rect 31754 41624 31760 41676
rect 31812 41664 31818 41676
rect 33413 41667 33471 41673
rect 33413 41664 33425 41667
rect 31812 41636 33425 41664
rect 31812 41624 31818 41636
rect 33413 41633 33425 41636
rect 33459 41633 33471 41667
rect 33413 41627 33471 41633
rect 33137 41599 33195 41605
rect 33137 41565 33149 41599
rect 33183 41596 33195 41599
rect 34992 41596 35020 41695
rect 35434 41692 35440 41704
rect 35492 41692 35498 41744
rect 38562 41692 38568 41744
rect 38620 41732 38626 41744
rect 39117 41735 39175 41741
rect 39117 41732 39129 41735
rect 38620 41704 39129 41732
rect 38620 41692 38626 41704
rect 39117 41701 39129 41704
rect 39163 41732 39175 41735
rect 39163 41704 40264 41732
rect 39163 41701 39175 41704
rect 39117 41695 39175 41701
rect 39390 41624 39396 41676
rect 39448 41664 39454 41676
rect 39485 41667 39543 41673
rect 39485 41664 39497 41667
rect 39448 41636 39497 41664
rect 39448 41624 39454 41636
rect 39485 41633 39497 41636
rect 39531 41633 39543 41667
rect 40034 41664 40040 41676
rect 39995 41636 40040 41664
rect 39485 41627 39543 41633
rect 40034 41624 40040 41636
rect 40092 41624 40098 41676
rect 40236 41673 40264 41704
rect 46584 41704 47440 41732
rect 40221 41667 40279 41673
rect 40221 41633 40233 41667
rect 40267 41664 40279 41667
rect 45649 41667 45707 41673
rect 45649 41664 45661 41667
rect 40267 41636 45661 41664
rect 40267 41633 40279 41636
rect 40221 41627 40279 41633
rect 45649 41633 45661 41636
rect 45695 41664 45707 41667
rect 45833 41667 45891 41673
rect 45833 41664 45845 41667
rect 45695 41636 45845 41664
rect 45695 41633 45707 41636
rect 45649 41627 45707 41633
rect 45833 41633 45845 41636
rect 45879 41633 45891 41667
rect 45833 41627 45891 41633
rect 46017 41667 46075 41673
rect 46017 41633 46029 41667
rect 46063 41664 46075 41667
rect 46106 41664 46112 41676
rect 46063 41636 46112 41664
rect 46063 41633 46075 41636
rect 46017 41627 46075 41633
rect 33183 41568 35020 41596
rect 33183 41565 33195 41568
rect 33137 41559 33195 41565
rect 35066 41556 35072 41608
rect 35124 41596 35130 41608
rect 39298 41596 39304 41608
rect 35124 41568 38516 41596
rect 39259 41568 39304 41596
rect 35124 41556 35130 41568
rect 27706 41528 27712 41540
rect 27619 41500 27712 41528
rect 7653 41491 7711 41497
rect 27706 41488 27712 41500
rect 27764 41528 27770 41540
rect 27801 41531 27859 41537
rect 27801 41528 27813 41531
rect 27764 41500 27813 41528
rect 27764 41488 27770 41500
rect 27801 41497 27813 41500
rect 27847 41528 27859 41531
rect 30742 41528 30748 41540
rect 27847 41500 30748 41528
rect 27847 41497 27859 41500
rect 27801 41491 27859 41497
rect 30742 41488 30748 41500
rect 30800 41488 30806 41540
rect 38488 41528 38516 41568
rect 39298 41556 39304 41568
rect 39356 41556 39362 41608
rect 41230 41556 41236 41608
rect 41288 41596 41294 41608
rect 46032 41596 46060 41627
rect 46106 41624 46112 41636
rect 46164 41624 46170 41676
rect 46584 41673 46612 41704
rect 47412 41676 47440 41704
rect 47670 41692 47676 41744
rect 47728 41732 47734 41744
rect 66625 41735 66683 41741
rect 47728 41704 65656 41732
rect 47728 41692 47734 41704
rect 46569 41667 46627 41673
rect 46569 41633 46581 41667
rect 46615 41633 46627 41667
rect 46569 41627 46627 41633
rect 46750 41624 46756 41676
rect 46808 41664 46814 41676
rect 47394 41664 47400 41676
rect 46808 41636 46853 41664
rect 47307 41636 47400 41664
rect 46808 41624 46814 41636
rect 47394 41624 47400 41636
rect 47452 41664 47458 41676
rect 48774 41664 48780 41676
rect 47452 41636 48780 41664
rect 47452 41624 47458 41636
rect 48774 41624 48780 41636
rect 48832 41664 48838 41676
rect 52181 41667 52239 41673
rect 48832 41636 52132 41664
rect 48832 41624 48838 41636
rect 41288 41568 46060 41596
rect 47121 41599 47179 41605
rect 41288 41556 41294 41568
rect 47121 41565 47133 41599
rect 47167 41596 47179 41599
rect 49602 41596 49608 41608
rect 47167 41568 49608 41596
rect 47167 41565 47179 41568
rect 47121 41559 47179 41565
rect 49602 41556 49608 41568
rect 49660 41556 49666 41608
rect 51997 41599 52055 41605
rect 51997 41565 52009 41599
rect 52043 41565 52055 41599
rect 51997 41559 52055 41565
rect 38562 41528 38568 41540
rect 38488 41500 38568 41528
rect 38562 41488 38568 41500
rect 38620 41488 38626 41540
rect 38746 41488 38752 41540
rect 38804 41528 38810 41540
rect 51629 41531 51687 41537
rect 51629 41528 51641 41531
rect 38804 41500 51641 41528
rect 38804 41488 38810 41500
rect 51629 41497 51641 41500
rect 51675 41528 51687 41531
rect 52012 41528 52040 41559
rect 51675 41500 52040 41528
rect 52104 41528 52132 41636
rect 52181 41633 52193 41667
rect 52227 41664 52239 41667
rect 52270 41664 52276 41676
rect 52227 41636 52276 41664
rect 52227 41633 52239 41636
rect 52181 41627 52239 41633
rect 52270 41624 52276 41636
rect 52328 41624 52334 41676
rect 52546 41624 52552 41676
rect 52604 41664 52610 41676
rect 52641 41667 52699 41673
rect 52641 41664 52653 41667
rect 52604 41636 52653 41664
rect 52604 41624 52610 41636
rect 52641 41633 52653 41636
rect 52687 41633 52699 41667
rect 52641 41627 52699 41633
rect 52733 41667 52791 41673
rect 52733 41633 52745 41667
rect 52779 41664 52791 41667
rect 53374 41664 53380 41676
rect 52779 41636 53380 41664
rect 52779 41633 52791 41636
rect 52733 41627 52791 41633
rect 53374 41624 53380 41636
rect 53432 41624 53438 41676
rect 58158 41624 58164 41676
rect 58216 41664 58222 41676
rect 60185 41667 60243 41673
rect 60185 41664 60197 41667
rect 58216 41636 60197 41664
rect 58216 41624 58222 41636
rect 60185 41633 60197 41636
rect 60231 41664 60243 41667
rect 60461 41667 60519 41673
rect 60461 41664 60473 41667
rect 60231 41636 60473 41664
rect 60231 41633 60243 41636
rect 60185 41627 60243 41633
rect 60461 41633 60473 41636
rect 60507 41664 60519 41667
rect 60826 41664 60832 41676
rect 60507 41636 60832 41664
rect 60507 41633 60519 41636
rect 60461 41627 60519 41633
rect 60826 41624 60832 41636
rect 60884 41624 60890 41676
rect 53285 41599 53343 41605
rect 53285 41565 53297 41599
rect 53331 41596 53343 41599
rect 53466 41596 53472 41608
rect 53331 41568 53472 41596
rect 53331 41565 53343 41568
rect 53285 41559 53343 41565
rect 53466 41556 53472 41568
rect 53524 41556 53530 41608
rect 65628 41596 65656 41704
rect 66625 41701 66637 41735
rect 66671 41732 66683 41735
rect 70486 41732 70492 41744
rect 66671 41704 70492 41732
rect 66671 41701 66683 41704
rect 66625 41695 66683 41701
rect 70486 41692 70492 41704
rect 70544 41692 70550 41744
rect 66806 41664 66812 41676
rect 66767 41636 66812 41664
rect 66806 41624 66812 41636
rect 66864 41624 66870 41676
rect 71866 41664 71872 41676
rect 66916 41636 71872 41664
rect 66916 41596 66944 41636
rect 71866 41624 71872 41636
rect 71924 41624 71930 41676
rect 72142 41624 72148 41676
rect 72200 41664 72206 41676
rect 72329 41667 72387 41673
rect 72329 41664 72341 41667
rect 72200 41636 72341 41664
rect 72200 41624 72206 41636
rect 72329 41633 72341 41636
rect 72375 41633 72387 41667
rect 72329 41627 72387 41633
rect 72418 41624 72424 41676
rect 72476 41664 72482 41676
rect 72513 41667 72571 41673
rect 72513 41664 72525 41667
rect 72476 41636 72525 41664
rect 72476 41624 72482 41636
rect 72513 41633 72525 41636
rect 72559 41664 72571 41667
rect 74258 41664 74264 41676
rect 72559 41636 74264 41664
rect 72559 41633 72571 41636
rect 72513 41627 72571 41633
rect 74258 41624 74264 41636
rect 74316 41624 74322 41676
rect 75825 41667 75883 41673
rect 75825 41633 75837 41667
rect 75871 41633 75883 41667
rect 75825 41627 75883 41633
rect 65628 41568 66944 41596
rect 71884 41596 71912 41624
rect 72786 41596 72792 41608
rect 71884 41568 72792 41596
rect 72786 41556 72792 41568
rect 72844 41596 72850 41608
rect 75840 41596 75868 41627
rect 76208 41605 76236 41772
rect 79778 41760 79784 41772
rect 79836 41760 79842 41812
rect 77386 41732 77392 41744
rect 77347 41704 77392 41732
rect 77386 41692 77392 41704
rect 77444 41692 77450 41744
rect 77110 41624 77116 41676
rect 77168 41664 77174 41676
rect 77404 41664 77432 41692
rect 77573 41667 77631 41673
rect 77573 41664 77585 41667
rect 77168 41636 77585 41664
rect 77168 41624 77174 41636
rect 77573 41633 77585 41636
rect 77619 41633 77631 41667
rect 77846 41664 77852 41676
rect 77807 41636 77852 41664
rect 77573 41627 77631 41633
rect 76193 41599 76251 41605
rect 76193 41596 76205 41599
rect 72844 41568 76205 41596
rect 72844 41556 72850 41568
rect 76193 41565 76205 41568
rect 76239 41565 76251 41599
rect 77588 41596 77616 41627
rect 77846 41624 77852 41636
rect 77904 41624 77910 41676
rect 83185 41599 83243 41605
rect 83185 41596 83197 41599
rect 77588 41568 83197 41596
rect 76193 41559 76251 41565
rect 83185 41565 83197 41568
rect 83231 41596 83243 41599
rect 83366 41596 83372 41608
rect 83231 41568 83372 41596
rect 83231 41565 83243 41568
rect 83185 41559 83243 41565
rect 83366 41556 83372 41568
rect 83424 41556 83430 41608
rect 83642 41596 83648 41608
rect 83603 41568 83648 41596
rect 83642 41556 83648 41568
rect 83700 41556 83706 41608
rect 76009 41531 76067 41537
rect 76009 41528 76021 41531
rect 52104 41500 76021 41528
rect 51675 41497 51687 41500
rect 51629 41491 51687 41497
rect 76009 41497 76021 41500
rect 76055 41528 76067 41531
rect 77478 41528 77484 41540
rect 76055 41500 77484 41528
rect 76055 41497 76067 41500
rect 76009 41491 76067 41497
rect 77478 41488 77484 41500
rect 77536 41488 77542 41540
rect 12437 41463 12495 41469
rect 12437 41429 12449 41463
rect 12483 41460 12495 41463
rect 12526 41460 12532 41472
rect 12483 41432 12532 41460
rect 12483 41429 12495 41432
rect 12437 41423 12495 41429
rect 12526 41420 12532 41432
rect 12584 41420 12590 41472
rect 26602 41420 26608 41472
rect 26660 41460 26666 41472
rect 26789 41463 26847 41469
rect 26789 41460 26801 41463
rect 26660 41432 26801 41460
rect 26660 41420 26666 41432
rect 26789 41429 26801 41432
rect 26835 41429 26847 41463
rect 27982 41460 27988 41472
rect 27943 41432 27988 41460
rect 26789 41423 26847 41429
rect 27982 41420 27988 41432
rect 28040 41420 28046 41472
rect 40494 41460 40500 41472
rect 40455 41432 40500 41460
rect 40494 41420 40500 41432
rect 40552 41420 40558 41472
rect 40865 41463 40923 41469
rect 40865 41429 40877 41463
rect 40911 41460 40923 41463
rect 41598 41460 41604 41472
rect 40911 41432 41604 41460
rect 40911 41429 40923 41432
rect 40865 41423 40923 41429
rect 41598 41420 41604 41432
rect 41656 41420 41662 41472
rect 45462 41460 45468 41472
rect 45423 41432 45468 41460
rect 45462 41420 45468 41432
rect 45520 41420 45526 41472
rect 51810 41460 51816 41472
rect 51771 41432 51816 41460
rect 51810 41420 51816 41432
rect 51868 41460 51874 41472
rect 52546 41460 52552 41472
rect 51868 41432 52552 41460
rect 51868 41420 51874 41432
rect 52546 41420 52552 41432
rect 52604 41420 52610 41472
rect 66622 41420 66628 41472
rect 66680 41460 66686 41472
rect 66901 41463 66959 41469
rect 66901 41460 66913 41463
rect 66680 41432 66913 41460
rect 66680 41420 66686 41432
rect 66901 41429 66913 41432
rect 66947 41429 66959 41463
rect 72602 41460 72608 41472
rect 72563 41432 72608 41460
rect 66901 41423 66959 41429
rect 72602 41420 72608 41432
rect 72660 41420 72666 41472
rect 78950 41460 78956 41472
rect 78911 41432 78956 41460
rect 78950 41420 78956 41432
rect 79008 41420 79014 41472
rect 84562 41420 84568 41472
rect 84620 41460 84626 41472
rect 84749 41463 84807 41469
rect 84749 41460 84761 41463
rect 84620 41432 84761 41460
rect 84620 41420 84626 41432
rect 84749 41429 84761 41432
rect 84795 41429 84807 41463
rect 84749 41423 84807 41429
rect 1104 41370 108008 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 65686 41370
rect 65738 41318 65750 41370
rect 65802 41318 65814 41370
rect 65866 41318 65878 41370
rect 65930 41318 96406 41370
rect 96458 41318 96470 41370
rect 96522 41318 96534 41370
rect 96586 41318 96598 41370
rect 96650 41318 108008 41370
rect 1104 41296 108008 41318
rect 4062 41216 4068 41268
rect 4120 41256 4126 41268
rect 7006 41256 7012 41268
rect 4120 41228 7012 41256
rect 4120 41216 4126 41228
rect 7006 41216 7012 41228
rect 7064 41216 7070 41268
rect 11054 41256 11060 41268
rect 7392 41228 11060 41256
rect 4433 41191 4491 41197
rect 4433 41157 4445 41191
rect 4479 41188 4491 41191
rect 4706 41188 4712 41200
rect 4479 41160 4712 41188
rect 4479 41157 4491 41160
rect 4433 41151 4491 41157
rect 4706 41148 4712 41160
rect 4764 41148 4770 41200
rect 3970 41120 3976 41132
rect 3931 41092 3976 41120
rect 3970 41080 3976 41092
rect 4028 41080 4034 41132
rect 2590 41012 2596 41064
rect 2648 41061 2654 41064
rect 2648 41052 2658 41061
rect 2869 41055 2927 41061
rect 2648 41024 2693 41052
rect 2648 41015 2658 41024
rect 2869 41021 2881 41055
rect 2915 41052 2927 41055
rect 4614 41052 4620 41064
rect 2915 41024 4620 41052
rect 2915 41021 2927 41024
rect 2869 41015 2927 41021
rect 2648 41012 2654 41015
rect 4614 41012 4620 41024
rect 4672 41012 4678 41064
rect 5445 41055 5503 41061
rect 5445 41021 5457 41055
rect 5491 41052 5503 41055
rect 5534 41052 5540 41064
rect 5491 41024 5540 41052
rect 5491 41021 5503 41024
rect 5445 41015 5503 41021
rect 5534 41012 5540 41024
rect 5592 41012 5598 41064
rect 5721 41055 5779 41061
rect 5721 41021 5733 41055
rect 5767 41021 5779 41055
rect 6822 41052 6828 41064
rect 6783 41024 6828 41052
rect 5721 41015 5779 41021
rect 3602 40944 3608 40996
rect 3660 40984 3666 40996
rect 5736 40984 5764 41015
rect 6822 41012 6828 41024
rect 6880 41012 6886 41064
rect 7392 41061 7420 41228
rect 11054 41216 11060 41228
rect 11112 41216 11118 41268
rect 11330 41256 11336 41268
rect 11291 41228 11336 41256
rect 11330 41216 11336 41228
rect 11388 41216 11394 41268
rect 11422 41216 11428 41268
rect 11480 41256 11486 41268
rect 16758 41256 16764 41268
rect 11480 41228 16764 41256
rect 11480 41216 11486 41228
rect 16758 41216 16764 41228
rect 16816 41216 16822 41268
rect 18414 41216 18420 41268
rect 18472 41256 18478 41268
rect 27706 41256 27712 41268
rect 18472 41228 27108 41256
rect 27667 41228 27712 41256
rect 18472 41216 18478 41228
rect 12437 41191 12495 41197
rect 10520 41160 11744 41188
rect 7377 41055 7435 41061
rect 7377 41021 7389 41055
rect 7423 41021 7435 41055
rect 7377 41015 7435 41021
rect 9861 41055 9919 41061
rect 9861 41021 9873 41055
rect 9907 41052 9919 41055
rect 10137 41055 10195 41061
rect 10137 41052 10149 41055
rect 9907 41024 10149 41052
rect 9907 41021 9919 41024
rect 9861 41015 9919 41021
rect 10137 41021 10149 41024
rect 10183 41021 10195 41055
rect 10137 41015 10195 41021
rect 10321 41055 10379 41061
rect 10321 41021 10333 41055
rect 10367 41021 10379 41055
rect 10520 41052 10548 41160
rect 11716 41129 11744 41160
rect 12437 41157 12449 41191
rect 12483 41188 12495 41191
rect 16574 41188 16580 41200
rect 12483 41160 16580 41188
rect 12483 41157 12495 41160
rect 12437 41151 12495 41157
rect 16574 41148 16580 41160
rect 16632 41148 16638 41200
rect 27080 41188 27108 41228
rect 27706 41216 27712 41228
rect 27764 41216 27770 41268
rect 29365 41259 29423 41265
rect 29365 41225 29377 41259
rect 29411 41256 29423 41259
rect 30558 41256 30564 41268
rect 29411 41228 30564 41256
rect 29411 41225 29423 41228
rect 29365 41219 29423 41225
rect 30558 41216 30564 41228
rect 30616 41216 30622 41268
rect 38838 41216 38844 41268
rect 38896 41256 38902 41268
rect 39945 41259 40003 41265
rect 39945 41256 39957 41259
rect 38896 41228 39957 41256
rect 38896 41216 38902 41228
rect 39945 41225 39957 41228
rect 39991 41256 40003 41259
rect 40037 41259 40095 41265
rect 40037 41256 40049 41259
rect 39991 41228 40049 41256
rect 39991 41225 40003 41228
rect 39945 41219 40003 41225
rect 40037 41225 40049 41228
rect 40083 41225 40095 41259
rect 40218 41256 40224 41268
rect 40179 41228 40224 41256
rect 40037 41219 40095 41225
rect 40218 41216 40224 41228
rect 40276 41216 40282 41268
rect 42058 41256 42064 41268
rect 41971 41228 42064 41256
rect 42058 41216 42064 41228
rect 42116 41256 42122 41268
rect 42116 41228 47348 41256
rect 42116 41216 42122 41228
rect 45462 41188 45468 41200
rect 27080 41160 45468 41188
rect 45462 41148 45468 41160
rect 45520 41188 45526 41200
rect 46750 41188 46756 41200
rect 45520 41160 46756 41188
rect 45520 41148 45526 41160
rect 46750 41148 46756 41160
rect 46808 41188 46814 41200
rect 46845 41191 46903 41197
rect 46845 41188 46857 41191
rect 46808 41160 46857 41188
rect 46808 41148 46814 41160
rect 46845 41157 46857 41160
rect 46891 41188 46903 41191
rect 47320 41188 47348 41228
rect 49602 41216 49608 41268
rect 49660 41256 49666 41268
rect 53377 41259 53435 41265
rect 53377 41256 53389 41259
rect 49660 41228 53389 41256
rect 49660 41216 49666 41228
rect 53377 41225 53389 41228
rect 53423 41225 53435 41259
rect 53377 41219 53435 41225
rect 55858 41216 55864 41268
rect 55916 41256 55922 41268
rect 72786 41256 72792 41268
rect 55916 41228 72648 41256
rect 72747 41228 72792 41256
rect 55916 41216 55922 41228
rect 59170 41188 59176 41200
rect 46891 41160 47256 41188
rect 47320 41160 59176 41188
rect 46891 41157 46903 41160
rect 46845 41151 46903 41157
rect 11701 41123 11759 41129
rect 11701 41089 11713 41123
rect 11747 41120 11759 41123
rect 17402 41120 17408 41132
rect 11747 41092 12756 41120
rect 11747 41089 11759 41092
rect 11701 41083 11759 41089
rect 12728 41064 12756 41092
rect 12820 41092 17408 41120
rect 10781 41055 10839 41061
rect 10781 41052 10793 41055
rect 10520 41024 10793 41052
rect 10321 41015 10379 41021
rect 10781 41021 10793 41024
rect 10827 41021 10839 41055
rect 10781 41015 10839 41021
rect 10873 41055 10931 41061
rect 10873 41021 10885 41055
rect 10919 41052 10931 41055
rect 12437 41055 12495 41061
rect 12437 41052 12449 41055
rect 10919 41024 12449 41052
rect 10919 41021 10931 41024
rect 10873 41015 10931 41021
rect 12437 41021 12449 41024
rect 12483 41021 12495 41055
rect 12710 41052 12716 41064
rect 12671 41024 12716 41052
rect 12437 41015 12495 41021
rect 10336 40984 10364 41015
rect 10888 40984 10916 41015
rect 12710 41012 12716 41024
rect 12768 41012 12774 41064
rect 12820 40984 12848 41092
rect 17402 41080 17408 41092
rect 17460 41080 17466 41132
rect 18690 41120 18696 41132
rect 18651 41092 18696 41120
rect 18690 41080 18696 41092
rect 18748 41080 18754 41132
rect 19426 41120 19432 41132
rect 19387 41092 19432 41120
rect 19426 41080 19432 41092
rect 19484 41080 19490 41132
rect 23750 41080 23756 41132
rect 23808 41120 23814 41132
rect 23937 41123 23995 41129
rect 23937 41120 23949 41123
rect 23808 41092 23949 41120
rect 23808 41080 23814 41092
rect 23937 41089 23949 41092
rect 23983 41089 23995 41123
rect 23937 41083 23995 41089
rect 25225 41123 25283 41129
rect 25225 41089 25237 41123
rect 25271 41120 25283 41123
rect 26421 41123 26479 41129
rect 26421 41120 26433 41123
rect 25271 41092 26433 41120
rect 25271 41089 25283 41092
rect 25225 41083 25283 41089
rect 26421 41089 26433 41092
rect 26467 41089 26479 41123
rect 26421 41083 26479 41089
rect 26510 41080 26516 41132
rect 26568 41120 26574 41132
rect 29365 41123 29423 41129
rect 29365 41120 29377 41123
rect 26568 41092 29377 41120
rect 26568 41080 26574 41092
rect 29365 41089 29377 41092
rect 29411 41089 29423 41123
rect 29733 41123 29791 41129
rect 29733 41120 29745 41123
rect 29365 41083 29423 41089
rect 29472 41092 29745 41120
rect 13446 41052 13452 41064
rect 13407 41024 13452 41052
rect 13446 41012 13452 41024
rect 13504 41012 13510 41064
rect 13633 41055 13691 41061
rect 13633 41021 13645 41055
rect 13679 41052 13691 41055
rect 13722 41052 13728 41064
rect 13679 41024 13728 41052
rect 13679 41021 13691 41024
rect 13633 41015 13691 41021
rect 13722 41012 13728 41024
rect 13780 41012 13786 41064
rect 13998 41052 14004 41064
rect 13959 41024 14004 41052
rect 13998 41012 14004 41024
rect 14056 41012 14062 41064
rect 14185 41055 14243 41061
rect 14185 41021 14197 41055
rect 14231 41021 14243 41055
rect 14185 41015 14243 41021
rect 3660 40956 5304 40984
rect 5736 40956 10272 40984
rect 10336 40956 10916 40984
rect 10980 40956 12848 40984
rect 12897 40987 12955 40993
rect 3660 40944 3666 40956
rect 5276 40925 5304 40956
rect 5261 40919 5319 40925
rect 5261 40885 5273 40919
rect 5307 40885 5319 40919
rect 5261 40879 5319 40885
rect 6917 40919 6975 40925
rect 6917 40885 6929 40919
rect 6963 40916 6975 40919
rect 7006 40916 7012 40928
rect 6963 40888 7012 40916
rect 6963 40885 6975 40888
rect 6917 40879 6975 40885
rect 7006 40876 7012 40888
rect 7064 40876 7070 40928
rect 7558 40876 7564 40928
rect 7616 40916 7622 40928
rect 9861 40919 9919 40925
rect 9861 40916 9873 40919
rect 7616 40888 9873 40916
rect 7616 40876 7622 40888
rect 9861 40885 9873 40888
rect 9907 40916 9919 40919
rect 9953 40919 10011 40925
rect 9953 40916 9965 40919
rect 9907 40888 9965 40916
rect 9907 40885 9919 40888
rect 9861 40879 9919 40885
rect 9953 40885 9965 40888
rect 9999 40885 10011 40919
rect 10244 40916 10272 40956
rect 10980 40916 11008 40956
rect 12897 40953 12909 40987
rect 12943 40984 12955 40987
rect 14200 40984 14228 41015
rect 19242 41012 19248 41064
rect 19300 41052 19306 41064
rect 19337 41055 19395 41061
rect 19337 41052 19349 41055
rect 19300 41024 19349 41052
rect 19300 41012 19306 41024
rect 19337 41021 19349 41024
rect 19383 41021 19395 41055
rect 19337 41015 19395 41021
rect 19705 41055 19763 41061
rect 19705 41021 19717 41055
rect 19751 41021 19763 41055
rect 19705 41015 19763 41021
rect 19889 41055 19947 41061
rect 19889 41021 19901 41055
rect 19935 41052 19947 41055
rect 19935 41024 24072 41052
rect 19935 41021 19947 41024
rect 19889 41015 19947 41021
rect 12943 40956 14228 40984
rect 12943 40953 12955 40956
rect 12897 40947 12955 40953
rect 10244 40888 11008 40916
rect 9953 40879 10011 40885
rect 11054 40876 11060 40928
rect 11112 40916 11118 40928
rect 12912 40916 12940 40947
rect 13078 40916 13084 40928
rect 11112 40888 12940 40916
rect 13039 40888 13084 40916
rect 11112 40876 11118 40888
rect 13078 40876 13084 40888
rect 13136 40876 13142 40928
rect 14200 40916 14228 40956
rect 19426 40944 19432 40996
rect 19484 40984 19490 40996
rect 19720 40984 19748 41015
rect 19484 40956 19748 40984
rect 24044 40984 24072 41024
rect 24118 41012 24124 41064
rect 24176 41052 24182 41064
rect 24670 41052 24676 41064
rect 24176 41024 24676 41052
rect 24176 41012 24182 41024
rect 24670 41012 24676 41024
rect 24728 41012 24734 41064
rect 24857 41055 24915 41061
rect 24857 41021 24869 41055
rect 24903 41021 24915 41055
rect 26142 41052 26148 41064
rect 26103 41024 26148 41052
rect 24857 41015 24915 41021
rect 24872 40984 24900 41015
rect 26142 41012 26148 41024
rect 26200 41012 26206 41064
rect 27982 41052 27988 41064
rect 26252 41024 27988 41052
rect 26252 40984 26280 41024
rect 27982 41012 27988 41024
rect 28040 41012 28046 41064
rect 24044 40956 26280 40984
rect 19484 40944 19490 40956
rect 21818 40916 21824 40928
rect 14200 40888 21824 40916
rect 21818 40876 21824 40888
rect 21876 40876 21882 40928
rect 23750 40916 23756 40928
rect 23711 40888 23756 40916
rect 23750 40876 23756 40888
rect 23808 40876 23814 40928
rect 26142 40876 26148 40928
rect 26200 40916 26206 40928
rect 27890 40916 27896 40928
rect 26200 40888 27896 40916
rect 26200 40876 26206 40888
rect 27890 40876 27896 40888
rect 27948 40876 27954 40928
rect 29178 40876 29184 40928
rect 29236 40916 29242 40928
rect 29472 40925 29500 41092
rect 29733 41089 29745 41092
rect 29779 41089 29791 41123
rect 29733 41083 29791 41089
rect 39485 41123 39543 41129
rect 39485 41089 39497 41123
rect 39531 41120 39543 41123
rect 40402 41120 40408 41132
rect 39531 41092 40408 41120
rect 39531 41089 39543 41092
rect 39485 41083 39543 41089
rect 40402 41080 40408 41092
rect 40460 41080 40466 41132
rect 40586 41080 40592 41132
rect 40644 41120 40650 41132
rect 41690 41120 41696 41132
rect 40644 41092 40908 41120
rect 41651 41092 41696 41120
rect 40644 41080 40650 41092
rect 29638 41012 29644 41064
rect 29696 41052 29702 41064
rect 29825 41055 29883 41061
rect 29825 41052 29837 41055
rect 29696 41024 29837 41052
rect 29696 41012 29702 41024
rect 29825 41021 29837 41024
rect 29871 41052 29883 41055
rect 30377 41055 30435 41061
rect 30377 41052 30389 41055
rect 29871 41024 30389 41052
rect 29871 41021 29883 41024
rect 29825 41015 29883 41021
rect 30377 41021 30389 41024
rect 30423 41021 30435 41055
rect 30558 41052 30564 41064
rect 30471 41024 30564 41052
rect 30377 41015 30435 41021
rect 30558 41012 30564 41024
rect 30616 41052 30622 41064
rect 31205 41055 31263 41061
rect 31205 41052 31217 41055
rect 30616 41024 31217 41052
rect 30616 41012 30622 41024
rect 31205 41021 31217 41024
rect 31251 41052 31263 41055
rect 31251 41024 33548 41052
rect 31251 41021 31263 41024
rect 31205 41015 31263 41021
rect 30929 40987 30987 40993
rect 30929 40953 30941 40987
rect 30975 40984 30987 40987
rect 33410 40984 33416 40996
rect 30975 40956 33416 40984
rect 30975 40953 30987 40956
rect 30929 40947 30987 40953
rect 33410 40944 33416 40956
rect 33468 40944 33474 40996
rect 33520 40984 33548 41024
rect 38010 41012 38016 41064
rect 38068 41052 38074 41064
rect 38197 41055 38255 41061
rect 38197 41052 38209 41055
rect 38068 41024 38209 41052
rect 38068 41012 38074 41024
rect 38197 41021 38209 41024
rect 38243 41021 38255 41055
rect 38197 41015 38255 41021
rect 38381 41055 38439 41061
rect 38381 41021 38393 41055
rect 38427 41052 38439 41055
rect 38746 41052 38752 41064
rect 38427 41024 38752 41052
rect 38427 41021 38439 41024
rect 38381 41015 38439 41021
rect 38746 41012 38752 41024
rect 38804 41012 38810 41064
rect 38841 41055 38899 41061
rect 38841 41021 38853 41055
rect 38887 41052 38899 41055
rect 39021 41055 39079 41061
rect 38887 41024 38976 41052
rect 38887 41021 38899 41024
rect 38841 41015 38899 41021
rect 38654 40984 38660 40996
rect 33520 40956 38660 40984
rect 38654 40944 38660 40956
rect 38712 40944 38718 40996
rect 38948 40984 38976 41024
rect 39021 41021 39033 41055
rect 39067 41052 39079 41055
rect 39390 41052 39396 41064
rect 39067 41024 39396 41052
rect 39067 41021 39079 41024
rect 39021 41015 39079 41021
rect 39390 41012 39396 41024
rect 39448 41012 39454 41064
rect 40497 41055 40555 41061
rect 40497 41052 40509 41055
rect 39960 41024 40509 41052
rect 39114 40984 39120 40996
rect 38948 40956 39120 40984
rect 39114 40944 39120 40956
rect 39172 40984 39178 40996
rect 39960 40984 39988 41024
rect 40497 41021 40509 41024
rect 40543 41021 40555 41055
rect 40497 41015 40555 41021
rect 40681 41055 40739 41061
rect 40681 41021 40693 41055
rect 40727 41021 40739 41055
rect 40880 41052 40908 41092
rect 41690 41080 41696 41092
rect 41748 41080 41754 41132
rect 47228 41129 47256 41160
rect 59170 41148 59176 41160
rect 59228 41148 59234 41200
rect 60826 41188 60832 41200
rect 60787 41160 60832 41188
rect 60826 41148 60832 41160
rect 60884 41148 60890 41200
rect 61102 41188 61108 41200
rect 61015 41160 61108 41188
rect 61102 41148 61108 41160
rect 61160 41188 61166 41200
rect 64322 41188 64328 41200
rect 61160 41160 64328 41188
rect 61160 41148 61166 41160
rect 64322 41148 64328 41160
rect 64380 41148 64386 41200
rect 65429 41191 65487 41197
rect 65429 41157 65441 41191
rect 65475 41188 65487 41191
rect 66438 41188 66444 41200
rect 65475 41160 66444 41188
rect 65475 41157 65487 41160
rect 65429 41151 65487 41157
rect 66438 41148 66444 41160
rect 66496 41148 66502 41200
rect 72237 41191 72295 41197
rect 72237 41157 72249 41191
rect 72283 41157 72295 41191
rect 72620 41188 72648 41228
rect 72786 41216 72792 41228
rect 72844 41216 72850 41268
rect 83185 41191 83243 41197
rect 83185 41188 83197 41191
rect 72620 41160 83197 41188
rect 72237 41151 72295 41157
rect 83185 41157 83197 41160
rect 83231 41188 83243 41191
rect 83734 41188 83740 41200
rect 83231 41160 83740 41188
rect 83231 41157 83243 41160
rect 83185 41151 83243 41157
rect 47213 41123 47271 41129
rect 47213 41089 47225 41123
rect 47259 41089 47271 41123
rect 47213 41083 47271 41089
rect 48501 41123 48559 41129
rect 48501 41089 48513 41123
rect 48547 41089 48559 41123
rect 48501 41083 48559 41089
rect 41141 41055 41199 41061
rect 41141 41052 41153 41055
rect 40880 41024 41153 41052
rect 40681 41015 40739 41021
rect 41141 41021 41153 41024
rect 41187 41021 41199 41055
rect 41141 41015 41199 41021
rect 39172 40956 39988 40984
rect 40037 40987 40095 40993
rect 39172 40944 39178 40956
rect 40037 40953 40049 40987
rect 40083 40984 40095 40987
rect 40586 40984 40592 40996
rect 40083 40956 40592 40984
rect 40083 40953 40095 40956
rect 40037 40947 40095 40953
rect 40586 40944 40592 40956
rect 40644 40944 40650 40996
rect 40696 40984 40724 41015
rect 41230 41012 41236 41064
rect 41288 41052 41294 41064
rect 41288 41024 41333 41052
rect 41288 41012 41294 41024
rect 41414 41012 41420 41064
rect 41472 41052 41478 41064
rect 47029 41055 47087 41061
rect 47029 41052 47041 41055
rect 41472 41024 47041 41052
rect 41472 41012 41478 41024
rect 47029 41021 47041 41024
rect 47075 41021 47087 41055
rect 47394 41052 47400 41064
rect 47355 41024 47400 41052
rect 47029 41015 47087 41021
rect 42058 40984 42064 40996
rect 40696 40956 42064 40984
rect 42058 40944 42064 40956
rect 42116 40944 42122 40996
rect 47044 40984 47072 41015
rect 47394 41012 47400 41024
rect 47452 41012 47458 41064
rect 47857 41055 47915 41061
rect 47857 41021 47869 41055
rect 47903 41021 47915 41055
rect 47857 41015 47915 41021
rect 47949 41055 48007 41061
rect 47949 41021 47961 41055
rect 47995 41021 48007 41055
rect 48516 41052 48544 41083
rect 53190 41080 53196 41132
rect 53248 41129 53254 41132
rect 53248 41123 53306 41129
rect 53248 41089 53260 41123
rect 53294 41089 53306 41123
rect 53466 41120 53472 41132
rect 53427 41092 53472 41120
rect 53248 41083 53306 41089
rect 53248 41080 53254 41083
rect 53466 41080 53472 41092
rect 53524 41080 53530 41132
rect 59262 41120 59268 41132
rect 59223 41092 59268 41120
rect 59262 41080 59268 41092
rect 59320 41080 59326 41132
rect 59538 41120 59544 41132
rect 59499 41092 59544 41120
rect 59538 41080 59544 41092
rect 59596 41080 59602 41132
rect 66349 41123 66407 41129
rect 66349 41089 66361 41123
rect 66395 41120 66407 41123
rect 66898 41120 66904 41132
rect 66395 41092 66904 41120
rect 66395 41089 66407 41092
rect 66349 41083 66407 41089
rect 66898 41080 66904 41092
rect 66956 41080 66962 41132
rect 71866 41080 71872 41132
rect 71924 41120 71930 41132
rect 72108 41123 72166 41129
rect 71924 41092 72004 41120
rect 71924 41080 71930 41092
rect 53101 41055 53159 41061
rect 53101 41052 53113 41055
rect 48516 41024 53113 41052
rect 47949 41015 48007 41021
rect 53101 41021 53113 41024
rect 53147 41021 53159 41055
rect 53101 41015 53159 41021
rect 58805 41055 58863 41061
rect 58805 41021 58817 41055
rect 58851 41052 58863 41055
rect 58894 41052 58900 41064
rect 58851 41024 58900 41052
rect 58851 41021 58863 41024
rect 58805 41015 58863 41021
rect 47872 40984 47900 41015
rect 47044 40956 47900 40984
rect 47964 40984 47992 41015
rect 58894 41012 58900 41024
rect 58952 41052 58958 41064
rect 59057 41055 59115 41061
rect 59057 41052 59069 41055
rect 58952 41024 59069 41052
rect 58952 41012 58958 41024
rect 59057 41021 59069 41024
rect 59103 41021 59115 41055
rect 65334 41052 65340 41064
rect 65295 41024 65340 41052
rect 59057 41015 59115 41021
rect 65334 41012 65340 41024
rect 65392 41052 65398 41064
rect 65613 41055 65671 41061
rect 65613 41052 65625 41055
rect 65392 41024 65625 41052
rect 65392 41012 65398 41024
rect 65613 41021 65625 41024
rect 65659 41052 65671 41055
rect 65978 41052 65984 41064
rect 65659 41024 65984 41052
rect 65659 41021 65671 41024
rect 65613 41015 65671 41021
rect 65978 41012 65984 41024
rect 66036 41012 66042 41064
rect 66622 41052 66628 41064
rect 66583 41024 66628 41052
rect 66622 41012 66628 41024
rect 66680 41012 66686 41064
rect 66824 41024 67220 41052
rect 48222 40984 48228 40996
rect 47964 40956 48228 40984
rect 29457 40919 29515 40925
rect 29457 40916 29469 40919
rect 29236 40888 29469 40916
rect 29236 40876 29242 40888
rect 29457 40885 29469 40888
rect 29503 40885 29515 40919
rect 38010 40916 38016 40928
rect 37971 40888 38016 40916
rect 29457 40879 29515 40885
rect 38010 40876 38016 40888
rect 38068 40876 38074 40928
rect 39298 40876 39304 40928
rect 39356 40916 39362 40928
rect 39574 40916 39580 40928
rect 39356 40888 39580 40916
rect 39356 40876 39362 40888
rect 39574 40876 39580 40888
rect 39632 40876 39638 40928
rect 39761 40919 39819 40925
rect 39761 40885 39773 40919
rect 39807 40916 39819 40919
rect 40218 40916 40224 40928
rect 39807 40888 40224 40916
rect 39807 40885 39819 40888
rect 39761 40879 39819 40885
rect 40218 40876 40224 40888
rect 40276 40876 40282 40928
rect 41046 40876 41052 40928
rect 41104 40916 41110 40928
rect 47964 40916 47992 40956
rect 48222 40944 48228 40956
rect 48280 40984 48286 40996
rect 48869 40987 48927 40993
rect 48869 40984 48881 40987
rect 48280 40956 48881 40984
rect 48280 40944 48286 40956
rect 48869 40953 48881 40956
rect 48915 40953 48927 40987
rect 66533 40987 66591 40993
rect 48869 40947 48927 40953
rect 53668 40956 59032 40984
rect 41104 40888 47992 40916
rect 41104 40876 41110 40888
rect 48130 40876 48136 40928
rect 48188 40916 48194 40928
rect 48685 40919 48743 40925
rect 48685 40916 48697 40919
rect 48188 40888 48697 40916
rect 48188 40876 48194 40888
rect 48685 40885 48697 40888
rect 48731 40916 48743 40919
rect 48774 40916 48780 40928
rect 48731 40888 48780 40916
rect 48731 40885 48743 40888
rect 48685 40879 48743 40885
rect 48774 40876 48780 40888
rect 48832 40876 48838 40928
rect 48884 40916 48912 40947
rect 53668 40916 53696 40956
rect 48884 40888 53696 40916
rect 53745 40919 53803 40925
rect 53745 40885 53757 40919
rect 53791 40916 53803 40919
rect 54478 40916 54484 40928
rect 53791 40888 54484 40916
rect 53791 40885 53803 40888
rect 53745 40879 53803 40885
rect 54478 40876 54484 40888
rect 54536 40876 54542 40928
rect 58710 40876 58716 40928
rect 58768 40916 58774 40928
rect 58897 40919 58955 40925
rect 58897 40916 58909 40919
rect 58768 40888 58909 40916
rect 58768 40876 58774 40888
rect 58897 40885 58909 40888
rect 58943 40885 58955 40919
rect 59004 40916 59032 40956
rect 66533 40953 66545 40987
rect 66579 40984 66591 40987
rect 66714 40984 66720 40996
rect 66579 40956 66720 40984
rect 66579 40953 66591 40956
rect 66533 40947 66591 40953
rect 66714 40944 66720 40956
rect 66772 40944 66778 40996
rect 66824 40916 66852 41024
rect 67082 40984 67088 40996
rect 67043 40956 67088 40984
rect 67082 40944 67088 40956
rect 67140 40944 67146 40996
rect 67192 40984 67220 41024
rect 67358 41012 67364 41064
rect 67416 41052 67422 41064
rect 71590 41052 71596 41064
rect 67416 41024 71596 41052
rect 67416 41012 67422 41024
rect 71590 41012 71596 41024
rect 71648 41012 71654 41064
rect 71976 41061 72004 41092
rect 72108 41089 72120 41123
rect 72154 41120 72166 41123
rect 72252 41120 72280 41151
rect 83734 41148 83740 41160
rect 83792 41148 83798 41200
rect 72418 41120 72424 41132
rect 72154 41089 72188 41120
rect 72252 41092 72424 41120
rect 72108 41083 72188 41089
rect 71961 41055 72019 41061
rect 71961 41021 71973 41055
rect 72007 41021 72019 41055
rect 71961 41015 72019 41021
rect 71682 40984 71688 40996
rect 67192 40956 71688 40984
rect 71682 40944 71688 40956
rect 71740 40944 71746 40996
rect 72160 40984 72188 41083
rect 72418 41080 72424 41092
rect 72476 41080 72482 41132
rect 72694 41120 72700 41132
rect 72655 41092 72700 41120
rect 72694 41080 72700 41092
rect 72752 41080 72758 41132
rect 76285 41123 76343 41129
rect 76285 41120 76297 41123
rect 75196 41092 76297 41120
rect 72326 41061 72332 41064
rect 72300 41055 72332 41061
rect 72300 41021 72312 41055
rect 72300 41015 72332 41021
rect 72326 41012 72332 41015
rect 72384 41012 72390 41064
rect 75196 41052 75224 41092
rect 76285 41089 76297 41092
rect 76331 41120 76343 41123
rect 77573 41123 77631 41129
rect 76331 41092 77340 41120
rect 76331 41089 76343 41092
rect 76285 41083 76343 41089
rect 76190 41052 76196 41064
rect 72436 41024 75224 41052
rect 76151 41024 76196 41052
rect 72436 40984 72464 41024
rect 76190 41012 76196 41024
rect 76248 41052 76254 41064
rect 76469 41055 76527 41061
rect 76469 41052 76481 41055
rect 76248 41024 76481 41052
rect 76248 41012 76254 41024
rect 76469 41021 76481 41024
rect 76515 41021 76527 41055
rect 77202 41052 77208 41064
rect 77163 41024 77208 41052
rect 76469 41015 76527 41021
rect 77202 41012 77208 41024
rect 77260 41012 77266 41064
rect 77312 41052 77340 41092
rect 77573 41089 77585 41123
rect 77619 41120 77631 41123
rect 77662 41120 77668 41132
rect 77619 41092 77668 41120
rect 77619 41089 77631 41092
rect 77573 41083 77631 41089
rect 77662 41080 77668 41092
rect 77720 41080 77726 41132
rect 77478 41052 77484 41064
rect 77312 41024 77484 41052
rect 77478 41012 77484 41024
rect 77536 41052 77542 41064
rect 77757 41055 77815 41061
rect 77757 41052 77769 41055
rect 77536 41024 77769 41052
rect 77536 41012 77542 41024
rect 77757 41021 77769 41024
rect 77803 41021 77815 41055
rect 77757 41015 77815 41021
rect 83001 41055 83059 41061
rect 83001 41021 83013 41055
rect 83047 41021 83059 41055
rect 83001 41015 83059 41021
rect 72160 40956 72464 40984
rect 72510 40944 72516 40996
rect 72568 40984 72574 40996
rect 83016 40984 83044 41015
rect 83369 40987 83427 40993
rect 83369 40984 83381 40987
rect 72568 40956 83381 40984
rect 72568 40944 72574 40956
rect 83369 40953 83381 40956
rect 83415 40984 83427 40987
rect 84102 40984 84108 40996
rect 83415 40956 84108 40984
rect 83415 40953 83427 40956
rect 83369 40947 83427 40953
rect 84102 40944 84108 40956
rect 84160 40944 84166 40996
rect 59004 40888 66852 40916
rect 58897 40879 58955 40885
rect 66898 40876 66904 40928
rect 66956 40916 66962 40928
rect 67269 40919 67327 40925
rect 67269 40916 67281 40919
rect 66956 40888 67281 40916
rect 66956 40876 66962 40888
rect 67269 40885 67281 40888
rect 67315 40916 67327 40919
rect 67634 40916 67640 40928
rect 67315 40888 67640 40916
rect 67315 40885 67327 40888
rect 67269 40879 67327 40885
rect 67634 40876 67640 40888
rect 67692 40876 67698 40928
rect 71774 40916 71780 40928
rect 71735 40888 71780 40916
rect 71774 40876 71780 40888
rect 71832 40876 71838 40928
rect 76190 40876 76196 40928
rect 76248 40916 76254 40928
rect 78950 40916 78956 40928
rect 76248 40888 78956 40916
rect 76248 40876 76254 40888
rect 78950 40876 78956 40888
rect 79008 40876 79014 40928
rect 1104 40826 108008 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 81046 40826
rect 81098 40774 81110 40826
rect 81162 40774 81174 40826
rect 81226 40774 81238 40826
rect 81290 40774 108008 40826
rect 1104 40752 108008 40774
rect 7285 40715 7343 40721
rect 7285 40681 7297 40715
rect 7331 40712 7343 40715
rect 7742 40712 7748 40724
rect 7331 40684 7748 40712
rect 7331 40681 7343 40684
rect 7285 40675 7343 40681
rect 7742 40672 7748 40684
rect 7800 40672 7806 40724
rect 10134 40672 10140 40724
rect 10192 40712 10198 40724
rect 11054 40712 11060 40724
rect 10192 40684 11060 40712
rect 10192 40672 10198 40684
rect 11054 40672 11060 40684
rect 11112 40672 11118 40724
rect 12621 40715 12679 40721
rect 12621 40681 12633 40715
rect 12667 40712 12679 40715
rect 12710 40712 12716 40724
rect 12667 40684 12716 40712
rect 12667 40681 12679 40684
rect 12621 40675 12679 40681
rect 12710 40672 12716 40684
rect 12768 40712 12774 40724
rect 13446 40712 13452 40724
rect 12768 40684 13452 40712
rect 12768 40672 12774 40684
rect 13446 40672 13452 40684
rect 13504 40712 13510 40724
rect 27249 40715 27307 40721
rect 13504 40684 27200 40712
rect 13504 40672 13510 40684
rect 5534 40604 5540 40656
rect 5592 40644 5598 40656
rect 13078 40644 13084 40656
rect 5592 40616 6868 40644
rect 5592 40604 5598 40616
rect 5736 40585 5764 40616
rect 6840 40588 6868 40616
rect 7576 40616 13084 40644
rect 5721 40579 5779 40585
rect 5721 40545 5733 40579
rect 5767 40545 5779 40579
rect 5721 40539 5779 40545
rect 5997 40579 6055 40585
rect 5997 40545 6009 40579
rect 6043 40545 6055 40579
rect 5997 40539 6055 40545
rect 3050 40468 3056 40520
rect 3108 40508 3114 40520
rect 5905 40511 5963 40517
rect 5905 40508 5917 40511
rect 3108 40480 5917 40508
rect 3108 40468 3114 40480
rect 5905 40477 5917 40480
rect 5951 40477 5963 40511
rect 6012 40508 6040 40539
rect 6822 40536 6828 40588
rect 6880 40576 6886 40588
rect 7576 40585 7604 40616
rect 13078 40604 13084 40616
rect 13136 40604 13142 40656
rect 13538 40604 13544 40656
rect 13596 40644 13602 40656
rect 15565 40647 15623 40653
rect 15565 40644 15577 40647
rect 13596 40616 15577 40644
rect 13596 40604 13602 40616
rect 15565 40613 15577 40616
rect 15611 40644 15623 40647
rect 15611 40616 15792 40644
rect 15611 40613 15623 40616
rect 15565 40607 15623 40613
rect 7009 40579 7067 40585
rect 7009 40576 7021 40579
rect 6880 40548 7021 40576
rect 6880 40536 6886 40548
rect 7009 40545 7021 40548
rect 7055 40545 7067 40579
rect 7009 40539 7067 40545
rect 7561 40579 7619 40585
rect 7561 40545 7573 40579
rect 7607 40545 7619 40579
rect 9493 40579 9551 40585
rect 9493 40576 9505 40579
rect 7561 40539 7619 40545
rect 7760 40548 9505 40576
rect 7760 40508 7788 40548
rect 9493 40545 9505 40548
rect 9539 40545 9551 40579
rect 10226 40576 10232 40588
rect 10187 40548 10232 40576
rect 9493 40539 9551 40545
rect 10226 40536 10232 40548
rect 10284 40536 10290 40588
rect 12526 40576 12532 40588
rect 12487 40548 12532 40576
rect 12526 40536 12532 40548
rect 12584 40536 12590 40588
rect 15764 40585 15792 40616
rect 19242 40604 19248 40656
rect 19300 40604 19306 40656
rect 20346 40644 20352 40656
rect 19904 40616 20352 40644
rect 15749 40579 15807 40585
rect 15749 40545 15761 40579
rect 15795 40545 15807 40579
rect 18785 40579 18843 40585
rect 18785 40576 18797 40579
rect 15749 40539 15807 40545
rect 15856 40548 18797 40576
rect 6012 40480 7788 40508
rect 5905 40471 5963 40477
rect 7834 40468 7840 40520
rect 7892 40508 7898 40520
rect 11422 40508 11428 40520
rect 7892 40480 11428 40508
rect 7892 40468 7898 40480
rect 11422 40468 11428 40480
rect 11480 40468 11486 40520
rect 15856 40508 15884 40548
rect 18785 40545 18797 40548
rect 18831 40545 18843 40579
rect 19260 40576 19288 40604
rect 19429 40579 19487 40585
rect 19429 40576 19441 40579
rect 19260 40548 19441 40576
rect 18785 40539 18843 40545
rect 19429 40545 19441 40548
rect 19475 40545 19487 40579
rect 19429 40539 19487 40545
rect 19518 40536 19524 40588
rect 19576 40576 19582 40588
rect 19797 40579 19855 40585
rect 19797 40576 19809 40579
rect 19576 40548 19809 40576
rect 19576 40536 19582 40548
rect 19797 40545 19809 40548
rect 19843 40545 19855 40579
rect 19797 40539 19855 40545
rect 16022 40508 16028 40520
rect 11532 40480 15884 40508
rect 15983 40480 16028 40508
rect 9493 40443 9551 40449
rect 9493 40409 9505 40443
rect 9539 40440 9551 40443
rect 11532 40440 11560 40480
rect 16022 40468 16028 40480
rect 16080 40468 16086 40520
rect 17405 40511 17463 40517
rect 17405 40477 17417 40511
rect 17451 40508 17463 40511
rect 18414 40508 18420 40520
rect 17451 40480 18420 40508
rect 17451 40477 17463 40480
rect 17405 40471 17463 40477
rect 18414 40468 18420 40480
rect 18472 40468 18478 40520
rect 19337 40511 19395 40517
rect 19337 40477 19349 40511
rect 19383 40508 19395 40511
rect 19904 40508 19932 40616
rect 20346 40604 20352 40616
rect 20404 40604 20410 40656
rect 26970 40604 26976 40656
rect 27028 40644 27034 40656
rect 27065 40647 27123 40653
rect 27065 40644 27077 40647
rect 27028 40616 27077 40644
rect 27028 40604 27034 40616
rect 27065 40613 27077 40616
rect 27111 40613 27123 40647
rect 27172 40644 27200 40684
rect 27249 40681 27261 40715
rect 27295 40712 27307 40715
rect 27338 40712 27344 40724
rect 27295 40684 27344 40712
rect 27295 40681 27307 40684
rect 27249 40675 27307 40681
rect 27338 40672 27344 40684
rect 27396 40672 27402 40724
rect 27430 40672 27436 40724
rect 27488 40712 27494 40724
rect 41506 40712 41512 40724
rect 27488 40684 41512 40712
rect 27488 40672 27494 40684
rect 41506 40672 41512 40684
rect 41564 40672 41570 40724
rect 41598 40672 41604 40724
rect 41656 40712 41662 40724
rect 55858 40712 55864 40724
rect 41656 40684 55864 40712
rect 41656 40672 41662 40684
rect 55858 40672 55864 40684
rect 55916 40672 55922 40724
rect 58434 40712 58440 40724
rect 58395 40684 58440 40712
rect 58434 40672 58440 40684
rect 58492 40672 58498 40724
rect 58894 40672 58900 40724
rect 58952 40712 58958 40724
rect 65426 40712 65432 40724
rect 58952 40684 65432 40712
rect 58952 40672 58958 40684
rect 65426 40672 65432 40684
rect 65484 40672 65490 40724
rect 71682 40672 71688 40724
rect 71740 40712 71746 40724
rect 76190 40712 76196 40724
rect 71740 40684 76196 40712
rect 71740 40672 71746 40684
rect 76190 40672 76196 40684
rect 76248 40672 76254 40724
rect 77665 40715 77723 40721
rect 77665 40681 77677 40715
rect 77711 40712 77723 40715
rect 77754 40712 77760 40724
rect 77711 40684 77760 40712
rect 77711 40681 77723 40684
rect 77665 40675 77723 40681
rect 77754 40672 77760 40684
rect 77812 40672 77818 40724
rect 84102 40672 84108 40724
rect 84160 40712 84166 40724
rect 84657 40715 84715 40721
rect 84657 40712 84669 40715
rect 84160 40684 84669 40712
rect 84160 40672 84166 40684
rect 84657 40681 84669 40684
rect 84703 40681 84715 40715
rect 84657 40675 84715 40681
rect 27172 40616 27384 40644
rect 27065 40607 27123 40613
rect 19981 40579 20039 40585
rect 19981 40545 19993 40579
rect 20027 40576 20039 40579
rect 20165 40579 20223 40585
rect 20165 40576 20177 40579
rect 20027 40548 20177 40576
rect 20027 40545 20039 40548
rect 19981 40539 20039 40545
rect 20165 40545 20177 40548
rect 20211 40576 20223 40579
rect 26605 40579 26663 40585
rect 20211 40548 26464 40576
rect 20211 40545 20223 40548
rect 20165 40539 20223 40545
rect 19383 40480 19932 40508
rect 19383 40477 19395 40480
rect 19337 40471 19395 40477
rect 21910 40468 21916 40520
rect 21968 40508 21974 40520
rect 22097 40511 22155 40517
rect 22097 40508 22109 40511
rect 21968 40480 22109 40508
rect 21968 40468 21974 40480
rect 22097 40477 22109 40480
rect 22143 40477 22155 40511
rect 22370 40508 22376 40520
rect 22331 40480 22376 40508
rect 22097 40471 22155 40477
rect 22370 40468 22376 40480
rect 22428 40468 22434 40520
rect 9539 40412 11560 40440
rect 26436 40440 26464 40548
rect 26605 40545 26617 40579
rect 26651 40576 26663 40579
rect 27246 40576 27252 40588
rect 26651 40548 27252 40576
rect 26651 40545 26663 40548
rect 26605 40539 26663 40545
rect 27246 40536 27252 40548
rect 27304 40536 27310 40588
rect 27356 40576 27384 40616
rect 28994 40604 29000 40656
rect 29052 40644 29058 40656
rect 29052 40616 30144 40644
rect 29052 40604 29058 40616
rect 27356 40548 29040 40576
rect 26513 40511 26571 40517
rect 26513 40477 26525 40511
rect 26559 40508 26571 40511
rect 27982 40508 27988 40520
rect 26559 40480 27988 40508
rect 26559 40477 26571 40480
rect 26513 40471 26571 40477
rect 27982 40468 27988 40480
rect 28040 40468 28046 40520
rect 29012 40508 29040 40548
rect 29454 40536 29460 40588
rect 29512 40576 29518 40588
rect 29564 40585 29592 40616
rect 30116 40585 30144 40616
rect 34146 40604 34152 40656
rect 34204 40644 34210 40656
rect 40218 40644 40224 40656
rect 34204 40616 40080 40644
rect 40179 40616 40224 40644
rect 34204 40604 34210 40616
rect 29549 40579 29607 40585
rect 29549 40576 29561 40579
rect 29512 40548 29561 40576
rect 29512 40536 29518 40548
rect 29549 40545 29561 40548
rect 29595 40545 29607 40579
rect 30009 40579 30067 40585
rect 30009 40576 30021 40579
rect 29549 40539 29607 40545
rect 29656 40548 30021 40576
rect 29086 40508 29092 40520
rect 29012 40480 29092 40508
rect 29086 40468 29092 40480
rect 29144 40468 29150 40520
rect 29178 40468 29184 40520
rect 29236 40508 29242 40520
rect 29365 40511 29423 40517
rect 29365 40508 29377 40511
rect 29236 40480 29377 40508
rect 29236 40468 29242 40480
rect 29365 40477 29377 40480
rect 29411 40477 29423 40511
rect 29365 40471 29423 40477
rect 29656 40440 29684 40548
rect 30009 40545 30021 40548
rect 30055 40545 30067 40579
rect 30009 40539 30067 40545
rect 30101 40579 30159 40585
rect 30101 40545 30113 40579
rect 30147 40545 30159 40579
rect 38838 40576 38844 40588
rect 38799 40548 38844 40576
rect 30101 40539 30159 40545
rect 38838 40536 38844 40548
rect 38896 40536 38902 40588
rect 39390 40576 39396 40588
rect 39351 40548 39396 40576
rect 39390 40536 39396 40548
rect 39448 40536 39454 40588
rect 39574 40576 39580 40588
rect 39535 40548 39580 40576
rect 39574 40536 39580 40548
rect 39632 40536 39638 40588
rect 40052 40576 40080 40616
rect 40218 40604 40224 40616
rect 40276 40604 40282 40656
rect 40405 40647 40463 40653
rect 40405 40613 40417 40647
rect 40451 40644 40463 40647
rect 40678 40644 40684 40656
rect 40451 40616 40684 40644
rect 40451 40613 40463 40616
rect 40405 40607 40463 40613
rect 40678 40604 40684 40616
rect 40736 40604 40742 40656
rect 40770 40604 40776 40656
rect 40828 40644 40834 40656
rect 40865 40647 40923 40653
rect 40865 40644 40877 40647
rect 40828 40616 40877 40644
rect 40828 40604 40834 40616
rect 40865 40613 40877 40616
rect 40911 40613 40923 40647
rect 40865 40607 40923 40613
rect 40954 40604 40960 40656
rect 41012 40644 41018 40656
rect 52730 40644 52736 40656
rect 41012 40616 52736 40644
rect 41012 40604 41018 40616
rect 52730 40604 52736 40616
rect 52788 40604 52794 40656
rect 52822 40604 52828 40656
rect 52880 40644 52886 40656
rect 58713 40647 58771 40653
rect 58713 40644 58725 40647
rect 52880 40616 58725 40644
rect 52880 40604 52886 40616
rect 58713 40613 58725 40616
rect 58759 40644 58771 40647
rect 58802 40644 58808 40656
rect 58759 40616 58808 40644
rect 58759 40613 58771 40616
rect 58713 40607 58771 40613
rect 58802 40604 58808 40616
rect 58860 40604 58866 40656
rect 60277 40647 60335 40653
rect 60277 40613 60289 40647
rect 60323 40644 60335 40647
rect 61562 40644 61568 40656
rect 60323 40616 61568 40644
rect 60323 40613 60335 40616
rect 60277 40607 60335 40613
rect 61562 40604 61568 40616
rect 61620 40604 61626 40656
rect 82725 40647 82783 40653
rect 82725 40613 82737 40647
rect 82771 40644 82783 40647
rect 83642 40644 83648 40656
rect 82771 40616 83648 40644
rect 82771 40613 82783 40616
rect 82725 40607 82783 40613
rect 83642 40604 83648 40616
rect 83700 40604 83706 40656
rect 44361 40579 44419 40585
rect 44361 40576 44373 40579
rect 40052 40548 44373 40576
rect 44361 40545 44373 40548
rect 44407 40576 44419 40579
rect 44450 40576 44456 40588
rect 44407 40548 44456 40576
rect 44407 40545 44419 40548
rect 44361 40539 44419 40545
rect 44450 40536 44456 40548
rect 44508 40536 44514 40588
rect 44729 40579 44787 40585
rect 44729 40545 44741 40579
rect 44775 40545 44787 40579
rect 44729 40539 44787 40545
rect 30653 40511 30711 40517
rect 30653 40477 30665 40511
rect 30699 40508 30711 40511
rect 31754 40508 31760 40520
rect 30699 40480 31760 40508
rect 30699 40477 30711 40480
rect 30653 40471 30711 40477
rect 31754 40468 31760 40480
rect 31812 40468 31818 40520
rect 32950 40468 32956 40520
rect 33008 40508 33014 40520
rect 33137 40511 33195 40517
rect 33137 40508 33149 40511
rect 33008 40480 33149 40508
rect 33008 40468 33014 40480
rect 33137 40477 33149 40480
rect 33183 40477 33195 40511
rect 33410 40508 33416 40520
rect 33371 40480 33416 40508
rect 33137 40471 33195 40477
rect 33410 40468 33416 40480
rect 33468 40468 33474 40520
rect 38562 40508 38568 40520
rect 38475 40480 38568 40508
rect 38562 40468 38568 40480
rect 38620 40508 38626 40520
rect 38657 40511 38715 40517
rect 38657 40508 38669 40511
rect 38620 40480 38669 40508
rect 38620 40468 38626 40480
rect 38657 40477 38669 40480
rect 38703 40477 38715 40511
rect 38657 40471 38715 40477
rect 39945 40511 40003 40517
rect 39945 40477 39957 40511
rect 39991 40508 40003 40511
rect 41233 40511 41291 40517
rect 41233 40508 41245 40511
rect 39991 40480 41245 40508
rect 39991 40477 40003 40480
rect 39945 40471 40003 40477
rect 41233 40477 41245 40480
rect 41279 40477 41291 40511
rect 41233 40471 41291 40477
rect 44545 40511 44603 40517
rect 44545 40477 44557 40511
rect 44591 40477 44603 40511
rect 44744 40508 44772 40539
rect 44818 40536 44824 40588
rect 44876 40576 44882 40588
rect 45189 40579 45247 40585
rect 45189 40576 45201 40579
rect 44876 40548 45201 40576
rect 44876 40536 44882 40548
rect 45189 40545 45201 40548
rect 45235 40545 45247 40579
rect 45189 40539 45247 40545
rect 45281 40579 45339 40585
rect 45281 40545 45293 40579
rect 45327 40576 45339 40579
rect 46566 40576 46572 40588
rect 45327 40548 46572 40576
rect 45327 40545 45339 40548
rect 45281 40539 45339 40545
rect 46566 40536 46572 40548
rect 46624 40536 46630 40588
rect 50908 40548 51120 40576
rect 44910 40508 44916 40520
rect 44744 40480 44916 40508
rect 44545 40471 44603 40477
rect 30837 40443 30895 40449
rect 30837 40440 30849 40443
rect 26436 40412 30849 40440
rect 9539 40409 9551 40412
rect 9493 40403 9551 40409
rect 30837 40409 30849 40412
rect 30883 40440 30895 40443
rect 40586 40440 40592 40452
rect 30883 40412 33180 40440
rect 30883 40409 30895 40412
rect 30837 40403 30895 40409
rect 9858 40332 9864 40384
rect 9916 40372 9922 40384
rect 10321 40375 10379 40381
rect 10321 40372 10333 40375
rect 9916 40344 10333 40372
rect 9916 40332 9922 40344
rect 10321 40341 10333 40344
rect 10367 40372 10379 40375
rect 12526 40372 12532 40384
rect 10367 40344 12532 40372
rect 10367 40341 10379 40344
rect 10321 40335 10379 40341
rect 12526 40332 12532 40344
rect 12584 40332 12590 40384
rect 21082 40332 21088 40384
rect 21140 40372 21146 40384
rect 21910 40372 21916 40384
rect 21140 40344 21916 40372
rect 21140 40332 21146 40344
rect 21910 40332 21916 40344
rect 21968 40332 21974 40384
rect 23658 40372 23664 40384
rect 23619 40344 23664 40372
rect 23658 40332 23664 40344
rect 23716 40332 23722 40384
rect 24670 40332 24676 40384
rect 24728 40372 24734 40384
rect 28994 40372 29000 40384
rect 24728 40344 29000 40372
rect 24728 40332 24734 40344
rect 28994 40332 29000 40344
rect 29052 40332 29058 40384
rect 29178 40372 29184 40384
rect 29139 40344 29184 40372
rect 29178 40332 29184 40344
rect 29236 40332 29242 40384
rect 32950 40372 32956 40384
rect 32911 40344 32956 40372
rect 32950 40332 32956 40344
rect 33008 40332 33014 40384
rect 33152 40372 33180 40412
rect 34072 40412 40592 40440
rect 34072 40372 34100 40412
rect 40586 40400 40592 40412
rect 40644 40400 40650 40452
rect 41141 40443 41199 40449
rect 41141 40409 41153 40443
rect 41187 40440 41199 40443
rect 44358 40440 44364 40452
rect 41187 40412 44364 40440
rect 41187 40409 41199 40412
rect 41141 40403 41199 40409
rect 44358 40400 44364 40412
rect 44416 40400 44422 40452
rect 34698 40372 34704 40384
rect 33152 40344 34100 40372
rect 34659 40344 34704 40372
rect 34698 40332 34704 40344
rect 34756 40332 34762 40384
rect 40494 40332 40500 40384
rect 40552 40372 40558 40384
rect 41003 40375 41061 40381
rect 41003 40372 41015 40375
rect 40552 40344 41015 40372
rect 40552 40332 40558 40344
rect 41003 40341 41015 40344
rect 41049 40341 41061 40375
rect 41506 40372 41512 40384
rect 41467 40344 41512 40372
rect 41003 40335 41061 40341
rect 41506 40332 41512 40344
rect 41564 40332 41570 40384
rect 41598 40332 41604 40384
rect 41656 40372 41662 40384
rect 44174 40372 44180 40384
rect 41656 40344 44180 40372
rect 41656 40332 41662 40344
rect 44174 40332 44180 40344
rect 44232 40332 44238 40384
rect 44560 40372 44588 40471
rect 44910 40468 44916 40480
rect 44968 40468 44974 40520
rect 45738 40468 45744 40520
rect 45796 40508 45802 40520
rect 46293 40511 46351 40517
rect 46293 40508 46305 40511
rect 45796 40480 46305 40508
rect 45796 40468 45802 40480
rect 46293 40477 46305 40480
rect 46339 40508 46351 40511
rect 48866 40508 48872 40520
rect 46339 40480 48872 40508
rect 46339 40477 46351 40480
rect 46293 40471 46351 40477
rect 48866 40468 48872 40480
rect 48924 40468 48930 40520
rect 44634 40400 44640 40452
rect 44692 40440 44698 40452
rect 50908 40440 50936 40548
rect 51092 40508 51120 40548
rect 52454 40536 52460 40588
rect 52512 40576 52518 40588
rect 52641 40579 52699 40585
rect 52641 40576 52653 40579
rect 52512 40548 52653 40576
rect 52512 40536 52518 40548
rect 52641 40545 52653 40548
rect 52687 40545 52699 40579
rect 52641 40539 52699 40545
rect 52914 40536 52920 40588
rect 52972 40576 52978 40588
rect 58066 40576 58072 40588
rect 52972 40548 58072 40576
rect 52972 40536 52978 40548
rect 58066 40536 58072 40548
rect 58124 40536 58130 40588
rect 58434 40536 58440 40588
rect 58492 40576 58498 40588
rect 58621 40579 58679 40585
rect 58621 40576 58633 40579
rect 58492 40548 58633 40576
rect 58492 40536 58498 40548
rect 58621 40545 58633 40548
rect 58667 40545 58679 40579
rect 58621 40539 58679 40545
rect 59170 40536 59176 40588
rect 59228 40576 59234 40588
rect 59722 40576 59728 40588
rect 59228 40548 59728 40576
rect 59228 40536 59234 40548
rect 59722 40536 59728 40548
rect 59780 40576 59786 40588
rect 60185 40579 60243 40585
rect 60185 40576 60197 40579
rect 59780 40548 60197 40576
rect 59780 40536 59786 40548
rect 60185 40545 60197 40548
rect 60231 40545 60243 40579
rect 60185 40539 60243 40545
rect 66073 40579 66131 40585
rect 66073 40545 66085 40579
rect 66119 40576 66131 40579
rect 67082 40576 67088 40588
rect 66119 40548 67088 40576
rect 66119 40545 66131 40548
rect 66073 40539 66131 40545
rect 67082 40536 67088 40548
rect 67140 40536 67146 40588
rect 77389 40579 77447 40585
rect 77389 40545 77401 40579
rect 77435 40545 77447 40579
rect 77389 40539 77447 40545
rect 52822 40508 52828 40520
rect 51092 40480 52828 40508
rect 52822 40468 52828 40480
rect 52880 40468 52886 40520
rect 53006 40508 53012 40520
rect 52967 40480 53012 40508
rect 53006 40468 53012 40480
rect 53064 40468 53070 40520
rect 53098 40468 53104 40520
rect 53156 40508 53162 40520
rect 65334 40508 65340 40520
rect 53156 40480 65340 40508
rect 53156 40468 53162 40480
rect 65334 40468 65340 40480
rect 65392 40468 65398 40520
rect 65613 40511 65671 40517
rect 65613 40477 65625 40511
rect 65659 40508 65671 40511
rect 65797 40511 65855 40517
rect 65797 40508 65809 40511
rect 65659 40480 65809 40508
rect 65659 40477 65671 40480
rect 65613 40471 65671 40477
rect 65797 40477 65809 40480
rect 65843 40508 65855 40511
rect 65843 40480 66760 40508
rect 65843 40477 65855 40480
rect 65797 40471 65855 40477
rect 52917 40443 52975 40449
rect 52917 40440 52929 40443
rect 44692 40412 50936 40440
rect 52012 40412 52929 40440
rect 44692 40400 44698 40412
rect 45554 40372 45560 40384
rect 44560 40344 45560 40372
rect 45554 40332 45560 40344
rect 45612 40332 45618 40384
rect 45738 40372 45744 40384
rect 45699 40344 45744 40372
rect 45738 40332 45744 40344
rect 45796 40332 45802 40384
rect 46014 40372 46020 40384
rect 45975 40344 46020 40372
rect 46014 40332 46020 40344
rect 46072 40332 46078 40384
rect 46477 40375 46535 40381
rect 46477 40341 46489 40375
rect 46523 40372 46535 40375
rect 46566 40372 46572 40384
rect 46523 40344 46572 40372
rect 46523 40341 46535 40344
rect 46477 40335 46535 40341
rect 46566 40332 46572 40344
rect 46624 40332 46630 40384
rect 49510 40332 49516 40384
rect 49568 40372 49574 40384
rect 52012 40372 52040 40412
rect 52917 40409 52929 40412
rect 52963 40409 52975 40443
rect 54294 40440 54300 40452
rect 52917 40403 52975 40409
rect 53208 40412 54300 40440
rect 49568 40344 52040 40372
rect 52806 40375 52864 40381
rect 49568 40332 49574 40344
rect 52806 40341 52818 40375
rect 52852 40372 52864 40375
rect 53208 40372 53236 40412
rect 54294 40400 54300 40412
rect 54352 40400 54358 40452
rect 63126 40400 63132 40452
rect 63184 40440 63190 40452
rect 65628 40440 65656 40471
rect 63184 40412 65656 40440
rect 66732 40440 66760 40480
rect 66806 40468 66812 40520
rect 66864 40508 66870 40520
rect 67177 40511 67235 40517
rect 67177 40508 67189 40511
rect 66864 40480 67189 40508
rect 66864 40468 66870 40480
rect 67177 40477 67189 40480
rect 67223 40477 67235 40511
rect 67177 40471 67235 40477
rect 67450 40468 67456 40520
rect 67508 40508 67514 40520
rect 71961 40511 72019 40517
rect 71961 40508 71973 40511
rect 67508 40480 71973 40508
rect 67508 40468 67514 40480
rect 71961 40477 71973 40480
rect 72007 40508 72019 40511
rect 72145 40511 72203 40517
rect 72145 40508 72157 40511
rect 72007 40480 72157 40508
rect 72007 40477 72019 40480
rect 71961 40471 72019 40477
rect 72145 40477 72157 40480
rect 72191 40477 72203 40511
rect 72418 40508 72424 40520
rect 72379 40480 72424 40508
rect 72145 40471 72203 40477
rect 72418 40468 72424 40480
rect 72476 40468 72482 40520
rect 72602 40468 72608 40520
rect 72660 40508 72666 40520
rect 77202 40508 77208 40520
rect 72660 40480 77208 40508
rect 72660 40468 72666 40480
rect 77202 40468 77208 40480
rect 77260 40508 77266 40520
rect 77404 40508 77432 40539
rect 77478 40536 77484 40588
rect 77536 40576 77542 40588
rect 77573 40579 77631 40585
rect 77573 40576 77585 40579
rect 77536 40548 77585 40576
rect 77536 40536 77542 40548
rect 77573 40545 77585 40548
rect 77619 40545 77631 40579
rect 83550 40576 83556 40588
rect 83511 40548 83556 40576
rect 77573 40539 77631 40545
rect 83550 40536 83556 40548
rect 83608 40536 83614 40588
rect 83734 40576 83740 40588
rect 83695 40548 83740 40576
rect 83734 40536 83740 40548
rect 83792 40576 83798 40588
rect 83829 40579 83887 40585
rect 83829 40576 83841 40579
rect 83792 40548 83841 40576
rect 83792 40536 83798 40548
rect 83829 40545 83841 40548
rect 83875 40545 83887 40579
rect 84562 40576 84568 40588
rect 84523 40548 84568 40576
rect 83829 40539 83887 40545
rect 84562 40536 84568 40548
rect 84620 40536 84626 40588
rect 83274 40508 83280 40520
rect 77260 40480 77432 40508
rect 83235 40480 83280 40508
rect 77260 40468 77266 40480
rect 83274 40468 83280 40480
rect 83332 40468 83338 40520
rect 67468 40440 67496 40468
rect 66732 40412 67496 40440
rect 63184 40400 63190 40412
rect 52852 40344 53236 40372
rect 53285 40375 53343 40381
rect 52852 40341 52864 40344
rect 52806 40335 52864 40341
rect 53285 40341 53297 40375
rect 53331 40372 53343 40375
rect 53926 40372 53932 40384
rect 53331 40344 53932 40372
rect 53331 40341 53343 40344
rect 53285 40335 53343 40341
rect 53926 40332 53932 40344
rect 53984 40332 53990 40384
rect 58710 40332 58716 40384
rect 58768 40372 58774 40384
rect 61010 40372 61016 40384
rect 58768 40344 61016 40372
rect 58768 40332 58774 40344
rect 61010 40332 61016 40344
rect 61068 40372 61074 40384
rect 61746 40372 61752 40384
rect 61068 40344 61752 40372
rect 61068 40332 61074 40344
rect 61746 40332 61752 40344
rect 61804 40332 61810 40384
rect 73522 40372 73528 40384
rect 73483 40344 73528 40372
rect 73522 40332 73528 40344
rect 73580 40332 73586 40384
rect 1104 40282 108008 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 65686 40282
rect 65738 40230 65750 40282
rect 65802 40230 65814 40282
rect 65866 40230 65878 40282
rect 65930 40230 96406 40282
rect 96458 40230 96470 40282
rect 96522 40230 96534 40282
rect 96586 40230 96598 40282
rect 96650 40230 108008 40282
rect 1104 40208 108008 40230
rect 3878 40128 3884 40180
rect 3936 40168 3942 40180
rect 10137 40171 10195 40177
rect 3936 40140 10088 40168
rect 3936 40128 3942 40140
rect 4798 40060 4804 40112
rect 4856 40100 4862 40112
rect 4982 40100 4988 40112
rect 4856 40072 4988 40100
rect 4856 40060 4862 40072
rect 4982 40060 4988 40072
rect 5040 40060 5046 40112
rect 10060 40032 10088 40140
rect 10137 40137 10149 40171
rect 10183 40168 10195 40171
rect 10226 40168 10232 40180
rect 10183 40140 10232 40168
rect 10183 40137 10195 40140
rect 10137 40131 10195 40137
rect 10226 40128 10232 40140
rect 10284 40128 10290 40180
rect 27338 40168 27344 40180
rect 12452 40140 27344 40168
rect 12452 40032 12480 40140
rect 27338 40128 27344 40140
rect 27396 40128 27402 40180
rect 27522 40128 27528 40180
rect 27580 40168 27586 40180
rect 27706 40168 27712 40180
rect 27580 40140 27712 40168
rect 27580 40128 27586 40140
rect 27706 40128 27712 40140
rect 27764 40128 27770 40180
rect 29454 40168 29460 40180
rect 29415 40140 29460 40168
rect 29454 40128 29460 40140
rect 29512 40128 29518 40180
rect 34698 40128 34704 40180
rect 34756 40168 34762 40180
rect 57790 40168 57796 40180
rect 34756 40140 57796 40168
rect 34756 40128 34762 40140
rect 57790 40128 57796 40140
rect 57848 40128 57854 40180
rect 58802 40168 58808 40180
rect 58763 40140 58808 40168
rect 58802 40128 58808 40140
rect 58860 40128 58866 40180
rect 72418 40128 72424 40180
rect 72476 40168 72482 40180
rect 72697 40171 72755 40177
rect 72697 40168 72709 40171
rect 72476 40140 72709 40168
rect 72476 40128 72482 40140
rect 72697 40137 72709 40140
rect 72743 40137 72755 40171
rect 74258 40168 74264 40180
rect 74219 40140 74264 40168
rect 72697 40131 72755 40137
rect 74258 40128 74264 40140
rect 74316 40128 74322 40180
rect 83734 40168 83740 40180
rect 83695 40140 83740 40168
rect 83734 40128 83740 40140
rect 83792 40128 83798 40180
rect 12526 40060 12532 40112
rect 12584 40100 12590 40112
rect 38562 40100 38568 40112
rect 12584 40072 38568 40100
rect 12584 40060 12590 40072
rect 38562 40060 38568 40072
rect 38620 40100 38626 40112
rect 40494 40100 40500 40112
rect 38620 40072 40500 40100
rect 38620 40060 38626 40072
rect 40494 40060 40500 40072
rect 40552 40060 40558 40112
rect 40773 40103 40831 40109
rect 40773 40069 40785 40103
rect 40819 40100 40831 40103
rect 45738 40100 45744 40112
rect 40819 40072 45744 40100
rect 40819 40069 40831 40072
rect 40773 40063 40831 40069
rect 45738 40060 45744 40072
rect 45796 40060 45802 40112
rect 48130 40100 48136 40112
rect 47412 40072 48136 40100
rect 16117 40035 16175 40041
rect 16117 40032 16129 40035
rect 10060 40004 12480 40032
rect 15672 40004 16129 40032
rect 4798 39924 4804 39976
rect 4856 39964 4862 39976
rect 8757 39967 8815 39973
rect 8757 39964 8769 39967
rect 4856 39936 8769 39964
rect 4856 39924 4862 39936
rect 8757 39933 8769 39936
rect 8803 39933 8815 39967
rect 8757 39927 8815 39933
rect 9033 39967 9091 39973
rect 9033 39933 9045 39967
rect 9079 39964 9091 39967
rect 9398 39964 9404 39976
rect 9079 39936 9404 39964
rect 9079 39933 9091 39936
rect 9033 39927 9091 39933
rect 9398 39924 9404 39936
rect 9456 39924 9462 39976
rect 15672 39973 15700 40004
rect 16117 40001 16129 40004
rect 16163 40032 16175 40035
rect 17126 40032 17132 40044
rect 16163 40004 17132 40032
rect 16163 40001 16175 40004
rect 16117 39995 16175 40001
rect 17126 39992 17132 40004
rect 17184 39992 17190 40044
rect 18414 40032 18420 40044
rect 18064 40004 18420 40032
rect 15657 39967 15715 39973
rect 15657 39933 15669 39967
rect 15703 39933 15715 39967
rect 15657 39927 15715 39933
rect 16853 39967 16911 39973
rect 16853 39933 16865 39967
rect 16899 39964 16911 39967
rect 17310 39964 17316 39976
rect 16899 39936 17316 39964
rect 16899 39933 16911 39936
rect 16853 39927 16911 39933
rect 17310 39924 17316 39936
rect 17368 39924 17374 39976
rect 18064 39973 18092 40004
rect 18414 39992 18420 40004
rect 18472 39992 18478 40044
rect 40678 40041 40684 40044
rect 40644 40035 40684 40041
rect 40644 40001 40656 40035
rect 40644 39995 40684 40001
rect 40678 39992 40684 39995
rect 40736 39992 40742 40044
rect 40865 40035 40923 40041
rect 40865 40001 40877 40035
rect 40911 40001 40923 40035
rect 40865 39995 40923 40001
rect 18049 39967 18107 39973
rect 18049 39933 18061 39967
rect 18095 39933 18107 39967
rect 23658 39964 23664 39976
rect 23619 39936 23664 39964
rect 18049 39927 18107 39933
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 28442 39924 28448 39976
rect 28500 39964 28506 39976
rect 29273 39967 29331 39973
rect 29273 39964 29285 39967
rect 28500 39936 29285 39964
rect 28500 39924 28506 39936
rect 29273 39933 29285 39936
rect 29319 39964 29331 39967
rect 29454 39964 29460 39976
rect 29319 39936 29460 39964
rect 29319 39933 29331 39936
rect 29273 39927 29331 39933
rect 29454 39924 29460 39936
rect 29512 39924 29518 39976
rect 40310 39964 40316 39976
rect 29656 39936 40316 39964
rect 15562 39856 15568 39908
rect 15620 39896 15626 39908
rect 18141 39899 18199 39905
rect 18141 39896 18153 39899
rect 15620 39868 18153 39896
rect 15620 39856 15626 39868
rect 18141 39865 18153 39868
rect 18187 39865 18199 39899
rect 18141 39859 18199 39865
rect 22738 39856 22744 39908
rect 22796 39896 22802 39908
rect 23753 39899 23811 39905
rect 23753 39896 23765 39899
rect 22796 39868 23765 39896
rect 22796 39856 22802 39868
rect 23753 39865 23765 39868
rect 23799 39896 23811 39899
rect 29656 39896 29684 39936
rect 40310 39924 40316 39936
rect 40368 39924 40374 39976
rect 40402 39924 40408 39976
rect 40460 39964 40466 39976
rect 40460 39936 40724 39964
rect 40460 39924 40466 39936
rect 23799 39868 29684 39896
rect 23799 39865 23811 39868
rect 23753 39859 23811 39865
rect 38930 39856 38936 39908
rect 38988 39896 38994 39908
rect 40497 39899 40555 39905
rect 40497 39896 40509 39899
rect 38988 39868 40509 39896
rect 38988 39856 38994 39868
rect 40497 39865 40509 39868
rect 40543 39865 40555 39899
rect 40696 39896 40724 39936
rect 40880 39896 40908 39995
rect 40954 39992 40960 40044
rect 41012 40032 41018 40044
rect 41690 40032 41696 40044
rect 41012 40004 41696 40032
rect 41012 39992 41018 40004
rect 41690 39992 41696 40004
rect 41748 39992 41754 40044
rect 44450 39992 44456 40044
rect 44508 40032 44514 40044
rect 44910 40032 44916 40044
rect 44508 40004 44916 40032
rect 44508 39992 44514 40004
rect 44910 39992 44916 40004
rect 44968 40032 44974 40044
rect 46014 40032 46020 40044
rect 44968 40004 46020 40032
rect 44968 39992 44974 40004
rect 46014 39992 46020 40004
rect 46072 39992 46078 40044
rect 46842 39924 46848 39976
rect 46900 39964 46906 39976
rect 47412 39973 47440 40072
rect 48130 40060 48136 40072
rect 48188 40100 48194 40112
rect 48685 40103 48743 40109
rect 48685 40100 48697 40103
rect 48188 40072 48697 40100
rect 48188 40060 48194 40072
rect 48685 40069 48697 40072
rect 48731 40069 48743 40103
rect 48685 40063 48743 40069
rect 48774 40060 48780 40112
rect 48832 40100 48838 40112
rect 53098 40100 53104 40112
rect 48832 40072 53104 40100
rect 48832 40060 48838 40072
rect 53098 40060 53104 40072
rect 53156 40060 53162 40112
rect 54110 40109 54116 40112
rect 54094 40103 54116 40109
rect 54094 40069 54106 40103
rect 54094 40063 54116 40069
rect 54110 40060 54116 40063
rect 54168 40060 54174 40112
rect 54386 40060 54392 40112
rect 54444 40100 54450 40112
rect 54444 40072 54800 40100
rect 54444 40060 54450 40072
rect 48501 40035 48559 40041
rect 48501 40001 48513 40035
rect 48547 40032 48559 40035
rect 52454 40032 52460 40044
rect 48547 40004 52460 40032
rect 48547 40001 48559 40004
rect 48501 39995 48559 40001
rect 52454 39992 52460 40004
rect 52512 39992 52518 40044
rect 54297 40035 54355 40041
rect 54297 40001 54309 40035
rect 54343 40032 54355 40035
rect 54662 40032 54668 40044
rect 54343 40004 54668 40032
rect 54343 40001 54355 40004
rect 54297 39995 54355 40001
rect 54662 39992 54668 40004
rect 54720 39992 54726 40044
rect 54772 40032 54800 40072
rect 54846 40060 54852 40112
rect 54904 40100 54910 40112
rect 54904 40072 54949 40100
rect 54904 40060 54910 40072
rect 59538 40060 59544 40112
rect 59596 40100 59602 40112
rect 82725 40103 82783 40109
rect 59596 40072 60136 40100
rect 59596 40060 59602 40072
rect 58621 40035 58679 40041
rect 58621 40032 58633 40035
rect 54772 40004 58633 40032
rect 58621 40001 58633 40004
rect 58667 40032 58679 40035
rect 60108 40032 60136 40072
rect 82725 40069 82737 40103
rect 82771 40100 82783 40103
rect 83274 40100 83280 40112
rect 82771 40072 83280 40100
rect 82771 40069 82783 40072
rect 82725 40063 82783 40069
rect 83274 40060 83280 40072
rect 83332 40060 83338 40112
rect 58667 40004 59308 40032
rect 60108 40004 72740 40032
rect 58667 40001 58679 40004
rect 58621 39995 58679 40001
rect 47213 39967 47271 39973
rect 47213 39964 47225 39967
rect 46900 39936 47225 39964
rect 46900 39924 46906 39936
rect 47213 39933 47225 39936
rect 47259 39933 47271 39967
rect 47213 39927 47271 39933
rect 47397 39967 47455 39973
rect 47397 39933 47409 39967
rect 47443 39933 47455 39967
rect 47397 39927 47455 39933
rect 47857 39967 47915 39973
rect 47857 39933 47869 39967
rect 47903 39933 47915 39967
rect 47857 39927 47915 39933
rect 47949 39967 48007 39973
rect 47949 39933 47961 39967
rect 47995 39933 48007 39967
rect 47949 39927 48007 39933
rect 40696 39868 40908 39896
rect 40497 39859 40555 39865
rect 44266 39856 44272 39908
rect 44324 39896 44330 39908
rect 47029 39899 47087 39905
rect 47029 39896 47041 39899
rect 44324 39868 47041 39896
rect 44324 39856 44330 39868
rect 47029 39865 47041 39868
rect 47075 39896 47087 39899
rect 47872 39896 47900 39927
rect 47075 39868 47900 39896
rect 47964 39896 47992 39927
rect 51074 39924 51080 39976
rect 51132 39964 51138 39976
rect 53374 39964 53380 39976
rect 51132 39936 53380 39964
rect 51132 39924 51138 39936
rect 53374 39924 53380 39936
rect 53432 39924 53438 39976
rect 53926 39964 53932 39976
rect 53887 39936 53932 39964
rect 53926 39924 53932 39936
rect 53984 39924 53990 39976
rect 54202 39973 54208 39976
rect 54159 39967 54208 39973
rect 54159 39933 54171 39967
rect 54205 39933 54208 39967
rect 54159 39927 54208 39933
rect 54202 39924 54208 39927
rect 54260 39924 54266 39976
rect 57790 39924 57796 39976
rect 57848 39964 57854 39976
rect 57977 39967 58035 39973
rect 57977 39964 57989 39967
rect 57848 39936 57989 39964
rect 57848 39924 57854 39936
rect 57977 39933 57989 39936
rect 58023 39933 58035 39967
rect 57977 39927 58035 39933
rect 58066 39924 58072 39976
rect 58124 39964 58130 39976
rect 58124 39936 58169 39964
rect 58124 39924 58130 39936
rect 58802 39924 58808 39976
rect 58860 39964 58866 39976
rect 58989 39967 59047 39973
rect 58989 39964 59001 39967
rect 58860 39936 59001 39964
rect 58860 39924 58866 39936
rect 58989 39933 59001 39936
rect 59035 39933 59047 39967
rect 59170 39964 59176 39976
rect 59131 39936 59176 39964
rect 58989 39927 59047 39933
rect 59170 39924 59176 39936
rect 59228 39924 59234 39976
rect 59280 39964 59308 40004
rect 59633 39967 59691 39973
rect 59633 39964 59645 39967
rect 59280 39936 59645 39964
rect 59633 39933 59645 39936
rect 59679 39933 59691 39967
rect 59633 39927 59691 39933
rect 59725 39967 59783 39973
rect 59725 39933 59737 39967
rect 59771 39933 59783 39967
rect 59725 39927 59783 39933
rect 48222 39896 48228 39908
rect 47964 39868 48228 39896
rect 47075 39865 47087 39868
rect 47029 39859 47087 39865
rect 48222 39856 48228 39868
rect 48280 39896 48286 39908
rect 48869 39899 48927 39905
rect 48869 39896 48881 39899
rect 48280 39868 48881 39896
rect 48280 39856 48286 39868
rect 48869 39865 48881 39868
rect 48915 39865 48927 39899
rect 48869 39859 48927 39865
rect 49050 39856 49056 39908
rect 49108 39896 49114 39908
rect 54386 39896 54392 39908
rect 49108 39868 54392 39896
rect 49108 39856 49114 39868
rect 54386 39856 54392 39868
rect 54444 39856 54450 39908
rect 59538 39896 59544 39908
rect 54496 39868 59544 39896
rect 10594 39828 10600 39840
rect 10555 39800 10600 39828
rect 10594 39788 10600 39800
rect 10652 39788 10658 39840
rect 15102 39788 15108 39840
rect 15160 39828 15166 39840
rect 15841 39831 15899 39837
rect 15841 39828 15853 39831
rect 15160 39800 15853 39828
rect 15160 39788 15166 39800
rect 15841 39797 15853 39800
rect 15887 39797 15899 39831
rect 15841 39791 15899 39797
rect 16574 39788 16580 39840
rect 16632 39828 16638 39840
rect 17037 39831 17095 39837
rect 17037 39828 17049 39831
rect 16632 39800 17049 39828
rect 16632 39788 16638 39800
rect 17037 39797 17049 39800
rect 17083 39797 17095 39831
rect 17310 39828 17316 39840
rect 17271 39800 17316 39828
rect 17037 39791 17095 39797
rect 17310 39788 17316 39800
rect 17368 39788 17374 39840
rect 19334 39788 19340 39840
rect 19392 39828 19398 39840
rect 24118 39828 24124 39840
rect 19392 39800 24124 39828
rect 19392 39788 19398 39800
rect 24118 39788 24124 39800
rect 24176 39788 24182 39840
rect 29454 39788 29460 39840
rect 29512 39828 29518 39840
rect 29733 39831 29791 39837
rect 29733 39828 29745 39831
rect 29512 39800 29745 39828
rect 29512 39788 29518 39800
rect 29733 39797 29745 39800
rect 29779 39828 29791 39831
rect 32398 39828 32404 39840
rect 29779 39800 32404 39828
rect 29779 39797 29791 39800
rect 29733 39791 29791 39797
rect 32398 39788 32404 39800
rect 32456 39788 32462 39840
rect 40862 39788 40868 39840
rect 40920 39828 40926 39840
rect 41141 39831 41199 39837
rect 41141 39828 41153 39831
rect 40920 39800 41153 39828
rect 40920 39788 40926 39800
rect 41141 39797 41153 39800
rect 41187 39797 41199 39831
rect 46842 39828 46848 39840
rect 46803 39800 46848 39828
rect 41141 39791 41199 39797
rect 46842 39788 46848 39800
rect 46900 39788 46906 39840
rect 46934 39788 46940 39840
rect 46992 39828 46998 39840
rect 54496 39828 54524 39868
rect 59538 39856 59544 39868
rect 59596 39856 59602 39908
rect 46992 39800 54524 39828
rect 54573 39831 54631 39837
rect 46992 39788 46998 39800
rect 54573 39797 54585 39831
rect 54619 39828 54631 39831
rect 56502 39828 56508 39840
rect 54619 39800 56508 39828
rect 54619 39797 54631 39800
rect 54573 39791 54631 39797
rect 56502 39788 56508 39800
rect 56560 39788 56566 39840
rect 57790 39788 57796 39840
rect 57848 39828 57854 39840
rect 59446 39828 59452 39840
rect 57848 39800 59452 39828
rect 57848 39788 57854 39800
rect 59446 39788 59452 39800
rect 59504 39788 59510 39840
rect 59740 39828 59768 39927
rect 60550 39924 60556 39976
rect 60608 39964 60614 39976
rect 71130 39964 71136 39976
rect 60608 39936 71136 39964
rect 60608 39924 60614 39936
rect 71130 39924 71136 39936
rect 71188 39924 71194 39976
rect 71225 39967 71283 39973
rect 71225 39933 71237 39967
rect 71271 39964 71283 39967
rect 72142 39964 72148 39976
rect 71271 39936 72148 39964
rect 71271 39933 71283 39936
rect 71225 39927 71283 39933
rect 72142 39924 72148 39936
rect 72200 39924 72206 39976
rect 72329 39967 72387 39973
rect 72329 39933 72341 39967
rect 72375 39933 72387 39967
rect 72510 39964 72516 39976
rect 72471 39936 72516 39964
rect 72329 39927 72387 39933
rect 60277 39899 60335 39905
rect 60277 39865 60289 39899
rect 60323 39896 60335 39899
rect 60826 39896 60832 39908
rect 60323 39868 60832 39896
rect 60323 39865 60335 39868
rect 60277 39859 60335 39865
rect 60826 39856 60832 39868
rect 60884 39856 60890 39908
rect 65150 39856 65156 39908
rect 65208 39896 65214 39908
rect 66070 39896 66076 39908
rect 65208 39868 66076 39896
rect 65208 39856 65214 39868
rect 66070 39856 66076 39868
rect 66128 39856 66134 39908
rect 67634 39856 67640 39908
rect 67692 39896 67698 39908
rect 72344 39896 72372 39927
rect 72510 39924 72516 39936
rect 72568 39924 72574 39976
rect 67692 39868 72372 39896
rect 67692 39856 67698 39868
rect 59998 39828 60004 39840
rect 59740 39800 60004 39828
rect 59998 39788 60004 39800
rect 60056 39828 60062 39840
rect 60553 39831 60611 39837
rect 60553 39828 60565 39831
rect 60056 39800 60565 39828
rect 60056 39788 60062 39800
rect 60553 39797 60565 39800
rect 60599 39828 60611 39831
rect 67358 39828 67364 39840
rect 60599 39800 67364 39828
rect 60599 39797 60611 39800
rect 60553 39791 60611 39797
rect 67358 39788 67364 39800
rect 67416 39788 67422 39840
rect 71317 39831 71375 39837
rect 71317 39797 71329 39831
rect 71363 39828 71375 39831
rect 71682 39828 71688 39840
rect 71363 39800 71688 39828
rect 71363 39797 71375 39800
rect 71317 39791 71375 39797
rect 71682 39788 71688 39800
rect 71740 39788 71746 39840
rect 72344 39828 72372 39868
rect 72421 39899 72479 39905
rect 72421 39865 72433 39899
rect 72467 39896 72479 39899
rect 72602 39896 72608 39908
rect 72467 39868 72608 39896
rect 72467 39865 72479 39868
rect 72421 39859 72479 39865
rect 72602 39856 72608 39868
rect 72660 39856 72666 39908
rect 72712 39896 72740 40004
rect 79686 39992 79692 40044
rect 79744 40032 79750 40044
rect 83369 40035 83427 40041
rect 83369 40032 83381 40035
rect 79744 40004 83381 40032
rect 79744 39992 79750 40004
rect 83369 40001 83381 40004
rect 83415 40032 83427 40035
rect 83550 40032 83556 40044
rect 83415 40004 83556 40032
rect 83415 40001 83427 40004
rect 83369 39995 83427 40001
rect 83550 39992 83556 40004
rect 83608 39992 83614 40044
rect 73522 39924 73528 39976
rect 73580 39964 73586 39976
rect 74169 39967 74227 39973
rect 74169 39964 74181 39967
rect 73580 39936 74181 39964
rect 73580 39924 73586 39936
rect 74169 39933 74181 39936
rect 74215 39933 74227 39967
rect 74169 39927 74227 39933
rect 77202 39924 77208 39976
rect 77260 39964 77266 39976
rect 77389 39967 77447 39973
rect 77389 39964 77401 39967
rect 77260 39936 77401 39964
rect 77260 39924 77266 39936
rect 77389 39933 77401 39936
rect 77435 39933 77447 39967
rect 77389 39927 77447 39933
rect 82170 39924 82176 39976
rect 82228 39964 82234 39976
rect 82449 39967 82507 39973
rect 82449 39964 82461 39967
rect 82228 39936 82461 39964
rect 82228 39924 82234 39936
rect 82262 39896 82268 39908
rect 72712 39868 82268 39896
rect 82262 39856 82268 39868
rect 82320 39856 82326 39908
rect 82372 39840 82400 39936
rect 82449 39933 82461 39936
rect 82495 39933 82507 39967
rect 82449 39927 82507 39933
rect 83185 39967 83243 39973
rect 83185 39933 83197 39967
rect 83231 39964 83243 39967
rect 83734 39964 83740 39976
rect 83231 39936 83740 39964
rect 83231 39933 83243 39936
rect 83185 39927 83243 39933
rect 83734 39924 83740 39936
rect 83792 39924 83798 39976
rect 73157 39831 73215 39837
rect 73157 39828 73169 39831
rect 72344 39800 73169 39828
rect 73157 39797 73169 39800
rect 73203 39828 73215 39831
rect 77570 39828 77576 39840
rect 73203 39800 77576 39828
rect 73203 39797 73215 39800
rect 73157 39791 73215 39797
rect 77570 39788 77576 39800
rect 77628 39828 77634 39840
rect 77754 39828 77760 39840
rect 77628 39800 77760 39828
rect 77628 39788 77634 39800
rect 77754 39788 77760 39800
rect 77812 39788 77818 39840
rect 82354 39828 82360 39840
rect 82315 39800 82360 39828
rect 82354 39788 82360 39800
rect 82412 39788 82418 39840
rect 1104 39738 108008 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 81046 39738
rect 81098 39686 81110 39738
rect 81162 39686 81174 39738
rect 81226 39686 81238 39738
rect 81290 39686 108008 39738
rect 1104 39664 108008 39686
rect 3786 39584 3792 39636
rect 3844 39624 3850 39636
rect 12066 39624 12072 39636
rect 3844 39596 12072 39624
rect 3844 39584 3850 39596
rect 12066 39584 12072 39596
rect 12124 39584 12130 39636
rect 22370 39624 22376 39636
rect 22331 39596 22376 39624
rect 22370 39584 22376 39596
rect 22428 39584 22434 39636
rect 22738 39624 22744 39636
rect 22699 39596 22744 39624
rect 22738 39584 22744 39596
rect 22796 39584 22802 39636
rect 24118 39584 24124 39636
rect 24176 39624 24182 39636
rect 38010 39624 38016 39636
rect 24176 39596 38016 39624
rect 24176 39584 24182 39596
rect 38010 39584 38016 39596
rect 38068 39624 38074 39636
rect 44266 39624 44272 39636
rect 38068 39596 44272 39624
rect 38068 39584 38074 39596
rect 44266 39584 44272 39596
rect 44324 39584 44330 39636
rect 44358 39584 44364 39636
rect 44416 39624 44422 39636
rect 45465 39627 45523 39633
rect 45465 39624 45477 39627
rect 44416 39596 45477 39624
rect 44416 39584 44422 39596
rect 45465 39593 45477 39596
rect 45511 39593 45523 39627
rect 45465 39587 45523 39593
rect 45833 39627 45891 39633
rect 45833 39593 45845 39627
rect 45879 39624 45891 39627
rect 46014 39624 46020 39636
rect 45879 39596 46020 39624
rect 45879 39593 45891 39596
rect 45833 39587 45891 39593
rect 46014 39584 46020 39596
rect 46072 39624 46078 39636
rect 46934 39624 46940 39636
rect 46072 39596 46940 39624
rect 46072 39584 46078 39596
rect 46934 39584 46940 39596
rect 46992 39584 46998 39636
rect 48038 39624 48044 39636
rect 47228 39596 48044 39624
rect 22756 39556 22784 39584
rect 32861 39559 32919 39565
rect 32861 39556 32873 39559
rect 21836 39528 22784 39556
rect 29748 39528 32873 39556
rect 4525 39491 4583 39497
rect 4525 39457 4537 39491
rect 4571 39488 4583 39491
rect 4614 39488 4620 39500
rect 4571 39460 4620 39488
rect 4571 39457 4583 39460
rect 4525 39451 4583 39457
rect 4614 39448 4620 39460
rect 4672 39448 4678 39500
rect 9122 39448 9128 39500
rect 9180 39488 9186 39500
rect 16117 39491 16175 39497
rect 9180 39460 14504 39488
rect 9180 39448 9186 39460
rect 4617 39287 4675 39293
rect 4617 39253 4629 39287
rect 4663 39284 4675 39287
rect 4706 39284 4712 39296
rect 4663 39256 4712 39284
rect 4663 39253 4675 39256
rect 4617 39247 4675 39253
rect 4706 39244 4712 39256
rect 4764 39284 4770 39296
rect 9122 39284 9128 39296
rect 4764 39256 9128 39284
rect 4764 39244 4770 39256
rect 9122 39244 9128 39256
rect 9180 39244 9186 39296
rect 14476 39284 14504 39460
rect 16117 39457 16129 39491
rect 16163 39488 16175 39491
rect 17957 39491 18015 39497
rect 17957 39488 17969 39491
rect 16163 39460 17969 39488
rect 16163 39457 16175 39460
rect 16117 39451 16175 39457
rect 17957 39457 17969 39460
rect 18003 39488 18015 39491
rect 21082 39488 21088 39500
rect 18003 39460 21088 39488
rect 18003 39457 18015 39460
rect 17957 39451 18015 39457
rect 21082 39448 21088 39460
rect 21140 39448 21146 39500
rect 21358 39488 21364 39500
rect 21319 39460 21364 39488
rect 21358 39448 21364 39460
rect 21416 39448 21422 39500
rect 21836 39497 21864 39528
rect 21821 39491 21879 39497
rect 21821 39457 21833 39491
rect 21867 39457 21879 39491
rect 21821 39451 21879 39457
rect 21913 39491 21971 39497
rect 21913 39457 21925 39491
rect 21959 39488 21971 39491
rect 21959 39460 22324 39488
rect 21959 39457 21971 39460
rect 21913 39451 21971 39457
rect 16390 39420 16396 39432
rect 16351 39392 16396 39420
rect 16390 39380 16396 39392
rect 16448 39380 16454 39432
rect 17773 39423 17831 39429
rect 17773 39389 17785 39423
rect 17819 39420 17831 39423
rect 17862 39420 17868 39432
rect 17819 39392 17868 39420
rect 17819 39389 17831 39392
rect 17773 39383 17831 39389
rect 17862 39380 17868 39392
rect 17920 39380 17926 39432
rect 21177 39423 21235 39429
rect 21177 39420 21189 39423
rect 21008 39392 21189 39420
rect 19242 39284 19248 39296
rect 14476 39256 19248 39284
rect 19242 39244 19248 39256
rect 19300 39244 19306 39296
rect 20714 39244 20720 39296
rect 20772 39284 20778 39296
rect 21008 39293 21036 39392
rect 21177 39389 21189 39392
rect 21223 39389 21235 39423
rect 21177 39383 21235 39389
rect 21358 39312 21364 39364
rect 21416 39352 21422 39364
rect 22296 39352 22324 39460
rect 27890 39448 27896 39500
rect 27948 39488 27954 39500
rect 29748 39497 29776 39528
rect 32861 39525 32873 39528
rect 32907 39556 32919 39559
rect 32950 39556 32956 39568
rect 32907 39528 32956 39556
rect 32907 39525 32919 39528
rect 32861 39519 32919 39525
rect 32950 39516 32956 39528
rect 33008 39556 33014 39568
rect 33008 39528 33088 39556
rect 33008 39516 33014 39528
rect 33060 39497 33088 39528
rect 44818 39516 44824 39568
rect 44876 39556 44882 39568
rect 46293 39559 46351 39565
rect 46293 39556 46305 39559
rect 44876 39528 46305 39556
rect 44876 39516 44882 39528
rect 46293 39525 46305 39528
rect 46339 39556 46351 39559
rect 46339 39528 46520 39556
rect 46339 39525 46351 39528
rect 46293 39519 46351 39525
rect 27985 39491 28043 39497
rect 27985 39488 27997 39491
rect 27948 39460 27997 39488
rect 27948 39448 27954 39460
rect 27985 39457 27997 39460
rect 28031 39488 28043 39491
rect 29733 39491 29791 39497
rect 29733 39488 29745 39491
rect 28031 39460 29745 39488
rect 28031 39457 28043 39460
rect 27985 39451 28043 39457
rect 29733 39457 29745 39460
rect 29779 39457 29791 39491
rect 29733 39451 29791 39457
rect 33045 39491 33103 39497
rect 33045 39457 33057 39491
rect 33091 39457 33103 39491
rect 39022 39488 39028 39500
rect 38983 39460 39028 39488
rect 33045 39451 33103 39457
rect 39022 39448 39028 39460
rect 39080 39448 39086 39500
rect 39482 39488 39488 39500
rect 39443 39460 39488 39488
rect 39482 39448 39488 39460
rect 39540 39448 39546 39500
rect 39577 39491 39635 39497
rect 39577 39457 39589 39491
rect 39623 39488 39635 39491
rect 39942 39488 39948 39500
rect 39623 39460 39948 39488
rect 39623 39457 39635 39460
rect 39577 39451 39635 39457
rect 39942 39448 39948 39460
rect 40000 39488 40006 39500
rect 40313 39491 40371 39497
rect 40313 39488 40325 39491
rect 40000 39460 40325 39488
rect 40000 39448 40006 39460
rect 40313 39457 40325 39460
rect 40359 39488 40371 39491
rect 43806 39488 43812 39500
rect 40359 39460 43812 39488
rect 40359 39457 40371 39460
rect 40313 39451 40371 39457
rect 43806 39448 43812 39460
rect 43864 39448 43870 39500
rect 44174 39488 44180 39500
rect 44135 39460 44180 39488
rect 44174 39448 44180 39460
rect 44232 39488 44238 39500
rect 44232 39460 44404 39488
rect 44232 39448 44238 39460
rect 28258 39420 28264 39432
rect 28219 39392 28264 39420
rect 28258 39380 28264 39392
rect 28316 39380 28322 39432
rect 33318 39420 33324 39432
rect 33279 39392 33324 39420
rect 33318 39380 33324 39392
rect 33376 39380 33382 39432
rect 38930 39420 38936 39432
rect 38891 39392 38936 39420
rect 38930 39380 38936 39392
rect 38988 39380 38994 39432
rect 44269 39423 44327 39429
rect 44269 39389 44281 39423
rect 44315 39389 44327 39423
rect 44376 39420 44404 39460
rect 44450 39448 44456 39500
rect 44508 39488 44514 39500
rect 44910 39488 44916 39500
rect 44508 39460 44553 39488
rect 44652 39460 44916 39488
rect 44508 39448 44514 39460
rect 44652 39420 44680 39460
rect 44910 39448 44916 39460
rect 44968 39448 44974 39500
rect 46492 39497 46520 39528
rect 45005 39491 45063 39497
rect 45005 39457 45017 39491
rect 45051 39488 45063 39491
rect 46477 39491 46535 39497
rect 45051 39460 46060 39488
rect 45051 39457 45063 39460
rect 45005 39451 45063 39457
rect 46032 39429 46060 39460
rect 46477 39457 46489 39491
rect 46523 39457 46535 39491
rect 46477 39451 46535 39457
rect 46661 39491 46719 39497
rect 46661 39457 46673 39491
rect 46707 39457 46719 39491
rect 46661 39451 46719 39457
rect 44376 39392 44680 39420
rect 46017 39423 46075 39429
rect 44269 39383 44327 39389
rect 46017 39389 46029 39423
rect 46063 39420 46075 39423
rect 46566 39420 46572 39432
rect 46063 39392 46572 39420
rect 46063 39389 46075 39392
rect 46017 39383 46075 39389
rect 26694 39352 26700 39364
rect 21416 39324 26700 39352
rect 21416 39312 21422 39324
rect 26694 39312 26700 39324
rect 26752 39312 26758 39364
rect 20993 39287 21051 39293
rect 20993 39284 21005 39287
rect 20772 39256 21005 39284
rect 20772 39244 20778 39256
rect 20993 39253 21005 39256
rect 21039 39253 21051 39287
rect 29546 39284 29552 39296
rect 29507 39256 29552 39284
rect 20993 39247 21051 39253
rect 29546 39244 29552 39256
rect 29604 39244 29610 39296
rect 34606 39284 34612 39296
rect 34567 39256 34612 39284
rect 34606 39244 34612 39256
rect 34664 39284 34670 39296
rect 39574 39284 39580 39296
rect 34664 39256 39580 39284
rect 34664 39244 34670 39256
rect 39574 39244 39580 39256
rect 39632 39244 39638 39296
rect 40034 39284 40040 39296
rect 39995 39256 40040 39284
rect 40034 39244 40040 39256
rect 40092 39244 40098 39296
rect 40589 39287 40647 39293
rect 40589 39253 40601 39287
rect 40635 39284 40647 39287
rect 40678 39284 40684 39296
rect 40635 39256 40684 39284
rect 40635 39253 40647 39256
rect 40589 39247 40647 39253
rect 40678 39244 40684 39256
rect 40736 39244 40742 39296
rect 42610 39244 42616 39296
rect 42668 39284 42674 39296
rect 43993 39287 44051 39293
rect 43993 39284 44005 39287
rect 42668 39256 44005 39284
rect 42668 39244 42674 39256
rect 43993 39253 44005 39256
rect 44039 39284 44051 39287
rect 44284 39284 44312 39383
rect 46566 39380 46572 39392
rect 46624 39420 46630 39432
rect 46676 39420 46704 39451
rect 47026 39448 47032 39500
rect 47084 39488 47090 39500
rect 47228 39497 47256 39596
rect 48038 39584 48044 39596
rect 48096 39624 48102 39636
rect 48225 39627 48283 39633
rect 48225 39624 48237 39627
rect 48096 39596 48237 39624
rect 48096 39584 48102 39596
rect 48225 39593 48237 39596
rect 48271 39624 48283 39627
rect 48271 39596 55904 39624
rect 48271 39593 48283 39596
rect 48225 39587 48283 39593
rect 48130 39516 48136 39568
rect 48188 39556 48194 39568
rect 48409 39559 48467 39565
rect 48409 39556 48421 39559
rect 48188 39528 48421 39556
rect 48188 39516 48194 39528
rect 48409 39525 48421 39528
rect 48455 39556 48467 39559
rect 48774 39556 48780 39568
rect 48455 39528 48780 39556
rect 48455 39525 48467 39528
rect 48409 39519 48467 39525
rect 48774 39516 48780 39528
rect 48832 39516 48838 39568
rect 48866 39516 48872 39568
rect 48924 39556 48930 39568
rect 54386 39556 54392 39568
rect 48924 39528 54392 39556
rect 48924 39516 48930 39528
rect 54386 39516 54392 39528
rect 54444 39516 54450 39568
rect 54478 39516 54484 39568
rect 54536 39556 54542 39568
rect 54573 39559 54631 39565
rect 54573 39556 54585 39559
rect 54536 39528 54585 39556
rect 54536 39516 54542 39528
rect 54573 39525 54585 39528
rect 54619 39525 54631 39559
rect 55214 39556 55220 39568
rect 54573 39519 54631 39525
rect 54680 39528 55220 39556
rect 47213 39491 47271 39497
rect 47213 39488 47225 39491
rect 47084 39460 47225 39488
rect 47084 39448 47090 39460
rect 47213 39457 47225 39460
rect 47259 39457 47271 39491
rect 47394 39488 47400 39500
rect 47355 39460 47400 39488
rect 47213 39451 47271 39457
rect 47394 39448 47400 39460
rect 47452 39448 47458 39500
rect 47578 39448 47584 39500
rect 47636 39488 47642 39500
rect 51810 39488 51816 39500
rect 47636 39460 51816 39488
rect 47636 39448 47642 39460
rect 51810 39448 51816 39460
rect 51868 39448 51874 39500
rect 52270 39488 52276 39500
rect 52231 39460 52276 39488
rect 52270 39448 52276 39460
rect 52328 39448 52334 39500
rect 52733 39491 52791 39497
rect 52733 39488 52745 39491
rect 52380 39460 52745 39488
rect 48130 39420 48136 39432
rect 46624 39392 46704 39420
rect 46624 39380 46630 39392
rect 46676 39352 46704 39392
rect 47596 39392 48136 39420
rect 47596 39352 47624 39392
rect 48130 39380 48136 39392
rect 48188 39380 48194 39432
rect 51718 39380 51724 39432
rect 51776 39420 51782 39432
rect 52089 39423 52147 39429
rect 52089 39420 52101 39423
rect 51776 39392 52101 39420
rect 51776 39380 51782 39392
rect 52089 39389 52101 39392
rect 52135 39420 52147 39423
rect 52380 39420 52408 39460
rect 52733 39457 52745 39460
rect 52779 39457 52791 39491
rect 52733 39451 52791 39457
rect 52822 39448 52828 39500
rect 52880 39488 52886 39500
rect 52880 39460 53696 39488
rect 52880 39448 52886 39460
rect 53668 39432 53696 39460
rect 53650 39420 53656 39432
rect 52135 39392 52408 39420
rect 53563 39392 53656 39420
rect 52135 39389 52147 39392
rect 52089 39383 52147 39389
rect 53650 39380 53656 39392
rect 53708 39420 53714 39432
rect 53837 39423 53895 39429
rect 53837 39420 53849 39423
rect 53708 39392 53849 39420
rect 53708 39380 53714 39392
rect 53837 39389 53849 39392
rect 53883 39420 53895 39423
rect 54680 39420 54708 39528
rect 55214 39516 55220 39528
rect 55272 39516 55278 39568
rect 55876 39556 55904 39596
rect 58434 39584 58440 39636
rect 58492 39624 58498 39636
rect 59909 39627 59967 39633
rect 59909 39624 59921 39627
rect 58492 39596 59921 39624
rect 58492 39584 58498 39596
rect 59909 39593 59921 39596
rect 59955 39624 59967 39627
rect 60366 39624 60372 39636
rect 59955 39596 60372 39624
rect 59955 39593 59967 39596
rect 59909 39587 59967 39593
rect 60366 39584 60372 39596
rect 60424 39584 60430 39636
rect 60826 39584 60832 39636
rect 60884 39624 60890 39636
rect 60884 39596 60964 39624
rect 60884 39584 60890 39596
rect 60734 39556 60740 39568
rect 55876 39528 60740 39556
rect 60734 39516 60740 39528
rect 60792 39516 60798 39568
rect 54846 39448 54852 39500
rect 54904 39488 54910 39500
rect 60826 39488 60832 39500
rect 54904 39460 60688 39488
rect 60787 39460 60832 39488
rect 54904 39448 54910 39460
rect 53883 39392 54708 39420
rect 53883 39389 53895 39392
rect 53837 39383 53895 39389
rect 54938 39380 54944 39432
rect 54996 39420 55002 39432
rect 54996 39392 55038 39420
rect 54996 39380 55002 39392
rect 55214 39380 55220 39432
rect 55272 39420 55278 39432
rect 60550 39420 60556 39432
rect 55272 39392 60556 39420
rect 55272 39380 55278 39392
rect 60550 39380 60556 39392
rect 60608 39380 60614 39432
rect 46676 39324 47624 39352
rect 47673 39355 47731 39361
rect 47673 39321 47685 39355
rect 47719 39352 47731 39355
rect 54202 39352 54208 39364
rect 47719 39324 54208 39352
rect 47719 39321 47731 39324
rect 47673 39315 47731 39321
rect 54202 39312 54208 39324
rect 54260 39312 54266 39364
rect 54570 39312 54576 39364
rect 54628 39352 54634 39364
rect 54711 39355 54769 39361
rect 54711 39352 54723 39355
rect 54628 39324 54723 39352
rect 54628 39312 54634 39324
rect 54711 39321 54723 39324
rect 54757 39321 54769 39355
rect 60090 39352 60096 39364
rect 54711 39315 54769 39321
rect 55140 39324 60096 39352
rect 47302 39284 47308 39296
rect 44039 39256 47308 39284
rect 44039 39253 44051 39256
rect 43993 39247 44051 39253
rect 47302 39244 47308 39256
rect 47360 39244 47366 39296
rect 47394 39244 47400 39296
rect 47452 39284 47458 39296
rect 47854 39284 47860 39296
rect 47452 39256 47860 39284
rect 47452 39244 47458 39256
rect 47854 39244 47860 39256
rect 47912 39284 47918 39296
rect 47949 39287 48007 39293
rect 47949 39284 47961 39287
rect 47912 39256 47961 39284
rect 47912 39244 47918 39256
rect 47949 39253 47961 39256
rect 47995 39253 48007 39287
rect 51718 39284 51724 39296
rect 51679 39256 51724 39284
rect 47949 39247 48007 39253
rect 51718 39244 51724 39256
rect 51776 39284 51782 39296
rect 51905 39287 51963 39293
rect 51905 39284 51917 39287
rect 51776 39256 51917 39284
rect 51776 39244 51782 39256
rect 51905 39253 51917 39256
rect 51951 39253 51963 39287
rect 51905 39247 51963 39253
rect 52270 39244 52276 39296
rect 52328 39284 52334 39296
rect 52822 39284 52828 39296
rect 52328 39256 52828 39284
rect 52328 39244 52334 39256
rect 52822 39244 52828 39256
rect 52880 39244 52886 39296
rect 53282 39284 53288 39296
rect 53243 39256 53288 39284
rect 53282 39244 53288 39256
rect 53340 39244 53346 39296
rect 54849 39287 54907 39293
rect 54849 39253 54861 39287
rect 54895 39284 54907 39287
rect 55140 39284 55168 39324
rect 60090 39312 60096 39324
rect 60148 39312 60154 39364
rect 60660 39352 60688 39460
rect 60826 39448 60832 39460
rect 60884 39448 60890 39500
rect 60936 39429 60964 39596
rect 67358 39584 67364 39636
rect 67416 39624 67422 39636
rect 69750 39624 69756 39636
rect 67416 39596 69756 39624
rect 67416 39584 67422 39596
rect 69750 39584 69756 39596
rect 69808 39584 69814 39636
rect 71682 39584 71688 39636
rect 71740 39624 71746 39636
rect 71740 39596 71912 39624
rect 71740 39584 71746 39596
rect 65981 39559 66039 39565
rect 65981 39525 65993 39559
rect 66027 39556 66039 39559
rect 66070 39556 66076 39568
rect 66027 39528 66076 39556
rect 66027 39525 66039 39528
rect 65981 39519 66039 39525
rect 66070 39516 66076 39528
rect 66128 39516 66134 39568
rect 71590 39516 71596 39568
rect 71648 39556 71654 39568
rect 71884 39556 71912 39596
rect 71958 39584 71964 39636
rect 72016 39624 72022 39636
rect 72237 39627 72295 39633
rect 72237 39624 72249 39627
rect 72016 39596 72249 39624
rect 72016 39584 72022 39596
rect 72237 39593 72249 39596
rect 72283 39593 72295 39627
rect 72237 39587 72295 39593
rect 72510 39584 72516 39636
rect 72568 39624 72574 39636
rect 73249 39627 73307 39633
rect 73249 39624 73261 39627
rect 72568 39596 73261 39624
rect 72568 39584 72574 39596
rect 73249 39593 73261 39596
rect 73295 39593 73307 39627
rect 77754 39624 77760 39636
rect 77715 39596 77760 39624
rect 73249 39587 73307 39593
rect 77754 39584 77760 39596
rect 77812 39584 77818 39636
rect 83366 39584 83372 39636
rect 83424 39624 83430 39636
rect 84013 39627 84071 39633
rect 84013 39624 84025 39627
rect 83424 39596 84025 39624
rect 83424 39584 83430 39596
rect 84013 39593 84025 39596
rect 84059 39593 84071 39627
rect 84013 39587 84071 39593
rect 72973 39559 73031 39565
rect 72973 39556 72985 39559
rect 71648 39528 71693 39556
rect 71884 39528 72985 39556
rect 71648 39516 71654 39528
rect 72973 39525 72985 39528
rect 73019 39525 73031 39559
rect 72973 39519 73031 39525
rect 61194 39488 61200 39500
rect 61155 39460 61200 39488
rect 61194 39448 61200 39460
rect 61252 39448 61258 39500
rect 61381 39491 61439 39497
rect 61381 39457 61393 39491
rect 61427 39488 61439 39491
rect 61562 39488 61568 39500
rect 61427 39460 61568 39488
rect 61427 39457 61439 39460
rect 61381 39451 61439 39457
rect 61562 39448 61568 39460
rect 61620 39488 61626 39500
rect 61930 39488 61936 39500
rect 61620 39460 61936 39488
rect 61620 39448 61626 39460
rect 61930 39448 61936 39460
rect 61988 39448 61994 39500
rect 65518 39448 65524 39500
rect 65576 39488 65582 39500
rect 65889 39491 65947 39497
rect 65889 39488 65901 39491
rect 65576 39460 65901 39488
rect 65576 39448 65582 39460
rect 65889 39457 65901 39460
rect 65935 39488 65947 39491
rect 66806 39488 66812 39500
rect 65935 39460 66812 39488
rect 65935 39457 65947 39460
rect 65889 39451 65947 39457
rect 66806 39448 66812 39460
rect 66864 39448 66870 39500
rect 66993 39491 67051 39497
rect 66993 39457 67005 39491
rect 67039 39488 67051 39491
rect 67085 39491 67143 39497
rect 67085 39488 67097 39491
rect 67039 39460 67097 39488
rect 67039 39457 67051 39460
rect 66993 39451 67051 39457
rect 67085 39457 67097 39460
rect 67131 39488 67143 39491
rect 67450 39488 67456 39500
rect 67131 39460 67456 39488
rect 67131 39457 67143 39460
rect 67085 39451 67143 39457
rect 67450 39448 67456 39460
rect 67508 39448 67514 39500
rect 71406 39448 71412 39500
rect 71464 39488 71470 39500
rect 71774 39488 71780 39500
rect 71464 39460 71780 39488
rect 71464 39448 71470 39460
rect 71774 39448 71780 39460
rect 71832 39448 71838 39500
rect 72142 39488 72148 39500
rect 72103 39460 72148 39488
rect 72142 39448 72148 39460
rect 72200 39448 72206 39500
rect 73157 39491 73215 39497
rect 73157 39488 73169 39491
rect 72804 39460 73169 39488
rect 60921 39423 60979 39429
rect 60921 39389 60933 39423
rect 60967 39389 60979 39423
rect 60921 39383 60979 39389
rect 67361 39423 67419 39429
rect 67361 39389 67373 39423
rect 67407 39420 67419 39423
rect 68830 39420 68836 39432
rect 67407 39392 68836 39420
rect 67407 39389 67419 39392
rect 67361 39383 67419 39389
rect 68830 39380 68836 39392
rect 68888 39380 68894 39432
rect 71590 39380 71596 39432
rect 71648 39420 71654 39432
rect 71958 39420 71964 39432
rect 71648 39392 71964 39420
rect 71648 39380 71654 39392
rect 71958 39380 71964 39392
rect 72016 39380 72022 39432
rect 66070 39352 66076 39364
rect 60660 39324 66076 39352
rect 66070 39312 66076 39324
rect 66128 39312 66134 39364
rect 71130 39312 71136 39364
rect 71188 39352 71194 39364
rect 72418 39352 72424 39364
rect 71188 39324 72424 39352
rect 71188 39312 71194 39324
rect 72418 39312 72424 39324
rect 72476 39352 72482 39364
rect 72804 39361 72832 39460
rect 73157 39457 73169 39460
rect 73203 39457 73215 39491
rect 77772 39488 77800 39584
rect 78125 39559 78183 39565
rect 78125 39525 78137 39559
rect 78171 39556 78183 39559
rect 79686 39556 79692 39568
rect 78171 39528 79692 39556
rect 78171 39525 78183 39528
rect 78125 39519 78183 39525
rect 79686 39516 79692 39528
rect 79744 39516 79750 39568
rect 77941 39491 77999 39497
rect 77941 39488 77953 39491
rect 77772 39460 77953 39488
rect 73157 39451 73215 39457
rect 77941 39457 77953 39460
rect 77987 39457 77999 39491
rect 78214 39488 78220 39500
rect 78175 39460 78220 39488
rect 77941 39451 77999 39457
rect 78214 39448 78220 39460
rect 78272 39448 78278 39500
rect 84028 39488 84056 39587
rect 84197 39491 84255 39497
rect 84197 39488 84209 39491
rect 84028 39460 84209 39488
rect 84197 39457 84209 39460
rect 84243 39488 84255 39491
rect 86310 39488 86316 39500
rect 84243 39460 86316 39488
rect 84243 39457 84255 39460
rect 84197 39451 84255 39457
rect 86310 39448 86316 39460
rect 86368 39448 86374 39500
rect 84378 39380 84384 39432
rect 84436 39420 84442 39432
rect 84473 39423 84531 39429
rect 84473 39420 84485 39423
rect 84436 39392 84485 39420
rect 84436 39380 84442 39392
rect 84473 39389 84485 39392
rect 84519 39389 84531 39423
rect 84473 39383 84531 39389
rect 72789 39355 72847 39361
rect 72789 39352 72801 39355
rect 72476 39324 72801 39352
rect 72476 39312 72482 39324
rect 72789 39321 72801 39324
rect 72835 39321 72847 39355
rect 72789 39315 72847 39321
rect 54895 39256 55168 39284
rect 55217 39287 55275 39293
rect 54895 39253 54907 39256
rect 54849 39247 54907 39253
rect 55217 39253 55229 39287
rect 55263 39284 55275 39287
rect 57882 39284 57888 39296
rect 55263 39256 57888 39284
rect 55263 39253 55275 39256
rect 55217 39247 55275 39253
rect 57882 39244 57888 39256
rect 57940 39244 57946 39296
rect 60274 39284 60280 39296
rect 60235 39256 60280 39284
rect 60274 39244 60280 39256
rect 60332 39244 60338 39296
rect 60366 39244 60372 39296
rect 60424 39284 60430 39296
rect 61194 39284 61200 39296
rect 60424 39256 61200 39284
rect 60424 39244 60430 39256
rect 61194 39244 61200 39256
rect 61252 39244 61258 39296
rect 66898 39244 66904 39296
rect 66956 39284 66962 39296
rect 68465 39287 68523 39293
rect 68465 39284 68477 39287
rect 66956 39256 68477 39284
rect 66956 39244 66962 39256
rect 68465 39253 68477 39256
rect 68511 39253 68523 39287
rect 71406 39284 71412 39296
rect 71367 39256 71412 39284
rect 68465 39247 68523 39253
rect 71406 39244 71412 39256
rect 71464 39244 71470 39296
rect 78398 39284 78404 39296
rect 78359 39256 78404 39284
rect 78398 39244 78404 39256
rect 78456 39244 78462 39296
rect 85390 39244 85396 39296
rect 85448 39284 85454 39296
rect 85577 39287 85635 39293
rect 85577 39284 85589 39287
rect 85448 39256 85589 39284
rect 85448 39244 85454 39256
rect 85577 39253 85589 39256
rect 85623 39253 85635 39287
rect 85577 39247 85635 39253
rect 1104 39194 108008 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 65686 39194
rect 65738 39142 65750 39194
rect 65802 39142 65814 39194
rect 65866 39142 65878 39194
rect 65930 39142 96406 39194
rect 96458 39142 96470 39194
rect 96522 39142 96534 39194
rect 96586 39142 96598 39194
rect 96650 39142 108008 39194
rect 1104 39120 108008 39142
rect 4525 39083 4583 39089
rect 4525 39049 4537 39083
rect 4571 39080 4583 39083
rect 4614 39080 4620 39092
rect 4571 39052 4620 39080
rect 4571 39049 4583 39052
rect 4525 39043 4583 39049
rect 4614 39040 4620 39052
rect 4672 39040 4678 39092
rect 4798 39080 4804 39092
rect 4759 39052 4804 39080
rect 4798 39040 4804 39052
rect 4856 39040 4862 39092
rect 9858 39080 9864 39092
rect 8680 39052 9864 39080
rect 2961 38947 3019 38953
rect 2961 38913 2973 38947
rect 3007 38944 3019 38947
rect 4798 38944 4804 38956
rect 3007 38916 4804 38944
rect 3007 38913 3019 38916
rect 2961 38907 3019 38913
rect 4798 38904 4804 38916
rect 4856 38904 4862 38956
rect 3237 38879 3295 38885
rect 3237 38845 3249 38879
rect 3283 38876 3295 38879
rect 4614 38876 4620 38888
rect 3283 38848 4620 38876
rect 3283 38845 3295 38848
rect 3237 38839 3295 38845
rect 4614 38836 4620 38848
rect 4672 38836 4678 38888
rect 8297 38879 8355 38885
rect 8297 38876 8309 38879
rect 8128 38848 8309 38876
rect 3510 38700 3516 38752
rect 3568 38740 3574 38752
rect 8128 38749 8156 38848
rect 8297 38845 8309 38848
rect 8343 38845 8355 38879
rect 8297 38839 8355 38845
rect 8481 38879 8539 38885
rect 8481 38845 8493 38879
rect 8527 38845 8539 38879
rect 8680 38876 8708 39052
rect 9858 39040 9864 39052
rect 9916 39040 9922 39092
rect 13538 39040 13544 39092
rect 13596 39080 13602 39092
rect 13814 39080 13820 39092
rect 13596 39052 13820 39080
rect 13596 39040 13602 39052
rect 13814 39040 13820 39052
rect 13872 39040 13878 39092
rect 14645 39083 14703 39089
rect 14645 39049 14657 39083
rect 14691 39080 14703 39083
rect 17126 39080 17132 39092
rect 14691 39052 17132 39080
rect 14691 39049 14703 39052
rect 14645 39043 14703 39049
rect 17126 39040 17132 39052
rect 17184 39040 17190 39092
rect 22186 39040 22192 39092
rect 22244 39080 22250 39092
rect 23753 39083 23811 39089
rect 23753 39080 23765 39083
rect 22244 39052 23765 39080
rect 22244 39040 22250 39052
rect 23753 39049 23765 39052
rect 23799 39080 23811 39083
rect 28442 39080 28448 39092
rect 23799 39052 28304 39080
rect 28403 39052 28448 39080
rect 23799 39049 23811 39052
rect 23753 39043 23811 39049
rect 9398 39012 9404 39024
rect 9359 38984 9404 39012
rect 9398 38972 9404 38984
rect 9456 38972 9462 39024
rect 10226 38972 10232 39024
rect 10284 39012 10290 39024
rect 15102 39012 15108 39024
rect 10284 38984 15108 39012
rect 10284 38972 10290 38984
rect 15102 38972 15108 38984
rect 15160 38972 15166 39024
rect 16022 39012 16028 39024
rect 15983 38984 16028 39012
rect 16022 38972 16028 38984
rect 16080 38972 16086 39024
rect 26694 38972 26700 39024
rect 26752 39012 26758 39024
rect 28169 39015 28227 39021
rect 28169 39012 28181 39015
rect 26752 38984 28181 39012
rect 26752 38972 26758 38984
rect 28169 38981 28181 38984
rect 28215 38981 28227 39015
rect 28276 39012 28304 39052
rect 28442 39040 28448 39052
rect 28500 39040 28506 39092
rect 29546 39040 29552 39092
rect 29604 39080 29610 39092
rect 53098 39080 53104 39092
rect 29604 39052 53104 39080
rect 29604 39040 29610 39052
rect 53098 39040 53104 39052
rect 53156 39040 53162 39092
rect 53282 39040 53288 39092
rect 53340 39080 53346 39092
rect 54481 39083 54539 39089
rect 54481 39080 54493 39083
rect 53340 39052 54493 39080
rect 53340 39040 53346 39052
rect 54481 39049 54493 39052
rect 54527 39049 54539 39083
rect 54662 39080 54668 39092
rect 54623 39052 54668 39080
rect 54481 39043 54539 39049
rect 54662 39040 54668 39052
rect 54720 39040 54726 39092
rect 72973 39083 73031 39089
rect 54772 39052 72924 39080
rect 42150 39012 42156 39024
rect 28276 38984 42156 39012
rect 28169 38975 28227 38981
rect 42150 38972 42156 38984
rect 42208 38972 42214 39024
rect 44910 38972 44916 39024
rect 44968 39012 44974 39024
rect 46106 39012 46112 39024
rect 44968 38984 46112 39012
rect 44968 38972 44974 38984
rect 46106 38972 46112 38984
rect 46164 38972 46170 39024
rect 46216 38984 53144 39012
rect 39022 38904 39028 38956
rect 39080 38944 39086 38956
rect 40402 38944 40408 38956
rect 39080 38916 40408 38944
rect 39080 38904 39086 38916
rect 40402 38904 40408 38916
rect 40460 38944 40466 38956
rect 40678 38944 40684 38956
rect 40460 38916 40684 38944
rect 40460 38904 40466 38916
rect 40678 38904 40684 38916
rect 40736 38944 40742 38956
rect 46216 38944 46244 38984
rect 40736 38916 46244 38944
rect 40736 38904 40742 38916
rect 46382 38904 46388 38956
rect 46440 38944 46446 38956
rect 48038 38944 48044 38956
rect 46440 38916 46485 38944
rect 47999 38916 48044 38944
rect 46440 38904 46446 38916
rect 48038 38904 48044 38916
rect 48096 38904 48102 38956
rect 48130 38904 48136 38956
rect 48188 38944 48194 38956
rect 53116 38944 53144 38984
rect 53374 38972 53380 39024
rect 53432 39012 53438 39024
rect 54343 39015 54401 39021
rect 54343 39012 54355 39015
rect 53432 38984 54355 39012
rect 53432 38972 53438 38984
rect 54343 38981 54355 38984
rect 54389 38981 54401 39015
rect 54343 38975 54401 38981
rect 54570 38944 54576 38956
rect 48188 38916 48233 38944
rect 53116 38916 54340 38944
rect 54531 38916 54576 38944
rect 48188 38904 48194 38916
rect 8941 38879 8999 38885
rect 8941 38876 8953 38879
rect 8680 38848 8953 38876
rect 8481 38839 8539 38845
rect 8941 38845 8953 38848
rect 8987 38845 8999 38879
rect 8941 38839 8999 38845
rect 9033 38879 9091 38885
rect 9033 38845 9045 38879
rect 9079 38876 9091 38879
rect 10226 38876 10232 38888
rect 9079 38848 10232 38876
rect 9079 38845 9091 38848
rect 9033 38839 9091 38845
rect 8496 38808 8524 38839
rect 9048 38808 9076 38839
rect 10226 38836 10232 38848
rect 10284 38836 10290 38888
rect 14001 38879 14059 38885
rect 14001 38845 14013 38879
rect 14047 38876 14059 38879
rect 14645 38879 14703 38885
rect 14645 38876 14657 38879
rect 14047 38848 14657 38876
rect 14047 38845 14059 38848
rect 14001 38839 14059 38845
rect 14645 38845 14657 38848
rect 14691 38845 14703 38879
rect 14645 38839 14703 38845
rect 14921 38879 14979 38885
rect 14921 38845 14933 38879
rect 14967 38845 14979 38879
rect 15102 38876 15108 38888
rect 15063 38848 15108 38876
rect 14921 38839 14979 38845
rect 8496 38780 9076 38808
rect 8113 38743 8171 38749
rect 8113 38740 8125 38743
rect 3568 38712 8125 38740
rect 3568 38700 3574 38712
rect 8113 38709 8125 38712
rect 8159 38709 8171 38743
rect 8113 38703 8171 38709
rect 14829 38743 14887 38749
rect 14829 38709 14841 38743
rect 14875 38740 14887 38743
rect 14936 38740 14964 38839
rect 15102 38836 15108 38848
rect 15160 38836 15166 38888
rect 15562 38876 15568 38888
rect 15523 38848 15568 38876
rect 15562 38836 15568 38848
rect 15620 38836 15626 38888
rect 15657 38879 15715 38885
rect 15657 38845 15669 38879
rect 15703 38876 15715 38879
rect 21358 38876 21364 38888
rect 15703 38848 21364 38876
rect 15703 38845 15715 38848
rect 15657 38839 15715 38845
rect 21358 38836 21364 38848
rect 21416 38836 21422 38888
rect 23658 38876 23664 38888
rect 23619 38848 23664 38876
rect 23658 38836 23664 38848
rect 23716 38836 23722 38888
rect 27985 38879 28043 38885
rect 27985 38845 27997 38879
rect 28031 38876 28043 38879
rect 28442 38876 28448 38888
rect 28031 38848 28448 38876
rect 28031 38845 28043 38848
rect 27985 38839 28043 38845
rect 28442 38836 28448 38848
rect 28500 38836 28506 38888
rect 36541 38879 36599 38885
rect 36541 38845 36553 38879
rect 36587 38876 36599 38879
rect 36725 38879 36783 38885
rect 36725 38876 36737 38879
rect 36587 38848 36737 38876
rect 36587 38845 36599 38848
rect 36541 38839 36599 38845
rect 36725 38845 36737 38848
rect 36771 38876 36783 38879
rect 44726 38876 44732 38888
rect 36771 38848 44732 38876
rect 36771 38845 36783 38848
rect 36725 38839 36783 38845
rect 44726 38836 44732 38848
rect 44784 38836 44790 38888
rect 46477 38879 46535 38885
rect 46477 38845 46489 38879
rect 46523 38876 46535 38879
rect 46566 38876 46572 38888
rect 46523 38848 46572 38876
rect 46523 38845 46535 38848
rect 46477 38839 46535 38845
rect 46566 38836 46572 38848
rect 46624 38836 46630 38888
rect 47026 38876 47032 38888
rect 46987 38848 47032 38876
rect 47026 38836 47032 38848
rect 47084 38836 47090 38888
rect 47118 38836 47124 38888
rect 47176 38876 47182 38888
rect 47213 38879 47271 38885
rect 47213 38876 47225 38879
rect 47176 38848 47225 38876
rect 47176 38836 47182 38848
rect 47213 38845 47225 38848
rect 47259 38845 47271 38879
rect 47213 38839 47271 38845
rect 51997 38879 52055 38885
rect 51997 38845 52009 38879
rect 52043 38845 52055 38879
rect 51997 38839 52055 38845
rect 52181 38879 52239 38885
rect 52181 38845 52193 38879
rect 52227 38876 52239 38879
rect 52270 38876 52276 38888
rect 52227 38848 52276 38876
rect 52227 38845 52239 38848
rect 52181 38839 52239 38845
rect 17862 38768 17868 38820
rect 17920 38808 17926 38820
rect 47581 38811 47639 38817
rect 17920 38780 36584 38808
rect 17920 38768 17926 38780
rect 15102 38740 15108 38752
rect 14875 38712 15108 38740
rect 14875 38709 14887 38712
rect 14829 38703 14887 38709
rect 15102 38700 15108 38712
rect 15160 38700 15166 38752
rect 36354 38740 36360 38752
rect 36315 38712 36360 38740
rect 36354 38700 36360 38712
rect 36412 38700 36418 38752
rect 36556 38740 36584 38780
rect 47581 38777 47593 38811
rect 47627 38808 47639 38811
rect 49234 38808 49240 38820
rect 47627 38780 49240 38808
rect 47627 38777 47639 38780
rect 47581 38771 47639 38777
rect 49234 38768 49240 38780
rect 49292 38768 49298 38820
rect 51442 38768 51448 38820
rect 51500 38808 51506 38820
rect 51537 38811 51595 38817
rect 51537 38808 51549 38811
rect 51500 38780 51549 38808
rect 51500 38768 51506 38780
rect 51537 38777 51549 38780
rect 51583 38808 51595 38811
rect 51905 38811 51963 38817
rect 51905 38808 51917 38811
rect 51583 38780 51917 38808
rect 51583 38777 51595 38780
rect 51537 38771 51595 38777
rect 51905 38777 51917 38780
rect 51951 38808 51963 38811
rect 52012 38808 52040 38839
rect 52270 38836 52276 38848
rect 52328 38836 52334 38888
rect 52641 38879 52699 38885
rect 52641 38845 52653 38879
rect 52687 38845 52699 38879
rect 52641 38839 52699 38845
rect 52733 38879 52791 38885
rect 52733 38845 52745 38879
rect 52779 38845 52791 38879
rect 53561 38879 53619 38885
rect 53561 38876 53573 38879
rect 52733 38839 52791 38845
rect 53024 38848 53573 38876
rect 52656 38808 52684 38839
rect 51951 38780 52684 38808
rect 52748 38808 52776 38839
rect 53024 38808 53052 38848
rect 53561 38845 53573 38848
rect 53607 38876 53619 38879
rect 53650 38876 53656 38888
rect 53607 38848 53656 38876
rect 53607 38845 53619 38848
rect 53561 38839 53619 38845
rect 53650 38836 53656 38848
rect 53708 38836 53714 38888
rect 54202 38876 54208 38888
rect 54163 38848 54208 38876
rect 54202 38836 54208 38848
rect 54260 38836 54266 38888
rect 54312 38876 54340 38916
rect 54570 38904 54576 38916
rect 54628 38904 54634 38956
rect 54772 38876 54800 39052
rect 58066 38972 58072 39024
rect 58124 39012 58130 39024
rect 58345 39015 58403 39021
rect 58345 39012 58357 39015
rect 58124 38984 58357 39012
rect 58124 38972 58130 38984
rect 58345 38981 58357 38984
rect 58391 38981 58403 39015
rect 59170 39012 59176 39024
rect 58345 38975 58403 38981
rect 58728 38984 59176 39012
rect 58360 38944 58388 38975
rect 58529 38947 58587 38953
rect 58529 38944 58541 38947
rect 58360 38916 58541 38944
rect 58529 38913 58541 38916
rect 58575 38913 58587 38947
rect 58529 38907 58587 38913
rect 58728 38885 58756 38984
rect 59170 38972 59176 38984
rect 59228 38972 59234 39024
rect 59446 38972 59452 39024
rect 59504 39012 59510 39024
rect 60553 39015 60611 39021
rect 60553 39012 60565 39015
rect 59504 38984 60565 39012
rect 59504 38972 59510 38984
rect 60553 38981 60565 38984
rect 60599 39012 60611 39015
rect 61470 39012 61476 39024
rect 60599 38984 61476 39012
rect 60599 38981 60611 38984
rect 60553 38975 60611 38981
rect 61470 38972 61476 38984
rect 61528 38972 61534 39024
rect 62117 39015 62175 39021
rect 62117 38981 62129 39015
rect 62163 39012 62175 39015
rect 68370 39012 68376 39024
rect 62163 38984 68376 39012
rect 62163 38981 62175 38984
rect 62117 38975 62175 38981
rect 59817 38947 59875 38953
rect 59817 38913 59829 38947
rect 59863 38944 59875 38947
rect 61289 38947 61347 38953
rect 61289 38944 61301 38947
rect 59863 38916 61301 38944
rect 59863 38913 59875 38916
rect 59817 38907 59875 38913
rect 61289 38913 61301 38916
rect 61335 38913 61347 38947
rect 62132 38944 62160 38975
rect 68370 38972 68376 38984
rect 68428 38972 68434 39024
rect 68830 39012 68836 39024
rect 68791 38984 68836 39012
rect 68830 38972 68836 38984
rect 68888 38972 68894 39024
rect 69750 38972 69756 39024
rect 69808 39012 69814 39024
rect 72896 39012 72924 39052
rect 72973 39049 72985 39083
rect 73019 39080 73031 39083
rect 73062 39080 73068 39092
rect 73019 39052 73068 39080
rect 73019 39049 73031 39052
rect 72973 39043 73031 39049
rect 73062 39040 73068 39052
rect 73120 39040 73126 39092
rect 77754 39080 77760 39092
rect 76024 39052 77760 39080
rect 76024 39012 76052 39052
rect 77754 39040 77760 39052
rect 77812 39080 77818 39092
rect 78677 39083 78735 39089
rect 78677 39080 78689 39083
rect 77812 39052 78689 39080
rect 77812 39040 77818 39052
rect 78677 39049 78689 39052
rect 78723 39049 78735 39083
rect 84378 39080 84384 39092
rect 84339 39052 84384 39080
rect 78677 39043 78735 39049
rect 84378 39040 84384 39052
rect 84436 39040 84442 39092
rect 86310 39080 86316 39092
rect 86271 39052 86316 39080
rect 86310 39040 86316 39052
rect 86368 39040 86374 39092
rect 69808 38984 72464 39012
rect 72896 38984 76052 39012
rect 77021 39015 77079 39021
rect 69808 38972 69814 38984
rect 61289 38907 61347 38913
rect 61396 38916 62160 38944
rect 64785 38947 64843 38953
rect 54312 38848 54800 38876
rect 58713 38879 58771 38885
rect 58713 38845 58725 38879
rect 58759 38845 58771 38879
rect 59078 38876 59084 38888
rect 58713 38839 58771 38845
rect 59004 38848 59084 38876
rect 52748 38780 53052 38808
rect 51951 38777 51963 38780
rect 51905 38771 51963 38777
rect 53098 38768 53104 38820
rect 53156 38808 53162 38820
rect 59004 38808 59032 38848
rect 59078 38836 59084 38848
rect 59136 38836 59142 38888
rect 59173 38879 59231 38885
rect 59173 38845 59185 38879
rect 59219 38845 59231 38879
rect 59173 38839 59231 38845
rect 59265 38879 59323 38885
rect 59265 38845 59277 38879
rect 59311 38845 59323 38879
rect 59265 38839 59323 38845
rect 53156 38780 59032 38808
rect 53156 38768 53162 38780
rect 46842 38740 46848 38752
rect 36556 38712 46848 38740
rect 46842 38700 46848 38712
rect 46900 38700 46906 38752
rect 47118 38700 47124 38752
rect 47176 38740 47182 38752
rect 47765 38743 47823 38749
rect 47765 38740 47777 38743
rect 47176 38712 47777 38740
rect 47176 38700 47182 38712
rect 47765 38709 47777 38712
rect 47811 38709 47823 38743
rect 47765 38703 47823 38709
rect 52730 38700 52736 38752
rect 52788 38740 52794 38752
rect 53193 38743 53251 38749
rect 53193 38740 53205 38743
rect 52788 38712 53205 38740
rect 52788 38700 52794 38712
rect 53193 38709 53205 38712
rect 53239 38709 53251 38743
rect 53193 38703 53251 38709
rect 54386 38700 54392 38752
rect 54444 38740 54450 38752
rect 58253 38743 58311 38749
rect 58253 38740 58265 38743
rect 54444 38712 58265 38740
rect 54444 38700 54450 38712
rect 58253 38709 58265 38712
rect 58299 38740 58311 38743
rect 59188 38740 59216 38839
rect 58299 38712 59216 38740
rect 59280 38740 59308 38839
rect 59446 38836 59452 38888
rect 59504 38876 59510 38888
rect 61396 38885 61424 38916
rect 64785 38913 64797 38947
rect 64831 38944 64843 38947
rect 65978 38944 65984 38956
rect 64831 38916 65984 38944
rect 64831 38913 64843 38916
rect 64785 38907 64843 38913
rect 65978 38904 65984 38916
rect 66036 38904 66042 38956
rect 66070 38904 66076 38956
rect 66128 38944 66134 38956
rect 69290 38944 69296 38956
rect 66128 38916 69296 38944
rect 66128 38904 66134 38916
rect 69290 38904 69296 38916
rect 69348 38904 69354 38956
rect 71406 38904 71412 38956
rect 71464 38944 71470 38956
rect 71464 38916 71912 38944
rect 71464 38904 71470 38916
rect 61381 38879 61439 38885
rect 59504 38848 61332 38876
rect 59504 38836 59510 38848
rect 59722 38768 59728 38820
rect 59780 38808 59786 38820
rect 60737 38811 60795 38817
rect 60737 38808 60749 38811
rect 59780 38780 60749 38808
rect 59780 38768 59786 38780
rect 60737 38777 60749 38780
rect 60783 38777 60795 38811
rect 61304 38808 61332 38848
rect 61381 38845 61393 38879
rect 61427 38845 61439 38879
rect 61381 38839 61439 38845
rect 61654 38836 61660 38888
rect 61712 38876 61718 38888
rect 61749 38879 61807 38885
rect 61749 38876 61761 38879
rect 61712 38848 61761 38876
rect 61712 38836 61718 38848
rect 61749 38845 61761 38848
rect 61795 38845 61807 38879
rect 61930 38876 61936 38888
rect 61891 38848 61936 38876
rect 61749 38839 61807 38845
rect 61930 38836 61936 38848
rect 61988 38836 61994 38888
rect 64966 38876 64972 38888
rect 64927 38848 64972 38876
rect 64966 38836 64972 38848
rect 65024 38836 65030 38888
rect 65150 38876 65156 38888
rect 65111 38848 65156 38876
rect 65150 38836 65156 38848
rect 65208 38836 65214 38888
rect 65518 38876 65524 38888
rect 65479 38848 65524 38876
rect 65518 38836 65524 38848
rect 65576 38836 65582 38888
rect 65613 38879 65671 38885
rect 65613 38845 65625 38879
rect 65659 38845 65671 38879
rect 66898 38876 66904 38888
rect 66859 38848 66904 38876
rect 65613 38839 65671 38845
rect 64230 38808 64236 38820
rect 61304 38780 64236 38808
rect 60737 38771 60795 38777
rect 64230 38768 64236 38780
rect 64288 38808 64294 38820
rect 64325 38811 64383 38817
rect 64325 38808 64337 38811
rect 64288 38780 64337 38808
rect 64288 38768 64294 38780
rect 64325 38777 64337 38780
rect 64371 38808 64383 38811
rect 65628 38808 65656 38839
rect 66898 38836 66904 38848
rect 66956 38876 66962 38888
rect 67177 38879 67235 38885
rect 67177 38876 67189 38879
rect 66956 38848 67189 38876
rect 66956 38836 66962 38848
rect 67177 38845 67189 38848
rect 67223 38845 67235 38879
rect 67177 38839 67235 38845
rect 68741 38879 68799 38885
rect 68741 38845 68753 38879
rect 68787 38876 68799 38879
rect 71041 38879 71099 38885
rect 71041 38876 71053 38879
rect 68787 38848 71053 38876
rect 68787 38845 68799 38848
rect 68741 38839 68799 38845
rect 71041 38845 71053 38848
rect 71087 38845 71099 38879
rect 71682 38876 71688 38888
rect 71643 38848 71688 38876
rect 71041 38839 71099 38845
rect 71682 38836 71688 38848
rect 71740 38836 71746 38888
rect 71777 38879 71835 38885
rect 71777 38845 71789 38879
rect 71823 38845 71835 38879
rect 71884 38876 71912 38916
rect 71958 38904 71964 38956
rect 72016 38944 72022 38956
rect 72145 38947 72203 38953
rect 72145 38944 72157 38947
rect 72016 38916 72157 38944
rect 72016 38904 72022 38916
rect 72145 38913 72157 38916
rect 72191 38944 72203 38947
rect 72329 38947 72387 38953
rect 72329 38944 72341 38947
rect 72191 38916 72341 38944
rect 72191 38913 72203 38916
rect 72145 38907 72203 38913
rect 72329 38913 72341 38916
rect 72375 38913 72387 38947
rect 72436 38944 72464 38984
rect 77021 38981 77033 39015
rect 77067 39012 77079 39015
rect 77110 39012 77116 39024
rect 77067 38984 77116 39012
rect 77067 38981 77079 38984
rect 77021 38975 77079 38981
rect 77110 38972 77116 38984
rect 77168 38972 77174 39024
rect 77389 38947 77447 38953
rect 72436 38916 77340 38944
rect 72329 38907 72387 38913
rect 72053 38879 72111 38885
rect 72053 38876 72065 38879
rect 71884 38848 72065 38876
rect 71777 38839 71835 38845
rect 72053 38845 72065 38848
rect 72099 38845 72111 38879
rect 72344 38876 72372 38907
rect 72786 38876 72792 38888
rect 72344 38848 72792 38876
rect 72053 38839 72111 38845
rect 64371 38780 65656 38808
rect 71792 38808 71820 38839
rect 72786 38836 72792 38848
rect 72844 38836 72850 38888
rect 73062 38876 73068 38888
rect 73023 38848 73068 38876
rect 73062 38836 73068 38848
rect 73120 38836 73126 38888
rect 77110 38876 77116 38888
rect 77071 38848 77116 38876
rect 77110 38836 77116 38848
rect 77168 38836 77174 38888
rect 77312 38876 77340 38916
rect 77389 38913 77401 38947
rect 77435 38944 77447 38947
rect 78398 38944 78404 38956
rect 77435 38916 78404 38944
rect 77435 38913 77447 38916
rect 77389 38907 77447 38913
rect 78398 38904 78404 38916
rect 78456 38904 78462 38956
rect 80149 38947 80207 38953
rect 80149 38913 80161 38947
rect 80195 38944 80207 38947
rect 87877 38947 87935 38953
rect 87877 38944 87889 38947
rect 80195 38916 87889 38944
rect 80195 38913 80207 38916
rect 80149 38907 80207 38913
rect 87877 38913 87889 38916
rect 87923 38913 87935 38947
rect 87877 38907 87935 38913
rect 79042 38876 79048 38888
rect 77312 38848 79048 38876
rect 79042 38836 79048 38848
rect 79100 38836 79106 38888
rect 79594 38836 79600 38888
rect 79652 38876 79658 38888
rect 79781 38879 79839 38885
rect 79781 38876 79793 38879
rect 79652 38848 79793 38876
rect 79652 38836 79658 38848
rect 79781 38845 79793 38848
rect 79827 38876 79839 38879
rect 80164 38876 80192 38907
rect 79827 38848 80192 38876
rect 79827 38845 79839 38848
rect 79781 38839 79839 38845
rect 82262 38836 82268 38888
rect 82320 38876 82326 38888
rect 83185 38879 83243 38885
rect 83185 38876 83197 38879
rect 82320 38848 83197 38876
rect 82320 38836 82326 38848
rect 83185 38845 83197 38848
rect 83231 38876 83243 38879
rect 83553 38879 83611 38885
rect 83553 38876 83565 38879
rect 83231 38848 83565 38876
rect 83231 38845 83243 38848
rect 83185 38839 83243 38845
rect 83553 38845 83565 38848
rect 83599 38845 83611 38879
rect 84286 38876 84292 38888
rect 84247 38848 84292 38876
rect 83553 38839 83611 38845
rect 83568 38808 83596 38839
rect 84286 38836 84292 38848
rect 84344 38836 84350 38888
rect 85390 38876 85396 38888
rect 85351 38848 85396 38876
rect 85390 38836 85396 38848
rect 85448 38836 85454 38888
rect 86310 38836 86316 38888
rect 86368 38876 86374 38888
rect 86497 38879 86555 38885
rect 86497 38876 86509 38879
rect 86368 38848 86509 38876
rect 86368 38836 86374 38848
rect 86497 38845 86509 38848
rect 86543 38845 86555 38879
rect 86770 38876 86776 38888
rect 86731 38848 86776 38876
rect 86497 38839 86555 38845
rect 86770 38836 86776 38848
rect 86828 38836 86834 38888
rect 84746 38808 84752 38820
rect 71792 38780 72648 38808
rect 83568 38780 84752 38808
rect 64371 38777 64383 38780
rect 64325 38771 64383 38777
rect 72620 38752 72648 38780
rect 84746 38768 84752 38780
rect 84804 38808 84810 38820
rect 85485 38811 85543 38817
rect 85485 38808 85497 38811
rect 84804 38780 85497 38808
rect 84804 38768 84810 38780
rect 85485 38777 85497 38780
rect 85531 38777 85543 38811
rect 85485 38771 85543 38777
rect 59998 38740 60004 38752
rect 59280 38712 60004 38740
rect 58299 38709 58311 38712
rect 58253 38703 58311 38709
rect 59998 38700 60004 38712
rect 60056 38700 60062 38752
rect 60090 38700 60096 38752
rect 60148 38740 60154 38752
rect 61378 38740 61384 38752
rect 60148 38712 61384 38740
rect 60148 38700 60154 38712
rect 61378 38700 61384 38712
rect 61436 38700 61442 38752
rect 64966 38700 64972 38752
rect 65024 38740 65030 38752
rect 65797 38743 65855 38749
rect 65797 38740 65809 38743
rect 65024 38712 65809 38740
rect 65024 38700 65030 38712
rect 65797 38709 65809 38712
rect 65843 38709 65855 38743
rect 65797 38703 65855 38709
rect 66993 38743 67051 38749
rect 66993 38709 67005 38743
rect 67039 38740 67051 38743
rect 68278 38740 68284 38752
rect 67039 38712 68284 38740
rect 67039 38709 67051 38712
rect 66993 38703 67051 38709
rect 68278 38700 68284 38712
rect 68336 38740 68342 38752
rect 70857 38743 70915 38749
rect 70857 38740 70869 38743
rect 68336 38712 70869 38740
rect 68336 38700 68342 38712
rect 70857 38709 70869 38712
rect 70903 38740 70915 38743
rect 71406 38740 71412 38752
rect 70903 38712 71412 38740
rect 70903 38709 70915 38712
rect 70857 38703 70915 38709
rect 71406 38700 71412 38712
rect 71464 38700 71470 38752
rect 72602 38740 72608 38752
rect 72563 38712 72608 38740
rect 72602 38700 72608 38712
rect 72660 38700 72666 38752
rect 73154 38740 73160 38752
rect 73115 38712 73160 38740
rect 73154 38700 73160 38712
rect 73212 38700 73218 38752
rect 79870 38740 79876 38752
rect 79831 38712 79876 38740
rect 79870 38700 79876 38712
rect 79928 38700 79934 38752
rect 83366 38740 83372 38752
rect 83327 38712 83372 38740
rect 83366 38700 83372 38712
rect 83424 38700 83430 38752
rect 1104 38650 108008 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 81046 38650
rect 81098 38598 81110 38650
rect 81162 38598 81174 38650
rect 81226 38598 81238 38650
rect 81290 38598 108008 38650
rect 1104 38576 108008 38598
rect 4062 38496 4068 38548
rect 4120 38536 4126 38548
rect 23750 38536 23756 38548
rect 4120 38508 23756 38536
rect 4120 38496 4126 38508
rect 23750 38496 23756 38508
rect 23808 38496 23814 38548
rect 28169 38539 28227 38545
rect 28169 38536 28181 38539
rect 27632 38508 28181 38536
rect 12250 38428 12256 38480
rect 12308 38468 12314 38480
rect 17589 38471 17647 38477
rect 17589 38468 17601 38471
rect 12308 38440 15608 38468
rect 12308 38428 12314 38440
rect 10594 38360 10600 38412
rect 10652 38400 10658 38412
rect 10781 38403 10839 38409
rect 10781 38400 10793 38403
rect 10652 38372 10793 38400
rect 10652 38360 10658 38372
rect 10781 38369 10793 38372
rect 10827 38400 10839 38403
rect 12621 38403 12679 38409
rect 10827 38372 12112 38400
rect 10827 38369 10839 38372
rect 10781 38363 10839 38369
rect 11054 38332 11060 38344
rect 11015 38304 11060 38332
rect 11054 38292 11060 38304
rect 11112 38292 11118 38344
rect 12084 38264 12112 38372
rect 12621 38369 12633 38403
rect 12667 38400 12679 38403
rect 13814 38400 13820 38412
rect 12667 38372 13820 38400
rect 12667 38369 12679 38372
rect 12621 38363 12679 38369
rect 12636 38264 12664 38363
rect 13814 38360 13820 38372
rect 13872 38360 13878 38412
rect 15458 38403 15516 38409
rect 15458 38369 15470 38403
rect 15504 38400 15516 38403
rect 15580 38400 15608 38440
rect 16224 38440 17601 38468
rect 16224 38412 16252 38440
rect 17589 38437 17601 38440
rect 17635 38437 17647 38471
rect 17862 38468 17868 38480
rect 17823 38440 17868 38468
rect 17589 38431 17647 38437
rect 17862 38428 17868 38440
rect 17920 38428 17926 38480
rect 20806 38428 20812 38480
rect 20864 38468 20870 38480
rect 21082 38468 21088 38480
rect 20864 38440 21088 38468
rect 20864 38428 20870 38440
rect 21082 38428 21088 38440
rect 21140 38468 21146 38480
rect 21269 38471 21327 38477
rect 21269 38468 21281 38471
rect 21140 38440 21281 38468
rect 21140 38428 21146 38440
rect 21269 38437 21281 38440
rect 21315 38437 21327 38471
rect 21269 38431 21327 38437
rect 23109 38471 23167 38477
rect 23109 38437 23121 38471
rect 23155 38468 23167 38471
rect 23658 38468 23664 38480
rect 23155 38440 23664 38468
rect 23155 38437 23167 38440
rect 23109 38431 23167 38437
rect 15838 38400 15844 38412
rect 15504 38372 15844 38400
rect 15504 38369 15516 38372
rect 15458 38363 15516 38369
rect 15838 38360 15844 38372
rect 15896 38360 15902 38412
rect 16022 38400 16028 38412
rect 15983 38372 16028 38400
rect 16022 38360 16028 38372
rect 16080 38360 16086 38412
rect 16206 38400 16212 38412
rect 16167 38372 16212 38400
rect 16206 38360 16212 38372
rect 16264 38360 16270 38412
rect 17497 38403 17555 38409
rect 17497 38369 17509 38403
rect 17543 38400 17555 38403
rect 17880 38400 17908 38428
rect 17543 38372 17908 38400
rect 21284 38400 21312 38431
rect 23658 38428 23664 38440
rect 23716 38428 23722 38480
rect 26234 38428 26240 38480
rect 26292 38468 26298 38480
rect 27632 38468 27660 38508
rect 28169 38505 28181 38508
rect 28215 38536 28227 38539
rect 28215 38508 36584 38536
rect 28215 38505 28227 38508
rect 28169 38499 28227 38505
rect 26292 38440 27660 38468
rect 26292 38428 26298 38440
rect 21453 38403 21511 38409
rect 21453 38400 21465 38403
rect 21284 38372 21465 38400
rect 17543 38369 17555 38372
rect 17497 38363 17555 38369
rect 21453 38369 21465 38372
rect 21499 38369 21511 38403
rect 21453 38363 21511 38369
rect 15289 38335 15347 38341
rect 15289 38332 15301 38335
rect 12084 38236 12664 38264
rect 15120 38304 15301 38332
rect 15120 38208 15148 38304
rect 15289 38301 15301 38304
rect 15335 38301 15347 38335
rect 15289 38295 15347 38301
rect 16390 38264 16396 38276
rect 16351 38236 16396 38264
rect 16390 38224 16396 38236
rect 16448 38224 16454 38276
rect 5074 38156 5080 38208
rect 5132 38196 5138 38208
rect 12250 38196 12256 38208
rect 5132 38168 12256 38196
rect 5132 38156 5138 38168
rect 12250 38156 12256 38168
rect 12308 38156 12314 38208
rect 12345 38199 12403 38205
rect 12345 38165 12357 38199
rect 12391 38196 12403 38199
rect 12434 38196 12440 38208
rect 12391 38168 12440 38196
rect 12391 38165 12403 38168
rect 12345 38159 12403 38165
rect 12434 38156 12440 38168
rect 12492 38156 12498 38208
rect 15102 38196 15108 38208
rect 15063 38168 15108 38196
rect 15102 38156 15108 38168
rect 15160 38156 15166 38208
rect 15838 38156 15844 38208
rect 15896 38196 15902 38208
rect 16761 38199 16819 38205
rect 16761 38196 16773 38199
rect 15896 38168 16773 38196
rect 15896 38156 15902 38168
rect 16761 38165 16773 38168
rect 16807 38165 16819 38199
rect 21468 38196 21496 38363
rect 26694 38360 26700 38412
rect 26752 38400 26758 38412
rect 26789 38403 26847 38409
rect 26789 38400 26801 38403
rect 26752 38372 26801 38400
rect 26752 38360 26758 38372
rect 26789 38369 26801 38372
rect 26835 38400 26847 38403
rect 27341 38403 27399 38409
rect 27341 38400 27353 38403
rect 26835 38372 27353 38400
rect 26835 38369 26847 38372
rect 26789 38363 26847 38369
rect 27341 38369 27353 38372
rect 27387 38369 27399 38403
rect 27341 38363 27399 38369
rect 27525 38403 27583 38409
rect 27525 38369 27537 38403
rect 27571 38400 27583 38403
rect 27632 38400 27660 38440
rect 27893 38471 27951 38477
rect 27893 38437 27905 38471
rect 27939 38468 27951 38471
rect 28258 38468 28264 38480
rect 27939 38440 28264 38468
rect 27939 38437 27951 38440
rect 27893 38431 27951 38437
rect 28258 38428 28264 38440
rect 28316 38428 28322 38480
rect 36556 38468 36584 38508
rect 37090 38496 37096 38548
rect 37148 38536 37154 38548
rect 40218 38536 40224 38548
rect 37148 38508 40224 38536
rect 37148 38496 37154 38508
rect 40218 38496 40224 38508
rect 40276 38496 40282 38548
rect 40402 38536 40408 38548
rect 40363 38508 40408 38536
rect 40402 38496 40408 38508
rect 40460 38496 40466 38548
rect 40954 38496 40960 38548
rect 41012 38536 41018 38548
rect 51810 38536 51816 38548
rect 41012 38508 51816 38536
rect 41012 38496 41018 38508
rect 51810 38496 51816 38508
rect 51868 38496 51874 38548
rect 53101 38539 53159 38545
rect 53101 38505 53113 38539
rect 53147 38536 53159 38539
rect 54938 38536 54944 38548
rect 53147 38508 54944 38536
rect 53147 38505 53159 38508
rect 53101 38499 53159 38505
rect 54938 38496 54944 38508
rect 54996 38496 55002 38548
rect 55030 38496 55036 38548
rect 55088 38536 55094 38548
rect 72418 38536 72424 38548
rect 55088 38508 72188 38536
rect 72379 38508 72424 38536
rect 55088 38496 55094 38508
rect 64509 38471 64567 38477
rect 64509 38468 64521 38471
rect 36556 38440 64521 38468
rect 64509 38437 64521 38440
rect 64555 38468 64567 38471
rect 64966 38468 64972 38480
rect 64555 38440 64972 38468
rect 64555 38437 64567 38440
rect 64509 38431 64567 38437
rect 64966 38428 64972 38440
rect 65024 38428 65030 38480
rect 71682 38468 71688 38480
rect 65168 38440 71688 38468
rect 27571 38372 27660 38400
rect 27571 38369 27583 38372
rect 27525 38363 27583 38369
rect 38470 38360 38476 38412
rect 38528 38400 38534 38412
rect 38933 38403 38991 38409
rect 38528 38372 38884 38400
rect 38528 38360 38534 38372
rect 21726 38332 21732 38344
rect 21687 38304 21732 38332
rect 21726 38292 21732 38304
rect 21784 38292 21790 38344
rect 26513 38335 26571 38341
rect 26513 38301 26525 38335
rect 26559 38332 26571 38335
rect 26605 38335 26663 38341
rect 26605 38332 26617 38335
rect 26559 38304 26617 38332
rect 26559 38301 26571 38304
rect 26513 38295 26571 38301
rect 26605 38301 26617 38304
rect 26651 38301 26663 38335
rect 33137 38335 33195 38341
rect 33137 38332 33149 38335
rect 26605 38295 26663 38301
rect 32968 38304 33149 38332
rect 23842 38224 23848 38276
rect 23900 38264 23906 38276
rect 32766 38264 32772 38276
rect 23900 38236 32772 38264
rect 23900 38224 23906 38236
rect 32766 38224 32772 38236
rect 32824 38224 32830 38276
rect 32968 38208 32996 38304
rect 33137 38301 33149 38304
rect 33183 38301 33195 38335
rect 33410 38332 33416 38344
rect 33371 38304 33416 38332
rect 33137 38295 33195 38301
rect 33410 38292 33416 38304
rect 33468 38292 33474 38344
rect 38746 38332 38752 38344
rect 38707 38304 38752 38332
rect 38746 38292 38752 38304
rect 38804 38292 38810 38344
rect 38856 38332 38884 38372
rect 38933 38369 38945 38403
rect 38979 38400 38991 38403
rect 39022 38400 39028 38412
rect 38979 38372 39028 38400
rect 38979 38369 38991 38372
rect 38933 38363 38991 38369
rect 39022 38360 39028 38372
rect 39080 38360 39086 38412
rect 39393 38403 39451 38409
rect 39393 38400 39405 38403
rect 39132 38372 39405 38400
rect 39132 38332 39160 38372
rect 39393 38369 39405 38372
rect 39439 38369 39451 38403
rect 39393 38363 39451 38369
rect 39485 38403 39543 38409
rect 39485 38369 39497 38403
rect 39531 38400 39543 38403
rect 39531 38372 39896 38400
rect 39531 38369 39543 38372
rect 39485 38363 39543 38369
rect 38856 38304 39160 38332
rect 39868 38332 39896 38372
rect 40218 38360 40224 38412
rect 40276 38400 40282 38412
rect 40681 38403 40739 38409
rect 40681 38400 40693 38403
rect 40276 38372 40693 38400
rect 40276 38360 40282 38372
rect 40681 38369 40693 38372
rect 40727 38400 40739 38403
rect 40773 38403 40831 38409
rect 40773 38400 40785 38403
rect 40727 38372 40785 38400
rect 40727 38369 40739 38372
rect 40681 38363 40739 38369
rect 40773 38369 40785 38372
rect 40819 38369 40831 38403
rect 40773 38363 40831 38369
rect 40957 38403 41015 38409
rect 40957 38369 40969 38403
rect 41003 38400 41015 38403
rect 41230 38400 41236 38412
rect 41003 38372 41236 38400
rect 41003 38369 41015 38372
rect 40957 38363 41015 38369
rect 41230 38360 41236 38372
rect 41288 38360 41294 38412
rect 49234 38360 49240 38412
rect 49292 38400 49298 38412
rect 52638 38409 52644 38412
rect 52457 38403 52515 38409
rect 52457 38400 52469 38403
rect 49292 38372 52469 38400
rect 49292 38360 49298 38372
rect 52457 38369 52469 38372
rect 52503 38369 52515 38403
rect 52457 38363 52515 38369
rect 52604 38403 52644 38409
rect 52604 38369 52616 38403
rect 52604 38363 52644 38369
rect 52638 38360 52644 38363
rect 52696 38360 52702 38412
rect 57882 38360 57888 38412
rect 57940 38400 57946 38412
rect 60185 38403 60243 38409
rect 60185 38400 60197 38403
rect 57940 38372 60197 38400
rect 57940 38360 57946 38372
rect 60185 38369 60197 38372
rect 60231 38369 60243 38403
rect 60185 38363 60243 38369
rect 60274 38360 60280 38412
rect 60332 38409 60338 38412
rect 60332 38403 60390 38409
rect 60332 38369 60344 38403
rect 60378 38369 60390 38403
rect 62206 38400 62212 38412
rect 60332 38363 60390 38369
rect 60568 38372 62212 38400
rect 60332 38360 60338 38363
rect 39942 38332 39948 38344
rect 39868 38304 39948 38332
rect 39942 38292 39948 38304
rect 40000 38292 40006 38344
rect 40034 38292 40040 38344
rect 40092 38332 40098 38344
rect 41325 38335 41383 38341
rect 41325 38332 41337 38335
rect 40092 38304 41337 38332
rect 40092 38292 40098 38304
rect 41325 38301 41337 38304
rect 41371 38301 41383 38335
rect 41325 38295 41383 38301
rect 46014 38292 46020 38344
rect 46072 38332 46078 38344
rect 52362 38332 52368 38344
rect 46072 38304 52368 38332
rect 46072 38292 46078 38304
rect 52362 38292 52368 38304
rect 52420 38292 52426 38344
rect 52825 38335 52883 38341
rect 52825 38301 52837 38335
rect 52871 38332 52883 38335
rect 53098 38332 53104 38344
rect 52871 38304 53104 38332
rect 52871 38301 52883 38304
rect 52825 38295 52883 38301
rect 53098 38292 53104 38304
rect 53156 38292 53162 38344
rect 58710 38292 58716 38344
rect 58768 38332 58774 38344
rect 59722 38332 59728 38344
rect 58768 38304 59728 38332
rect 58768 38292 58774 38304
rect 59722 38292 59728 38304
rect 59780 38292 59786 38344
rect 60568 38341 60596 38372
rect 62206 38360 62212 38372
rect 62264 38360 62270 38412
rect 64230 38400 64236 38412
rect 64191 38372 64236 38400
rect 64230 38360 64236 38372
rect 64288 38400 64294 38412
rect 64417 38403 64475 38409
rect 64417 38400 64429 38403
rect 64288 38372 64429 38400
rect 64288 38360 64294 38372
rect 64417 38369 64429 38372
rect 64463 38369 64475 38403
rect 64417 38363 64475 38369
rect 60553 38335 60611 38341
rect 60553 38301 60565 38335
rect 60599 38301 60611 38335
rect 60553 38295 60611 38301
rect 60734 38292 60740 38344
rect 60792 38332 60798 38344
rect 65168 38332 65196 38440
rect 71682 38428 71688 38440
rect 71740 38428 71746 38480
rect 65613 38403 65671 38409
rect 65613 38400 65625 38403
rect 60792 38304 65196 38332
rect 65260 38372 65625 38400
rect 60792 38292 60798 38304
rect 34701 38267 34759 38273
rect 34701 38233 34713 38267
rect 34747 38264 34759 38267
rect 34790 38264 34796 38276
rect 34747 38236 34796 38264
rect 34747 38233 34759 38236
rect 34701 38227 34759 38233
rect 34790 38224 34796 38236
rect 34848 38264 34854 38276
rect 39114 38264 39120 38276
rect 34848 38236 39120 38264
rect 34848 38224 34854 38236
rect 39114 38224 39120 38236
rect 39172 38224 39178 38276
rect 39850 38264 39856 38276
rect 39811 38236 39856 38264
rect 39850 38224 39856 38236
rect 39908 38224 39914 38276
rect 40862 38264 40868 38276
rect 39960 38236 40868 38264
rect 24670 38196 24676 38208
rect 21468 38168 24676 38196
rect 16761 38159 16819 38165
rect 24670 38156 24676 38168
rect 24728 38156 24734 38208
rect 25498 38156 25504 38208
rect 25556 38196 25562 38208
rect 26237 38199 26295 38205
rect 26237 38196 26249 38199
rect 25556 38168 26249 38196
rect 25556 38156 25562 38168
rect 26237 38165 26249 38168
rect 26283 38196 26295 38199
rect 26513 38199 26571 38205
rect 26513 38196 26525 38199
rect 26283 38168 26525 38196
rect 26283 38165 26295 38168
rect 26237 38159 26295 38165
rect 26513 38165 26525 38168
rect 26559 38165 26571 38199
rect 32950 38196 32956 38208
rect 32911 38168 32956 38196
rect 26513 38159 26571 38165
rect 32950 38156 32956 38168
rect 33008 38196 33014 38208
rect 38286 38196 38292 38208
rect 33008 38168 38292 38196
rect 33008 38156 33014 38168
rect 38286 38156 38292 38168
rect 38344 38156 38350 38208
rect 38838 38156 38844 38208
rect 38896 38196 38902 38208
rect 39960 38196 39988 38236
rect 40862 38224 40868 38236
rect 40920 38224 40926 38276
rect 52730 38264 52736 38276
rect 52691 38236 52736 38264
rect 52730 38224 52736 38236
rect 52788 38224 52794 38276
rect 65260 38273 65288 38372
rect 65613 38369 65625 38372
rect 65659 38369 65671 38403
rect 65613 38363 65671 38369
rect 72160 38332 72188 38508
rect 72418 38496 72424 38508
rect 72476 38496 72482 38548
rect 76650 38536 76656 38548
rect 76563 38508 76656 38536
rect 76650 38496 76656 38508
rect 76708 38536 76714 38548
rect 77110 38536 77116 38548
rect 76708 38508 77116 38536
rect 76708 38496 76714 38508
rect 77110 38496 77116 38508
rect 77168 38496 77174 38548
rect 79042 38496 79048 38548
rect 79100 38536 79106 38548
rect 79781 38539 79839 38545
rect 79781 38536 79793 38539
rect 79100 38508 79793 38536
rect 79100 38496 79106 38508
rect 79781 38505 79793 38508
rect 79827 38536 79839 38539
rect 79962 38536 79968 38548
rect 79827 38508 79968 38536
rect 79827 38505 79839 38508
rect 79781 38499 79839 38505
rect 79962 38496 79968 38508
rect 80020 38496 80026 38548
rect 83366 38496 83372 38548
rect 83424 38536 83430 38548
rect 84381 38539 84439 38545
rect 84381 38536 84393 38539
rect 83424 38508 84393 38536
rect 83424 38496 83430 38508
rect 84381 38505 84393 38508
rect 84427 38505 84439 38539
rect 84381 38499 84439 38505
rect 73522 38468 73528 38480
rect 72252 38440 73528 38468
rect 72252 38409 72280 38440
rect 73522 38428 73528 38440
rect 73580 38428 73586 38480
rect 79134 38468 79140 38480
rect 77588 38440 79140 38468
rect 72237 38403 72295 38409
rect 72237 38369 72249 38403
rect 72283 38369 72295 38403
rect 72237 38363 72295 38369
rect 73154 38360 73160 38412
rect 73212 38400 73218 38412
rect 73341 38403 73399 38409
rect 73341 38400 73353 38403
rect 73212 38372 73353 38400
rect 73212 38360 73218 38372
rect 73341 38369 73353 38372
rect 73387 38369 73399 38403
rect 73341 38363 73399 38369
rect 76006 38360 76012 38412
rect 76064 38400 76070 38412
rect 77588 38409 77616 38440
rect 79134 38428 79140 38440
rect 79192 38428 79198 38480
rect 79686 38468 79692 38480
rect 79647 38440 79692 38468
rect 79686 38428 79692 38440
rect 79744 38428 79750 38480
rect 83093 38471 83151 38477
rect 83093 38437 83105 38471
rect 83139 38468 83151 38471
rect 84286 38468 84292 38480
rect 83139 38440 84292 38468
rect 83139 38437 83151 38440
rect 83093 38431 83151 38437
rect 84286 38428 84292 38440
rect 84344 38428 84350 38480
rect 76837 38403 76895 38409
rect 76837 38400 76849 38403
rect 76064 38372 76849 38400
rect 76064 38360 76070 38372
rect 76837 38369 76849 38372
rect 76883 38369 76895 38403
rect 76837 38363 76895 38369
rect 77573 38403 77631 38409
rect 77573 38369 77585 38403
rect 77619 38369 77631 38403
rect 77941 38403 77999 38409
rect 77941 38400 77953 38403
rect 77573 38363 77631 38369
rect 77680 38372 77953 38400
rect 77478 38332 77484 38344
rect 72160 38304 77484 38332
rect 77478 38292 77484 38304
rect 77536 38332 77542 38344
rect 77680 38332 77708 38372
rect 77941 38369 77953 38372
rect 77987 38400 77999 38403
rect 78309 38403 78367 38409
rect 78309 38400 78321 38403
rect 77987 38372 78321 38400
rect 77987 38369 77999 38372
rect 77941 38363 77999 38369
rect 78309 38369 78321 38372
rect 78355 38400 78367 38403
rect 78585 38403 78643 38409
rect 78585 38400 78597 38403
rect 78355 38372 78597 38400
rect 78355 38369 78367 38372
rect 78309 38363 78367 38369
rect 78585 38369 78597 38372
rect 78631 38369 78643 38403
rect 78585 38363 78643 38369
rect 78953 38403 79011 38409
rect 78953 38369 78965 38403
rect 78999 38400 79011 38403
rect 79778 38400 79784 38412
rect 78999 38372 79784 38400
rect 78999 38369 79011 38372
rect 78953 38363 79011 38369
rect 77536 38304 77708 38332
rect 77757 38335 77815 38341
rect 77536 38292 77542 38304
rect 77757 38301 77769 38335
rect 77803 38332 77815 38335
rect 78214 38332 78220 38344
rect 77803 38304 78220 38332
rect 77803 38301 77815 38304
rect 77757 38295 77815 38301
rect 78214 38292 78220 38304
rect 78272 38292 78278 38344
rect 59909 38267 59967 38273
rect 59909 38264 59921 38267
rect 52840 38236 59921 38264
rect 38896 38168 39988 38196
rect 38896 38156 38902 38168
rect 40034 38156 40040 38208
rect 40092 38196 40098 38208
rect 40221 38199 40279 38205
rect 40221 38196 40233 38199
rect 40092 38168 40233 38196
rect 40092 38156 40098 38168
rect 40221 38165 40233 38168
rect 40267 38165 40279 38199
rect 40221 38159 40279 38165
rect 40681 38199 40739 38205
rect 40681 38165 40693 38199
rect 40727 38196 40739 38199
rect 41095 38199 41153 38205
rect 41095 38196 41107 38199
rect 40727 38168 41107 38196
rect 40727 38165 40739 38168
rect 40681 38159 40739 38165
rect 41095 38165 41107 38168
rect 41141 38165 41153 38199
rect 41095 38159 41153 38165
rect 41230 38156 41236 38208
rect 41288 38196 41294 38208
rect 41601 38199 41659 38205
rect 41288 38168 41333 38196
rect 41288 38156 41294 38168
rect 41601 38165 41613 38199
rect 41647 38196 41659 38199
rect 52840 38196 52868 38236
rect 59909 38233 59921 38236
rect 59955 38264 59967 38267
rect 60461 38267 60519 38273
rect 60461 38264 60473 38267
rect 59955 38236 60473 38264
rect 59955 38233 59967 38236
rect 59909 38227 59967 38233
rect 60461 38233 60473 38236
rect 60507 38233 60519 38267
rect 65245 38267 65303 38273
rect 65245 38264 65257 38267
rect 60461 38227 60519 38233
rect 60568 38236 65257 38264
rect 41647 38168 52868 38196
rect 41647 38165 41659 38168
rect 41601 38159 41659 38165
rect 55306 38156 55312 38208
rect 55364 38196 55370 38208
rect 60568 38196 60596 38236
rect 65245 38233 65257 38236
rect 65291 38233 65303 38267
rect 66254 38264 66260 38276
rect 65245 38227 65303 38233
rect 65352 38236 66260 38264
rect 60826 38196 60832 38208
rect 55364 38168 60596 38196
rect 60787 38168 60832 38196
rect 55364 38156 55370 38168
rect 60826 38156 60832 38168
rect 60884 38156 60890 38208
rect 62206 38156 62212 38208
rect 62264 38196 62270 38208
rect 65352 38196 65380 38236
rect 66254 38224 66260 38236
rect 66312 38224 66318 38276
rect 73338 38224 73344 38276
rect 73396 38264 73402 38276
rect 73525 38267 73583 38273
rect 73525 38264 73537 38267
rect 73396 38236 73537 38264
rect 73396 38224 73402 38236
rect 73525 38233 73537 38236
rect 73571 38233 73583 38267
rect 78600 38264 78628 38363
rect 79778 38360 79784 38372
rect 79836 38360 79842 38412
rect 80330 38360 80336 38412
rect 80388 38400 80394 38412
rect 80517 38403 80575 38409
rect 80517 38400 80529 38403
rect 80388 38372 80529 38400
rect 80388 38360 80394 38372
rect 80517 38369 80529 38372
rect 80563 38369 80575 38403
rect 80517 38363 80575 38369
rect 80609 38403 80667 38409
rect 80609 38369 80621 38403
rect 80655 38400 80667 38403
rect 80882 38400 80888 38412
rect 80655 38372 80888 38400
rect 80655 38369 80667 38372
rect 80609 38363 80667 38369
rect 80882 38360 80888 38372
rect 80940 38400 80946 38412
rect 83737 38403 83795 38409
rect 83737 38400 83749 38403
rect 80940 38372 83749 38400
rect 80940 38360 80946 38372
rect 83737 38369 83749 38372
rect 83783 38369 83795 38403
rect 83737 38363 83795 38369
rect 84105 38403 84163 38409
rect 84105 38369 84117 38403
rect 84151 38400 84163 38403
rect 84396 38400 84424 38499
rect 84151 38372 84424 38400
rect 84151 38369 84163 38372
rect 84105 38363 84163 38369
rect 79042 38292 79048 38344
rect 79100 38341 79106 38344
rect 79100 38335 79158 38341
rect 79100 38301 79112 38335
rect 79146 38301 79158 38335
rect 79100 38295 79158 38301
rect 79321 38335 79379 38341
rect 79321 38301 79333 38335
rect 79367 38301 79379 38335
rect 79321 38295 79379 38301
rect 83645 38335 83703 38341
rect 83645 38301 83657 38335
rect 83691 38301 83703 38335
rect 84194 38332 84200 38344
rect 84155 38304 84200 38332
rect 83645 38295 83703 38301
rect 79100 38292 79106 38295
rect 78950 38264 78956 38276
rect 78600 38236 78956 38264
rect 73525 38227 73583 38233
rect 78950 38224 78956 38236
rect 79008 38264 79014 38276
rect 79229 38267 79287 38273
rect 79229 38264 79241 38267
rect 79008 38236 79241 38264
rect 79008 38224 79014 38236
rect 79229 38233 79241 38236
rect 79275 38233 79287 38267
rect 79229 38227 79287 38233
rect 62264 38168 65380 38196
rect 62264 38156 62270 38168
rect 65426 38156 65432 38208
rect 65484 38196 65490 38208
rect 78766 38196 78772 38208
rect 65484 38168 65529 38196
rect 78727 38168 78772 38196
rect 65484 38156 65490 38168
rect 78766 38156 78772 38168
rect 78824 38196 78830 38208
rect 79336 38196 79364 38295
rect 79410 38224 79416 38276
rect 79468 38264 79474 38276
rect 82909 38267 82967 38273
rect 82909 38264 82921 38267
rect 79468 38236 82921 38264
rect 79468 38224 79474 38236
rect 82909 38233 82921 38236
rect 82955 38264 82967 38267
rect 83660 38264 83688 38295
rect 84194 38292 84200 38304
rect 84252 38292 84258 38344
rect 85390 38264 85396 38276
rect 82955 38236 85396 38264
rect 82955 38233 82967 38236
rect 82909 38227 82967 38233
rect 85390 38224 85396 38236
rect 85448 38224 85454 38276
rect 78824 38168 79364 38196
rect 78824 38156 78830 38168
rect 79962 38156 79968 38208
rect 80020 38196 80026 38208
rect 83366 38196 83372 38208
rect 80020 38168 83372 38196
rect 80020 38156 80026 38168
rect 83366 38156 83372 38168
rect 83424 38156 83430 38208
rect 1104 38106 108008 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 65686 38106
rect 65738 38054 65750 38106
rect 65802 38054 65814 38106
rect 65866 38054 65878 38106
rect 65930 38054 96406 38106
rect 96458 38054 96470 38106
rect 96522 38054 96534 38106
rect 96586 38054 96598 38106
rect 96650 38054 108008 38106
rect 1104 38032 108008 38054
rect 4341 37995 4399 38001
rect 4341 37961 4353 37995
rect 4387 37992 4399 37995
rect 4614 37992 4620 38004
rect 4387 37964 4620 37992
rect 4387 37961 4399 37964
rect 4341 37955 4399 37961
rect 4614 37952 4620 37964
rect 4672 37952 4678 38004
rect 4706 37952 4712 38004
rect 4764 37992 4770 38004
rect 4893 37995 4951 38001
rect 4764 37964 4809 37992
rect 4764 37952 4770 37964
rect 4893 37961 4905 37995
rect 4939 37992 4951 37995
rect 5074 37992 5080 38004
rect 4939 37964 5080 37992
rect 4939 37961 4951 37964
rect 4893 37955 4951 37961
rect 5074 37952 5080 37964
rect 5132 37952 5138 38004
rect 10689 37995 10747 38001
rect 10689 37961 10701 37995
rect 10735 37992 10747 37995
rect 11054 37992 11060 38004
rect 10735 37964 11060 37992
rect 10735 37961 10747 37964
rect 10689 37955 10747 37961
rect 11054 37952 11060 37964
rect 11112 37952 11118 38004
rect 22186 37992 22192 38004
rect 22147 37964 22192 37992
rect 22186 37952 22192 37964
rect 22244 37952 22250 38004
rect 23661 37995 23719 38001
rect 23661 37961 23673 37995
rect 23707 37992 23719 37995
rect 51718 37992 51724 38004
rect 23707 37964 51724 37992
rect 23707 37961 23719 37964
rect 23661 37955 23719 37961
rect 51718 37952 51724 37964
rect 51776 37952 51782 38004
rect 52917 37995 52975 38001
rect 52917 37961 52929 37995
rect 52963 37992 52975 37995
rect 54570 37992 54576 38004
rect 52963 37964 54576 37992
rect 52963 37961 52975 37964
rect 52917 37955 52975 37961
rect 54570 37952 54576 37964
rect 54628 37952 54634 38004
rect 58710 37952 58716 38004
rect 58768 38001 58774 38004
rect 58768 37995 58817 38001
rect 58768 37961 58771 37995
rect 58805 37961 58817 37995
rect 58768 37955 58817 37961
rect 58768 37952 58774 37955
rect 58894 37952 58900 38004
rect 58952 37992 58958 38004
rect 58952 37964 58997 37992
rect 58952 37952 58958 37964
rect 60826 37952 60832 38004
rect 60884 37992 60890 38004
rect 70118 37992 70124 38004
rect 60884 37964 70124 37992
rect 60884 37952 60890 37964
rect 70118 37952 70124 37964
rect 70176 37952 70182 38004
rect 72237 37995 72295 38001
rect 72237 37961 72249 37995
rect 72283 37992 72295 37995
rect 72326 37992 72332 38004
rect 72283 37964 72332 37992
rect 72283 37961 72295 37964
rect 72237 37955 72295 37961
rect 72326 37952 72332 37964
rect 72384 37992 72390 38004
rect 73062 37992 73068 38004
rect 72384 37964 73068 37992
rect 72384 37952 72390 37964
rect 73062 37952 73068 37964
rect 73120 37952 73126 38004
rect 77478 37992 77484 38004
rect 77439 37964 77484 37992
rect 77478 37952 77484 37964
rect 77536 37952 77542 38004
rect 77754 37992 77760 38004
rect 77715 37964 77760 37992
rect 77754 37952 77760 37964
rect 77812 37952 77818 38004
rect 86681 37995 86739 38001
rect 86681 37961 86693 37995
rect 86727 37992 86739 37995
rect 86770 37992 86776 38004
rect 86727 37964 86776 37992
rect 86727 37961 86739 37964
rect 86681 37955 86739 37961
rect 86770 37952 86776 37964
rect 86828 37952 86834 38004
rect 4724 37924 4752 37952
rect 3528 37896 4752 37924
rect 3053 37859 3111 37865
rect 3053 37825 3065 37859
rect 3099 37856 3111 37859
rect 3237 37859 3295 37865
rect 3237 37856 3249 37859
rect 3099 37828 3249 37856
rect 3099 37825 3111 37828
rect 3053 37819 3111 37825
rect 3237 37825 3249 37828
rect 3283 37856 3295 37859
rect 3283 37828 3464 37856
rect 3283 37825 3295 37828
rect 3237 37819 3295 37825
rect 3436 37800 3464 37828
rect 3329 37791 3387 37797
rect 3329 37757 3341 37791
rect 3375 37757 3387 37791
rect 3329 37751 3387 37757
rect 3344 37720 3372 37751
rect 3418 37748 3424 37800
rect 3476 37748 3482 37800
rect 3528 37788 3556 37896
rect 15838 37884 15844 37936
rect 15896 37924 15902 37936
rect 16393 37927 16451 37933
rect 16393 37924 16405 37927
rect 15896 37896 16405 37924
rect 15896 37884 15902 37896
rect 16393 37893 16405 37896
rect 16439 37893 16451 37927
rect 21726 37924 21732 37936
rect 21687 37896 21732 37924
rect 16393 37887 16451 37893
rect 21726 37884 21732 37896
rect 21784 37884 21790 37936
rect 22646 37884 22652 37936
rect 22704 37924 22710 37936
rect 27614 37924 27620 37936
rect 22704 37896 27620 37924
rect 22704 37884 22710 37896
rect 27614 37884 27620 37896
rect 27672 37884 27678 37936
rect 29104 37896 36492 37924
rect 10962 37816 10968 37868
rect 11020 37856 11026 37868
rect 11057 37859 11115 37865
rect 11057 37856 11069 37859
rect 11020 37828 11069 37856
rect 11020 37816 11026 37828
rect 11057 37825 11069 37828
rect 11103 37856 11115 37859
rect 12526 37856 12532 37868
rect 11103 37828 12532 37856
rect 11103 37825 11115 37828
rect 11057 37819 11115 37825
rect 12526 37816 12532 37828
rect 12584 37816 12590 37868
rect 16022 37816 16028 37868
rect 16080 37856 16086 37868
rect 16080 37828 20852 37856
rect 16080 37816 16086 37828
rect 3789 37791 3847 37797
rect 3789 37788 3801 37791
rect 3528 37760 3801 37788
rect 3789 37757 3801 37760
rect 3835 37757 3847 37791
rect 3789 37751 3847 37757
rect 3881 37791 3939 37797
rect 3881 37757 3893 37791
rect 3927 37788 3939 37791
rect 5074 37788 5080 37800
rect 3927 37760 5080 37788
rect 3927 37757 3939 37760
rect 3881 37751 3939 37757
rect 3896 37720 3924 37751
rect 5074 37748 5080 37760
rect 5132 37748 5138 37800
rect 5626 37788 5632 37800
rect 5587 37760 5632 37788
rect 5626 37748 5632 37760
rect 5684 37748 5690 37800
rect 9493 37791 9551 37797
rect 9493 37788 9505 37791
rect 9324 37760 9505 37788
rect 5718 37720 5724 37732
rect 3344 37692 3924 37720
rect 5679 37692 5724 37720
rect 5718 37680 5724 37692
rect 5776 37680 5782 37732
rect 3786 37612 3792 37664
rect 3844 37652 3850 37664
rect 9324 37661 9352 37760
rect 9493 37757 9505 37760
rect 9539 37757 9551 37791
rect 9493 37751 9551 37757
rect 9677 37791 9735 37797
rect 9677 37757 9689 37791
rect 9723 37757 9735 37791
rect 10226 37788 10232 37800
rect 10187 37760 10232 37788
rect 9677 37751 9735 37757
rect 9692 37720 9720 37751
rect 10226 37748 10232 37760
rect 10284 37748 10290 37800
rect 10413 37791 10471 37797
rect 10413 37757 10425 37791
rect 10459 37788 10471 37791
rect 10980 37788 11008 37816
rect 10459 37760 11008 37788
rect 10459 37757 10471 37760
rect 10413 37751 10471 37757
rect 12434 37748 12440 37800
rect 12492 37788 12498 37800
rect 16117 37791 16175 37797
rect 12492 37760 12537 37788
rect 12492 37748 12498 37760
rect 16117 37757 16129 37791
rect 16163 37788 16175 37791
rect 16209 37791 16267 37797
rect 16209 37788 16221 37791
rect 16163 37760 16221 37788
rect 16163 37757 16175 37760
rect 16117 37751 16175 37757
rect 16209 37757 16221 37760
rect 16255 37757 16267 37791
rect 16209 37751 16267 37757
rect 20349 37791 20407 37797
rect 20349 37757 20361 37791
rect 20395 37788 20407 37791
rect 20625 37791 20683 37797
rect 20625 37788 20637 37791
rect 20395 37760 20637 37788
rect 20395 37757 20407 37760
rect 20349 37751 20407 37757
rect 20625 37757 20637 37760
rect 20671 37788 20683 37791
rect 20714 37788 20720 37800
rect 20671 37760 20720 37788
rect 20671 37757 20683 37760
rect 20625 37751 20683 37757
rect 20714 37748 20720 37760
rect 20772 37748 20778 37800
rect 20824 37797 20852 37828
rect 23658 37816 23664 37868
rect 23716 37856 23722 37868
rect 25317 37859 25375 37865
rect 25317 37856 25329 37859
rect 23716 37828 25329 37856
rect 23716 37816 23722 37828
rect 25317 37825 25329 37828
rect 25363 37856 25375 37859
rect 25498 37856 25504 37868
rect 25363 37828 25504 37856
rect 25363 37825 25375 37828
rect 25317 37819 25375 37825
rect 25498 37816 25504 37828
rect 25556 37816 25562 37868
rect 25590 37816 25596 37868
rect 25648 37856 25654 37868
rect 25648 37828 25820 37856
rect 25648 37816 25654 37828
rect 20809 37791 20867 37797
rect 20809 37757 20821 37791
rect 20855 37788 20867 37791
rect 21358 37788 21364 37800
rect 20855 37760 21364 37788
rect 20855 37757 20867 37760
rect 20809 37751 20867 37757
rect 21358 37748 21364 37760
rect 21416 37748 21422 37800
rect 21545 37791 21603 37797
rect 21545 37757 21557 37791
rect 21591 37788 21603 37791
rect 22186 37788 22192 37800
rect 21591 37760 22192 37788
rect 21591 37757 21603 37760
rect 21545 37751 21603 37757
rect 22186 37748 22192 37760
rect 22244 37748 22250 37800
rect 23937 37791 23995 37797
rect 23937 37757 23949 37791
rect 23983 37757 23995 37791
rect 25685 37791 25743 37797
rect 25685 37788 25697 37791
rect 23937 37751 23995 37757
rect 24136 37760 25697 37788
rect 10244 37720 10272 37748
rect 9692 37692 10272 37720
rect 10502 37680 10508 37732
rect 10560 37720 10566 37732
rect 23661 37723 23719 37729
rect 23661 37720 23673 37723
rect 10560 37692 23673 37720
rect 10560 37680 10566 37692
rect 23661 37689 23673 37692
rect 23707 37689 23719 37723
rect 23661 37683 23719 37689
rect 23750 37680 23756 37732
rect 23808 37720 23814 37732
rect 23952 37720 23980 37751
rect 23808 37692 23980 37720
rect 23808 37680 23814 37692
rect 9309 37655 9367 37661
rect 9309 37652 9321 37655
rect 3844 37624 9321 37652
rect 3844 37612 3850 37624
rect 9309 37621 9321 37624
rect 9355 37621 9367 37655
rect 9309 37615 9367 37621
rect 16117 37655 16175 37661
rect 16117 37621 16129 37655
rect 16163 37652 16175 37655
rect 16669 37655 16727 37661
rect 16669 37652 16681 37655
rect 16163 37624 16681 37652
rect 16163 37621 16175 37624
rect 16117 37615 16175 37621
rect 16669 37621 16681 37624
rect 16715 37652 16727 37655
rect 17310 37652 17316 37664
rect 16715 37624 17316 37652
rect 16715 37621 16727 37624
rect 16669 37615 16727 37621
rect 17310 37612 17316 37624
rect 17368 37652 17374 37664
rect 17862 37652 17868 37664
rect 17368 37624 17868 37652
rect 17368 37612 17374 37624
rect 17862 37612 17868 37624
rect 17920 37612 17926 37664
rect 20070 37612 20076 37664
rect 20128 37652 20134 37664
rect 20349 37655 20407 37661
rect 20349 37652 20361 37655
rect 20128 37624 20361 37652
rect 20128 37612 20134 37624
rect 20349 37621 20361 37624
rect 20395 37652 20407 37655
rect 20441 37655 20499 37661
rect 20441 37652 20453 37655
rect 20395 37624 20453 37652
rect 20395 37621 20407 37624
rect 20349 37615 20407 37621
rect 20441 37621 20453 37624
rect 20487 37621 20499 37655
rect 20441 37615 20499 37621
rect 21358 37612 21364 37664
rect 21416 37652 21422 37664
rect 24136 37661 24164 37760
rect 25685 37757 25697 37760
rect 25731 37757 25743 37791
rect 25792 37788 25820 37828
rect 26142 37788 26148 37800
rect 25792 37760 26148 37788
rect 25685 37751 25743 37757
rect 25700 37720 25728 37751
rect 26142 37748 26148 37760
rect 26200 37748 26206 37800
rect 26237 37791 26295 37797
rect 26237 37757 26249 37791
rect 26283 37757 26295 37791
rect 26237 37751 26295 37757
rect 26252 37720 26280 37751
rect 27706 37748 27712 37800
rect 27764 37788 27770 37800
rect 29104 37788 29132 37896
rect 36354 37856 36360 37868
rect 33152 37828 36360 37856
rect 33152 37797 33180 37828
rect 36354 37816 36360 37828
rect 36412 37816 36418 37868
rect 27764 37760 29132 37788
rect 33137 37791 33195 37797
rect 27764 37748 27770 37760
rect 33137 37757 33149 37791
rect 33183 37757 33195 37791
rect 33137 37751 33195 37757
rect 33597 37791 33655 37797
rect 33597 37757 33609 37791
rect 33643 37788 33655 37791
rect 34606 37788 34612 37800
rect 33643 37760 34612 37788
rect 33643 37757 33655 37760
rect 33597 37751 33655 37757
rect 34606 37748 34612 37760
rect 34664 37748 34670 37800
rect 34790 37748 34796 37800
rect 34848 37788 34854 37800
rect 34885 37791 34943 37797
rect 34885 37788 34897 37791
rect 34848 37760 34897 37788
rect 34848 37748 34854 37760
rect 34885 37757 34897 37760
rect 34931 37757 34943 37791
rect 36464 37788 36492 37896
rect 36630 37884 36636 37936
rect 36688 37924 36694 37936
rect 38979 37927 39037 37933
rect 38979 37924 38991 37927
rect 36688 37896 38991 37924
rect 36688 37884 36694 37896
rect 38979 37893 38991 37896
rect 39025 37893 39037 37927
rect 38979 37887 39037 37893
rect 39117 37927 39175 37933
rect 39117 37893 39129 37927
rect 39163 37893 39175 37927
rect 51442 37924 51448 37936
rect 39117 37887 39175 37893
rect 39960 37896 51448 37924
rect 37274 37816 37280 37868
rect 37332 37856 37338 37868
rect 39132 37856 39160 37887
rect 37332 37828 39160 37856
rect 39209 37859 39267 37865
rect 37332 37816 37338 37828
rect 39209 37825 39221 37859
rect 39255 37856 39267 37859
rect 39850 37856 39856 37868
rect 39255 37828 39856 37856
rect 39255 37825 39267 37828
rect 39209 37819 39267 37825
rect 39850 37816 39856 37828
rect 39908 37816 39914 37868
rect 39960 37788 39988 37896
rect 51442 37884 51448 37896
rect 51500 37884 51506 37936
rect 52362 37884 52368 37936
rect 52420 37924 52426 37936
rect 58437 37927 58495 37933
rect 58437 37924 58449 37927
rect 52420 37896 58449 37924
rect 52420 37884 52426 37896
rect 58437 37893 58449 37896
rect 58483 37924 58495 37927
rect 58618 37924 58624 37936
rect 58483 37896 58624 37924
rect 58483 37893 58495 37896
rect 58437 37887 58495 37893
rect 58618 37884 58624 37896
rect 58676 37884 58682 37936
rect 81345 37927 81403 37933
rect 81345 37924 81357 37927
rect 58912 37896 81357 37924
rect 53285 37859 53343 37865
rect 53285 37825 53297 37859
rect 53331 37856 53343 37859
rect 53374 37856 53380 37868
rect 53331 37828 53380 37856
rect 53331 37825 53343 37828
rect 53285 37819 53343 37825
rect 36464 37760 39988 37788
rect 46109 37791 46167 37797
rect 34885 37751 34943 37757
rect 46109 37757 46121 37791
rect 46155 37788 46167 37791
rect 46566 37788 46572 37800
rect 46155 37760 46572 37788
rect 46155 37757 46167 37760
rect 46109 37751 46167 37757
rect 46566 37748 46572 37760
rect 46624 37788 46630 37800
rect 51721 37791 51779 37797
rect 51721 37788 51733 37791
rect 46624 37760 51733 37788
rect 46624 37748 46630 37760
rect 51721 37757 51733 37760
rect 51767 37757 51779 37791
rect 51721 37751 51779 37757
rect 51905 37791 51963 37797
rect 51905 37757 51917 37791
rect 51951 37788 51963 37791
rect 51994 37788 52000 37800
rect 51951 37760 52000 37788
rect 51951 37757 51963 37760
rect 51905 37751 51963 37757
rect 51994 37748 52000 37760
rect 52052 37748 52058 37800
rect 52362 37788 52368 37800
rect 52323 37760 52368 37788
rect 52362 37748 52368 37760
rect 52420 37748 52426 37800
rect 52457 37791 52515 37797
rect 52457 37757 52469 37791
rect 52503 37788 52515 37791
rect 52546 37788 52552 37800
rect 52503 37760 52552 37788
rect 52503 37757 52515 37760
rect 52457 37751 52515 37757
rect 52546 37748 52552 37760
rect 52604 37788 52610 37800
rect 53300 37788 53328 37819
rect 53374 37816 53380 37828
rect 53432 37856 53438 37868
rect 58912 37856 58940 37896
rect 81345 37893 81357 37896
rect 81391 37924 81403 37927
rect 85574 37924 85580 37936
rect 81391 37896 85580 37924
rect 81391 37893 81403 37896
rect 81345 37887 81403 37893
rect 85574 37884 85580 37896
rect 85632 37884 85638 37936
rect 53432 37828 58940 37856
rect 58986 37859 59044 37865
rect 53432 37816 53438 37828
rect 58986 37825 58998 37859
rect 59032 37856 59044 37859
rect 59032 37828 64092 37856
rect 59032 37825 59044 37828
rect 58986 37819 59044 37825
rect 52604 37760 53328 37788
rect 53469 37791 53527 37797
rect 52604 37748 52610 37760
rect 53469 37757 53481 37791
rect 53515 37788 53527 37791
rect 53558 37788 53564 37800
rect 53515 37760 53564 37788
rect 53515 37757 53527 37760
rect 53469 37751 53527 37757
rect 53558 37748 53564 37760
rect 53616 37788 53622 37800
rect 55030 37788 55036 37800
rect 53616 37760 55036 37788
rect 53616 37748 53622 37760
rect 55030 37748 55036 37760
rect 55088 37748 55094 37800
rect 55876 37760 60964 37788
rect 25700 37692 26280 37720
rect 26789 37723 26847 37729
rect 26789 37689 26801 37723
rect 26835 37720 26847 37723
rect 27154 37720 27160 37732
rect 26835 37692 27160 37720
rect 26835 37689 26847 37692
rect 26789 37683 26847 37689
rect 27154 37680 27160 37692
rect 27212 37680 27218 37732
rect 38838 37720 38844 37732
rect 32232 37692 35112 37720
rect 38799 37692 38844 37720
rect 24121 37655 24179 37661
rect 24121 37652 24133 37655
rect 21416 37624 24133 37652
rect 21416 37612 21422 37624
rect 24121 37621 24133 37624
rect 24167 37621 24179 37655
rect 24121 37615 24179 37621
rect 26142 37612 26148 37664
rect 26200 37652 26206 37664
rect 26973 37655 27031 37661
rect 26973 37652 26985 37655
rect 26200 37624 26985 37652
rect 26200 37612 26206 37624
rect 26973 37621 26985 37624
rect 27019 37652 27031 37655
rect 32232 37652 32260 37692
rect 27019 37624 32260 37652
rect 27019 37621 27031 37624
rect 26973 37615 27031 37621
rect 32306 37612 32312 37664
rect 32364 37652 32370 37664
rect 32950 37652 32956 37664
rect 32364 37624 32956 37652
rect 32364 37612 32370 37624
rect 32950 37612 32956 37624
rect 33008 37612 33014 37664
rect 33686 37652 33692 37664
rect 33647 37624 33692 37652
rect 33686 37612 33692 37624
rect 33744 37612 33750 37664
rect 34974 37652 34980 37664
rect 34935 37624 34980 37652
rect 34974 37612 34980 37624
rect 35032 37612 35038 37664
rect 35084 37652 35112 37692
rect 38838 37680 38844 37692
rect 38896 37680 38902 37732
rect 39577 37723 39635 37729
rect 39577 37689 39589 37723
rect 39623 37720 39635 37723
rect 46014 37720 46020 37732
rect 39623 37692 46020 37720
rect 39623 37689 39635 37692
rect 39577 37683 39635 37689
rect 46014 37680 46020 37692
rect 46072 37680 46078 37732
rect 55876 37720 55904 37760
rect 46124 37692 55904 37720
rect 46124 37652 46152 37692
rect 56502 37680 56508 37732
rect 56560 37720 56566 37732
rect 58621 37723 58679 37729
rect 58621 37720 58633 37723
rect 56560 37692 58633 37720
rect 56560 37680 56566 37692
rect 58621 37689 58633 37692
rect 58667 37689 58679 37723
rect 60936 37720 60964 37760
rect 61010 37748 61016 37800
rect 61068 37788 61074 37800
rect 61105 37791 61163 37797
rect 61105 37788 61117 37791
rect 61068 37760 61117 37788
rect 61068 37748 61074 37760
rect 61105 37757 61117 37760
rect 61151 37757 61163 37791
rect 61105 37751 61163 37757
rect 63310 37748 63316 37800
rect 63368 37788 63374 37800
rect 63497 37791 63555 37797
rect 63497 37788 63509 37791
rect 63368 37760 63509 37788
rect 63368 37748 63374 37760
rect 63497 37757 63509 37760
rect 63543 37757 63555 37791
rect 64064 37788 64092 37828
rect 64690 37816 64696 37868
rect 64748 37856 64754 37868
rect 65429 37859 65487 37865
rect 65429 37856 65441 37859
rect 64748 37828 65441 37856
rect 64748 37816 64754 37828
rect 65429 37825 65441 37828
rect 65475 37825 65487 37859
rect 65429 37819 65487 37825
rect 79870 37816 79876 37868
rect 79928 37856 79934 37868
rect 79928 37828 81204 37856
rect 79928 37816 79934 37828
rect 64874 37788 64880 37800
rect 64064 37760 64880 37788
rect 63497 37751 63555 37757
rect 64874 37748 64880 37760
rect 64932 37748 64938 37800
rect 64969 37791 65027 37797
rect 64969 37757 64981 37791
rect 65015 37757 65027 37791
rect 65150 37788 65156 37800
rect 65111 37760 65156 37788
rect 64969 37751 65027 37757
rect 63589 37723 63647 37729
rect 63589 37720 63601 37723
rect 60936 37692 63601 37720
rect 58621 37683 58679 37689
rect 63589 37689 63601 37692
rect 63635 37720 63647 37723
rect 64325 37723 64383 37729
rect 64325 37720 64337 37723
rect 63635 37692 64337 37720
rect 63635 37689 63647 37692
rect 63589 37683 63647 37689
rect 64325 37689 64337 37692
rect 64371 37720 64383 37723
rect 64984 37720 65012 37751
rect 65150 37748 65156 37760
rect 65208 37748 65214 37800
rect 65518 37788 65524 37800
rect 65479 37760 65524 37788
rect 65518 37748 65524 37760
rect 65576 37748 65582 37800
rect 72326 37788 72332 37800
rect 72287 37760 72332 37788
rect 72326 37748 72332 37760
rect 72384 37748 72390 37800
rect 72436 37760 73108 37788
rect 64371 37692 65012 37720
rect 64371 37689 64383 37692
rect 64325 37683 64383 37689
rect 65058 37680 65064 37732
rect 65116 37720 65122 37732
rect 66438 37720 66444 37732
rect 65116 37692 66444 37720
rect 65116 37680 65122 37692
rect 66438 37680 66444 37692
rect 66496 37680 66502 37732
rect 68554 37680 68560 37732
rect 68612 37720 68618 37732
rect 72436 37720 72464 37760
rect 68612 37692 72464 37720
rect 73080 37720 73108 37760
rect 73154 37748 73160 37800
rect 73212 37788 73218 37800
rect 74169 37791 74227 37797
rect 74169 37788 74181 37791
rect 73212 37760 74181 37788
rect 73212 37748 73218 37760
rect 74169 37757 74181 37760
rect 74215 37757 74227 37791
rect 74169 37751 74227 37757
rect 77389 37791 77447 37797
rect 77389 37757 77401 37791
rect 77435 37788 77447 37791
rect 77754 37788 77760 37800
rect 77435 37760 77760 37788
rect 77435 37757 77447 37760
rect 77389 37751 77447 37757
rect 77754 37748 77760 37760
rect 77812 37748 77818 37800
rect 79778 37788 79784 37800
rect 79739 37760 79784 37788
rect 79778 37748 79784 37760
rect 79836 37748 79842 37800
rect 79962 37788 79968 37800
rect 79923 37760 79968 37788
rect 79962 37748 79968 37760
rect 80020 37788 80026 37800
rect 81176 37797 81204 37828
rect 80425 37791 80483 37797
rect 80425 37788 80437 37791
rect 80020 37760 80437 37788
rect 80020 37748 80026 37760
rect 80425 37757 80437 37760
rect 80471 37757 80483 37791
rect 80425 37751 80483 37757
rect 81161 37791 81219 37797
rect 81161 37757 81173 37791
rect 81207 37757 81219 37791
rect 86586 37788 86592 37800
rect 86547 37760 86592 37788
rect 81161 37751 81219 37757
rect 86586 37748 86592 37760
rect 86644 37748 86650 37800
rect 79318 37720 79324 37732
rect 73080 37692 79324 37720
rect 68612 37680 68618 37692
rect 79318 37680 79324 37692
rect 79376 37680 79382 37732
rect 79796 37720 79824 37748
rect 80330 37720 80336 37732
rect 79796 37692 80192 37720
rect 80291 37692 80336 37720
rect 35084 37624 46152 37652
rect 46198 37612 46204 37664
rect 46256 37652 46262 37664
rect 46256 37624 46301 37652
rect 46256 37612 46262 37624
rect 51994 37612 52000 37664
rect 52052 37652 52058 37664
rect 53558 37652 53564 37664
rect 52052 37624 53564 37652
rect 52052 37612 52058 37624
rect 53558 37612 53564 37624
rect 53616 37612 53622 37664
rect 59265 37655 59323 37661
rect 59265 37621 59277 37655
rect 59311 37652 59323 37655
rect 60182 37652 60188 37664
rect 59311 37624 60188 37652
rect 59311 37621 59323 37624
rect 59265 37615 59323 37621
rect 60182 37612 60188 37624
rect 60240 37612 60246 37664
rect 60918 37652 60924 37664
rect 60831 37624 60924 37652
rect 60918 37612 60924 37624
rect 60976 37652 60982 37664
rect 63126 37652 63132 37664
rect 60976 37624 63132 37652
rect 60976 37612 60982 37624
rect 63126 37612 63132 37624
rect 63184 37612 63190 37664
rect 63310 37652 63316 37664
rect 63271 37624 63316 37652
rect 63310 37612 63316 37624
rect 63368 37652 63374 37664
rect 64141 37655 64199 37661
rect 64141 37652 64153 37655
rect 63368 37624 64153 37652
rect 63368 37612 63374 37624
rect 64141 37621 64153 37624
rect 64187 37652 64199 37655
rect 64690 37652 64696 37664
rect 64187 37624 64696 37652
rect 64187 37621 64199 37624
rect 64141 37615 64199 37621
rect 64690 37612 64696 37624
rect 64748 37612 64754 37664
rect 64785 37655 64843 37661
rect 64785 37621 64797 37655
rect 64831 37652 64843 37655
rect 66162 37652 66168 37664
rect 64831 37624 66168 37652
rect 64831 37621 64843 37624
rect 64785 37615 64843 37621
rect 66162 37612 66168 37624
rect 66220 37612 66226 37664
rect 72510 37652 72516 37664
rect 72471 37624 72516 37652
rect 72510 37612 72516 37624
rect 72568 37612 72574 37664
rect 72602 37612 72608 37664
rect 72660 37652 72666 37664
rect 74353 37655 74411 37661
rect 74353 37652 74365 37655
rect 72660 37624 74365 37652
rect 72660 37612 72666 37624
rect 74353 37621 74365 37624
rect 74399 37652 74411 37655
rect 79410 37652 79416 37664
rect 74399 37624 79416 37652
rect 74399 37621 74411 37624
rect 74353 37615 74411 37621
rect 79410 37612 79416 37624
rect 79468 37612 79474 37664
rect 80164 37652 80192 37692
rect 80330 37680 80336 37692
rect 80388 37680 80394 37732
rect 84194 37652 84200 37664
rect 80164 37624 84200 37652
rect 84194 37612 84200 37624
rect 84252 37612 84258 37664
rect 1104 37562 108008 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 81046 37562
rect 81098 37510 81110 37562
rect 81162 37510 81174 37562
rect 81226 37510 81238 37562
rect 81290 37510 108008 37562
rect 1104 37488 108008 37510
rect 4798 37448 4804 37460
rect 4172 37420 4804 37448
rect 4172 37321 4200 37420
rect 4798 37408 4804 37420
rect 4856 37448 4862 37460
rect 5537 37451 5595 37457
rect 4856 37420 5304 37448
rect 4856 37408 4862 37420
rect 5276 37380 5304 37420
rect 5537 37417 5549 37451
rect 5583 37448 5595 37451
rect 5626 37448 5632 37460
rect 5583 37420 5632 37448
rect 5583 37417 5595 37420
rect 5537 37411 5595 37417
rect 5626 37408 5632 37420
rect 5684 37408 5690 37460
rect 10962 37448 10968 37460
rect 10923 37420 10968 37448
rect 10962 37408 10968 37420
rect 11020 37408 11026 37460
rect 11054 37408 11060 37460
rect 11112 37448 11118 37460
rect 11241 37451 11299 37457
rect 11241 37448 11253 37451
rect 11112 37420 11253 37448
rect 11112 37408 11118 37420
rect 11241 37417 11253 37420
rect 11287 37448 11299 37451
rect 11287 37420 21036 37448
rect 11287 37417 11299 37420
rect 11241 37411 11299 37417
rect 5905 37383 5963 37389
rect 5905 37380 5917 37383
rect 5276 37352 5917 37380
rect 5905 37349 5917 37352
rect 5951 37349 5963 37383
rect 5905 37343 5963 37349
rect 5994 37340 6000 37392
rect 6052 37380 6058 37392
rect 20901 37383 20959 37389
rect 20901 37380 20913 37383
rect 6052 37352 11008 37380
rect 6052 37340 6058 37352
rect 4157 37315 4215 37321
rect 4157 37281 4169 37315
rect 4203 37281 4215 37315
rect 4157 37275 4215 37281
rect 5718 37272 5724 37324
rect 5776 37312 5782 37324
rect 9493 37315 9551 37321
rect 9493 37312 9505 37315
rect 5776 37284 9505 37312
rect 5776 37272 5782 37284
rect 9493 37281 9505 37284
rect 9539 37312 9551 37315
rect 10318 37312 10324 37324
rect 9539 37284 10180 37312
rect 10279 37284 10324 37312
rect 9539 37281 9551 37284
rect 9493 37275 9551 37281
rect 4433 37247 4491 37253
rect 4433 37213 4445 37247
rect 4479 37244 4491 37247
rect 4798 37244 4804 37256
rect 4479 37216 4804 37244
rect 4479 37213 4491 37216
rect 4433 37207 4491 37213
rect 4798 37204 4804 37216
rect 4856 37204 4862 37256
rect 9674 37244 9680 37256
rect 9635 37216 9680 37244
rect 9674 37204 9680 37216
rect 9732 37204 9738 37256
rect 10152 37244 10180 37284
rect 10318 37272 10324 37284
rect 10376 37272 10382 37324
rect 10689 37315 10747 37321
rect 10689 37281 10701 37315
rect 10735 37281 10747 37315
rect 10870 37312 10876 37324
rect 10831 37284 10876 37312
rect 10689 37275 10747 37281
rect 10413 37247 10471 37253
rect 10413 37244 10425 37247
rect 10152 37216 10425 37244
rect 10413 37213 10425 37216
rect 10459 37244 10471 37247
rect 10502 37244 10508 37256
rect 10459 37216 10508 37244
rect 10459 37213 10471 37216
rect 10413 37207 10471 37213
rect 10502 37204 10508 37216
rect 10560 37204 10566 37256
rect 10704 37244 10732 37275
rect 10870 37272 10876 37284
rect 10928 37272 10934 37324
rect 10980 37312 11008 37352
rect 11164 37352 20913 37380
rect 11164 37312 11192 37352
rect 20901 37349 20913 37352
rect 20947 37349 20959 37383
rect 20901 37343 20959 37349
rect 10980 37284 11192 37312
rect 15289 37315 15347 37321
rect 15289 37281 15301 37315
rect 15335 37312 15347 37315
rect 15473 37315 15531 37321
rect 15335 37284 15424 37312
rect 15335 37281 15347 37284
rect 15289 37275 15347 37281
rect 11054 37244 11060 37256
rect 10704 37216 11060 37244
rect 11054 37204 11060 37216
rect 11112 37204 11118 37256
rect 15396 37244 15424 37284
rect 15473 37281 15485 37315
rect 15519 37312 15531 37315
rect 15562 37312 15568 37324
rect 15519 37284 15568 37312
rect 15519 37281 15531 37284
rect 15473 37275 15531 37281
rect 15562 37272 15568 37284
rect 15620 37272 15626 37324
rect 16025 37315 16083 37321
rect 16025 37312 16037 37315
rect 15672 37284 16037 37312
rect 15672 37244 15700 37284
rect 16025 37281 16037 37284
rect 16071 37312 16083 37315
rect 16114 37312 16120 37324
rect 16071 37284 16120 37312
rect 16071 37281 16083 37284
rect 16025 37275 16083 37281
rect 16114 37272 16120 37284
rect 16172 37272 16178 37324
rect 17126 37272 17132 37324
rect 17184 37312 17190 37324
rect 20717 37315 20775 37321
rect 20717 37312 20729 37315
rect 17184 37284 20729 37312
rect 17184 37272 17190 37284
rect 20717 37281 20729 37284
rect 20763 37281 20775 37315
rect 20717 37275 20775 37281
rect 20806 37272 20812 37324
rect 20864 37272 20870 37324
rect 15396 37216 15700 37244
rect 20533 37179 20591 37185
rect 20533 37145 20545 37179
rect 20579 37176 20591 37179
rect 20824 37176 20852 37272
rect 21008 37244 21036 37420
rect 30374 37408 30380 37460
rect 30432 37448 30438 37460
rect 32858 37448 32864 37460
rect 30432 37420 32864 37448
rect 30432 37408 30438 37420
rect 32858 37408 32864 37420
rect 32916 37408 32922 37460
rect 63310 37448 63316 37460
rect 32968 37420 63316 37448
rect 22186 37380 22192 37392
rect 21376 37352 22192 37380
rect 21376 37321 21404 37352
rect 22186 37340 22192 37352
rect 22244 37340 22250 37392
rect 22281 37383 22339 37389
rect 22281 37349 22293 37383
rect 22327 37380 22339 37383
rect 22738 37380 22744 37392
rect 22327 37352 22744 37380
rect 22327 37349 22339 37352
rect 22281 37343 22339 37349
rect 21361 37315 21419 37321
rect 21361 37281 21373 37315
rect 21407 37281 21419 37315
rect 21361 37275 21419 37281
rect 21450 37272 21456 37324
rect 21508 37312 21514 37324
rect 21545 37315 21603 37321
rect 21545 37312 21557 37315
rect 21508 37284 21557 37312
rect 21508 37272 21514 37284
rect 21545 37281 21557 37284
rect 21591 37281 21603 37315
rect 21545 37275 21603 37281
rect 21913 37315 21971 37321
rect 21913 37281 21925 37315
rect 21959 37312 21971 37315
rect 22097 37315 22155 37321
rect 21959 37284 21993 37312
rect 21959 37281 21971 37284
rect 21913 37275 21971 37281
rect 22097 37281 22109 37315
rect 22143 37312 22155 37315
rect 22296 37312 22324 37343
rect 22738 37340 22744 37352
rect 22796 37340 22802 37392
rect 28537 37383 28595 37389
rect 28537 37349 28549 37383
rect 28583 37380 28595 37383
rect 32968 37380 32996 37420
rect 63310 37408 63316 37420
rect 63368 37408 63374 37460
rect 63957 37451 64015 37457
rect 63957 37417 63969 37451
rect 64003 37448 64015 37451
rect 66070 37448 66076 37460
rect 64003 37420 66076 37448
rect 64003 37417 64015 37420
rect 63957 37411 64015 37417
rect 66070 37408 66076 37420
rect 66128 37408 66134 37460
rect 66254 37448 66260 37460
rect 66215 37420 66260 37448
rect 66254 37408 66260 37420
rect 66312 37408 66318 37460
rect 71682 37408 71688 37460
rect 71740 37448 71746 37460
rect 72421 37451 72479 37457
rect 72421 37448 72433 37451
rect 71740 37420 72433 37448
rect 71740 37408 71746 37420
rect 72421 37417 72433 37420
rect 72467 37417 72479 37451
rect 72421 37411 72479 37417
rect 73525 37451 73583 37457
rect 73525 37417 73537 37451
rect 73571 37448 73583 37451
rect 73614 37448 73620 37460
rect 73571 37420 73620 37448
rect 73571 37417 73583 37420
rect 73525 37411 73583 37417
rect 73614 37408 73620 37420
rect 73672 37408 73678 37460
rect 78950 37448 78956 37460
rect 78911 37420 78956 37448
rect 78950 37408 78956 37420
rect 79008 37408 79014 37460
rect 80164 37420 84148 37448
rect 33410 37380 33416 37392
rect 28583 37352 32996 37380
rect 33371 37352 33416 37380
rect 28583 37349 28595 37352
rect 28537 37343 28595 37349
rect 33410 37340 33416 37352
rect 33468 37340 33474 37392
rect 33689 37383 33747 37389
rect 33689 37349 33701 37383
rect 33735 37380 33747 37383
rect 34974 37380 34980 37392
rect 33735 37352 34980 37380
rect 33735 37349 33747 37352
rect 33689 37343 33747 37349
rect 22143 37284 22324 37312
rect 22143 37281 22155 37284
rect 22097 37275 22155 37281
rect 21818 37244 21824 37256
rect 21008 37216 21824 37244
rect 21818 37204 21824 37216
rect 21876 37244 21882 37256
rect 21928 37244 21956 37275
rect 22370 37272 22376 37324
rect 22428 37312 22434 37324
rect 27154 37312 27160 37324
rect 22428 37284 22473 37312
rect 27115 37284 27160 37312
rect 22428 37272 22434 37284
rect 27154 37272 27160 37284
rect 27212 37272 27218 37324
rect 32309 37315 32367 37321
rect 32309 37281 32321 37315
rect 32355 37312 32367 37315
rect 32861 37315 32919 37321
rect 32861 37312 32873 37315
rect 32355 37284 32873 37312
rect 32355 37281 32367 37284
rect 32309 37275 32367 37281
rect 32861 37281 32873 37284
rect 32907 37312 32919 37315
rect 32950 37312 32956 37324
rect 32907 37284 32956 37312
rect 32907 37281 32919 37284
rect 32861 37275 32919 37281
rect 32950 37272 32956 37284
rect 33008 37272 33014 37324
rect 33042 37272 33048 37324
rect 33100 37312 33106 37324
rect 33704 37312 33732 37343
rect 34974 37340 34980 37352
rect 35032 37340 35038 37392
rect 38286 37380 38292 37392
rect 38247 37352 38292 37380
rect 38286 37340 38292 37352
rect 38344 37340 38350 37392
rect 46566 37380 46572 37392
rect 46527 37352 46572 37380
rect 46566 37340 46572 37352
rect 46624 37340 46630 37392
rect 46658 37340 46664 37392
rect 46716 37380 46722 37392
rect 50982 37380 50988 37392
rect 46716 37352 50988 37380
rect 46716 37340 46722 37352
rect 50982 37340 50988 37352
rect 51040 37340 51046 37392
rect 53098 37380 53104 37392
rect 53059 37352 53104 37380
rect 53098 37340 53104 37352
rect 53156 37340 53162 37392
rect 53374 37380 53380 37392
rect 53335 37352 53380 37380
rect 53374 37340 53380 37352
rect 53432 37340 53438 37392
rect 53558 37380 53564 37392
rect 53519 37352 53564 37380
rect 53558 37340 53564 37352
rect 53616 37340 53622 37392
rect 59722 37340 59728 37392
rect 59780 37380 59786 37392
rect 60277 37383 60335 37389
rect 60277 37380 60289 37383
rect 59780 37352 60289 37380
rect 59780 37340 59786 37352
rect 60277 37349 60289 37352
rect 60323 37349 60335 37383
rect 60277 37343 60335 37349
rect 63126 37340 63132 37392
rect 63184 37380 63190 37392
rect 66990 37380 66996 37392
rect 63184 37352 64828 37380
rect 63184 37340 63190 37352
rect 34330 37312 34336 37324
rect 33100 37284 33732 37312
rect 34291 37284 34336 37312
rect 33100 37272 33106 37284
rect 34330 37272 34336 37284
rect 34388 37272 34394 37324
rect 40129 37315 40187 37321
rect 34532 37284 40080 37312
rect 22557 37247 22615 37253
rect 22557 37244 22569 37247
rect 21876 37216 22569 37244
rect 21876 37204 21882 37216
rect 22557 37213 22569 37216
rect 22603 37213 22615 37247
rect 22557 37207 22615 37213
rect 26786 37204 26792 37256
rect 26844 37244 26850 37256
rect 26881 37247 26939 37253
rect 26881 37244 26893 37247
rect 26844 37216 26893 37244
rect 26844 37204 26850 37216
rect 26881 37213 26893 37216
rect 26927 37244 26939 37247
rect 27890 37244 27896 37256
rect 26927 37216 27896 37244
rect 26927 37213 26939 37216
rect 26881 37207 26939 37213
rect 27890 37204 27896 37216
rect 27948 37244 27954 37256
rect 28629 37247 28687 37253
rect 28629 37244 28641 37247
rect 27948 37216 28641 37244
rect 27948 37204 27954 37216
rect 28629 37213 28641 37216
rect 28675 37213 28687 37247
rect 28629 37207 28687 37213
rect 32125 37247 32183 37253
rect 32125 37213 32137 37247
rect 32171 37213 32183 37247
rect 32125 37207 32183 37213
rect 20579 37148 20852 37176
rect 20579 37145 20591 37148
rect 20533 37139 20591 37145
rect 4062 37068 4068 37120
rect 4120 37108 4126 37120
rect 7926 37108 7932 37120
rect 4120 37080 7932 37108
rect 4120 37068 4126 37080
rect 7926 37068 7932 37080
rect 7984 37068 7990 37120
rect 14274 37068 14280 37120
rect 14332 37108 14338 37120
rect 15565 37111 15623 37117
rect 15565 37108 15577 37111
rect 14332 37080 15577 37108
rect 14332 37068 14338 37080
rect 15565 37077 15577 37080
rect 15611 37077 15623 37111
rect 15565 37071 15623 37077
rect 31941 37111 31999 37117
rect 31941 37077 31953 37111
rect 31987 37108 31999 37111
rect 32140 37108 32168 37207
rect 32950 37136 32956 37188
rect 33008 37176 33014 37188
rect 34532 37185 34560 37284
rect 38470 37244 38476 37256
rect 38431 37216 38476 37244
rect 38470 37204 38476 37216
rect 38528 37204 38534 37256
rect 38746 37244 38752 37256
rect 38707 37216 38752 37244
rect 38746 37204 38752 37216
rect 38804 37204 38810 37256
rect 40052 37244 40080 37284
rect 40129 37281 40141 37315
rect 40175 37312 40187 37315
rect 40954 37312 40960 37324
rect 40175 37284 40960 37312
rect 40175 37281 40187 37284
rect 40129 37275 40187 37281
rect 40954 37272 40960 37284
rect 41012 37272 41018 37324
rect 44542 37312 44548 37324
rect 44503 37284 44548 37312
rect 44542 37272 44548 37284
rect 44600 37272 44606 37324
rect 44818 37272 44824 37324
rect 44876 37321 44882 37324
rect 44876 37312 44887 37321
rect 51810 37312 51816 37324
rect 44876 37284 44921 37312
rect 51771 37284 51816 37312
rect 44876 37275 44887 37284
rect 44876 37272 44882 37275
rect 51810 37272 51816 37284
rect 51868 37272 51874 37324
rect 51994 37312 52000 37324
rect 51955 37284 52000 37312
rect 51994 37272 52000 37284
rect 52052 37272 52058 37324
rect 52546 37312 52552 37324
rect 52507 37284 52552 37312
rect 52546 37272 52552 37284
rect 52604 37272 52610 37324
rect 52733 37315 52791 37321
rect 52733 37281 52745 37315
rect 52779 37312 52791 37315
rect 60182 37312 60188 37324
rect 52779 37284 53144 37312
rect 60143 37284 60188 37312
rect 52779 37281 52791 37284
rect 52733 37275 52791 37281
rect 53116 37256 53144 37284
rect 60182 37272 60188 37284
rect 60240 37272 60246 37324
rect 64325 37315 64383 37321
rect 64325 37281 64337 37315
rect 64371 37312 64383 37315
rect 64598 37312 64604 37324
rect 64371 37284 64604 37312
rect 64371 37281 64383 37284
rect 64325 37275 64383 37281
rect 64598 37272 64604 37284
rect 64656 37272 64662 37324
rect 64800 37321 64828 37352
rect 65812 37352 66996 37380
rect 64693 37315 64751 37321
rect 64693 37281 64705 37315
rect 64739 37281 64751 37315
rect 64693 37275 64751 37281
rect 64785 37315 64843 37321
rect 64785 37281 64797 37315
rect 64831 37281 64843 37315
rect 64785 37275 64843 37281
rect 65061 37315 65119 37321
rect 65061 37281 65073 37315
rect 65107 37312 65119 37315
rect 65334 37312 65340 37324
rect 65107 37284 65340 37312
rect 65107 37281 65119 37284
rect 65061 37275 65119 37281
rect 42150 37244 42156 37256
rect 40052 37216 42156 37244
rect 42150 37204 42156 37216
rect 42208 37204 42214 37256
rect 44910 37244 44916 37256
rect 44871 37216 44916 37244
rect 44910 37204 44916 37216
rect 44968 37204 44974 37256
rect 45186 37244 45192 37256
rect 45147 37216 45192 37244
rect 45186 37204 45192 37216
rect 45244 37204 45250 37256
rect 53098 37204 53104 37256
rect 53156 37204 53162 37256
rect 64141 37247 64199 37253
rect 64141 37213 64153 37247
rect 64187 37213 64199 37247
rect 64708 37244 64736 37275
rect 65334 37272 65340 37284
rect 65392 37312 65398 37324
rect 65812 37321 65840 37352
rect 66990 37340 66996 37352
rect 67048 37340 67054 37392
rect 78766 37380 78772 37392
rect 67100 37352 78772 37380
rect 65797 37315 65855 37321
rect 65392 37284 65748 37312
rect 65392 37272 65398 37284
rect 65242 37244 65248 37256
rect 64708 37216 65248 37244
rect 64141 37207 64199 37213
rect 34517 37179 34575 37185
rect 34517 37176 34529 37179
rect 33008 37148 34529 37176
rect 33008 37136 33014 37148
rect 34517 37145 34529 37148
rect 34563 37145 34575 37179
rect 34517 37139 34575 37145
rect 32214 37108 32220 37120
rect 31987 37080 32220 37108
rect 31987 37077 31999 37080
rect 31941 37071 31999 37077
rect 32214 37068 32220 37080
rect 32272 37068 32278 37120
rect 32766 37068 32772 37120
rect 32824 37108 32830 37120
rect 34149 37111 34207 37117
rect 34149 37108 34161 37111
rect 32824 37080 34161 37108
rect 32824 37068 32830 37080
rect 34149 37077 34161 37080
rect 34195 37108 34207 37111
rect 34330 37108 34336 37120
rect 34195 37080 34336 37108
rect 34195 37077 34207 37080
rect 34149 37071 34207 37077
rect 34330 37068 34336 37080
rect 34388 37068 34394 37120
rect 38378 37068 38384 37120
rect 38436 37108 38442 37120
rect 38930 37108 38936 37120
rect 38436 37080 38936 37108
rect 38436 37068 38442 37080
rect 38930 37068 38936 37080
rect 38988 37108 38994 37120
rect 41049 37111 41107 37117
rect 41049 37108 41061 37111
rect 38988 37080 41061 37108
rect 38988 37068 38994 37080
rect 41049 37077 41061 37080
rect 41095 37077 41107 37111
rect 41049 37071 41107 37077
rect 44637 37111 44695 37117
rect 44637 37077 44649 37111
rect 44683 37108 44695 37111
rect 44726 37108 44732 37120
rect 44683 37080 44732 37108
rect 44683 37077 44695 37080
rect 44637 37071 44695 37077
rect 44726 37068 44732 37080
rect 44784 37068 44790 37120
rect 46750 37108 46756 37120
rect 46711 37080 46756 37108
rect 46750 37068 46756 37080
rect 46808 37068 46814 37120
rect 63218 37068 63224 37120
rect 63276 37108 63282 37120
rect 63497 37111 63555 37117
rect 63497 37108 63509 37111
rect 63276 37080 63509 37108
rect 63276 37068 63282 37080
rect 63497 37077 63509 37080
rect 63543 37108 63555 37111
rect 64156 37108 64184 37207
rect 65242 37204 65248 37216
rect 65300 37204 65306 37256
rect 65720 37244 65748 37284
rect 65797 37281 65809 37315
rect 65843 37281 65855 37315
rect 65797 37275 65855 37281
rect 65978 37272 65984 37324
rect 66036 37312 66042 37324
rect 66073 37315 66131 37321
rect 66073 37312 66085 37315
rect 66036 37284 66085 37312
rect 66036 37272 66042 37284
rect 66073 37281 66085 37284
rect 66119 37281 66131 37315
rect 67100 37312 67128 37352
rect 78766 37340 78772 37352
rect 78824 37380 78830 37392
rect 79137 37383 79195 37389
rect 79137 37380 79149 37383
rect 78824 37352 79149 37380
rect 78824 37340 78830 37352
rect 79137 37349 79149 37352
rect 79183 37349 79195 37383
rect 79318 37380 79324 37392
rect 79279 37352 79324 37380
rect 79137 37343 79195 37349
rect 70118 37312 70124 37324
rect 66073 37275 66131 37281
rect 66180 37284 67128 37312
rect 70079 37284 70124 37312
rect 66180 37244 66208 37284
rect 70118 37272 70124 37284
rect 70176 37272 70182 37324
rect 70213 37315 70271 37321
rect 70213 37281 70225 37315
rect 70259 37312 70271 37315
rect 71130 37312 71136 37324
rect 70259 37284 71136 37312
rect 70259 37281 70271 37284
rect 70213 37275 70271 37281
rect 71130 37272 71136 37284
rect 71188 37272 71194 37324
rect 72237 37315 72295 37321
rect 72237 37281 72249 37315
rect 72283 37312 72295 37315
rect 72510 37312 72516 37324
rect 72283 37284 72516 37312
rect 72283 37281 72295 37284
rect 72237 37275 72295 37281
rect 72510 37272 72516 37284
rect 72568 37312 72574 37324
rect 72568 37284 73108 37312
rect 72568 37272 72574 37284
rect 65720 37216 66208 37244
rect 73080 37244 73108 37284
rect 73154 37272 73160 37324
rect 73212 37312 73218 37324
rect 73341 37315 73399 37321
rect 73341 37312 73353 37315
rect 73212 37284 73353 37312
rect 73212 37272 73218 37284
rect 73341 37281 73353 37284
rect 73387 37281 73399 37315
rect 77202 37312 77208 37324
rect 73341 37275 73399 37281
rect 73448 37284 77208 37312
rect 73448 37244 73476 37284
rect 77202 37272 77208 37284
rect 77260 37272 77266 37324
rect 73080 37216 73476 37244
rect 79152 37244 79180 37343
rect 79318 37340 79324 37352
rect 79376 37380 79382 37392
rect 80164 37389 80192 37420
rect 80149 37383 80207 37389
rect 80149 37380 80161 37383
rect 79376 37352 80161 37380
rect 79376 37340 79382 37352
rect 80149 37349 80161 37352
rect 80195 37349 80207 37383
rect 80882 37380 80888 37392
rect 80843 37352 80888 37380
rect 80149 37343 80207 37349
rect 80882 37340 80888 37352
rect 80940 37340 80946 37392
rect 79468 37315 79526 37321
rect 79468 37281 79480 37315
rect 79514 37312 79526 37315
rect 79870 37312 79876 37324
rect 79514 37284 79876 37312
rect 79514 37281 79526 37284
rect 79468 37275 79526 37281
rect 79870 37272 79876 37284
rect 79928 37272 79934 37324
rect 81069 37315 81127 37321
rect 81069 37281 81081 37315
rect 81115 37312 81127 37315
rect 81342 37312 81348 37324
rect 81115 37284 81348 37312
rect 81115 37281 81127 37284
rect 81069 37275 81127 37281
rect 79686 37244 79692 37256
rect 79152 37216 79692 37244
rect 79686 37204 79692 37216
rect 79744 37204 79750 37256
rect 79778 37204 79784 37256
rect 79836 37244 79842 37256
rect 81084 37244 81112 37275
rect 81342 37272 81348 37284
rect 81400 37312 81406 37324
rect 81529 37315 81587 37321
rect 81529 37312 81541 37315
rect 81400 37284 81541 37312
rect 81400 37272 81406 37284
rect 81529 37281 81541 37284
rect 81575 37281 81587 37315
rect 84120 37312 84148 37420
rect 84194 37408 84200 37460
rect 84252 37448 84258 37460
rect 86129 37451 86187 37457
rect 86129 37448 86141 37451
rect 84252 37420 86141 37448
rect 84252 37408 84258 37420
rect 86129 37417 86141 37420
rect 86175 37417 86187 37451
rect 86129 37411 86187 37417
rect 85574 37380 85580 37392
rect 85535 37352 85580 37380
rect 85574 37340 85580 37352
rect 85632 37380 85638 37392
rect 85632 37352 85988 37380
rect 85632 37340 85638 37352
rect 85960 37324 85988 37352
rect 86512 37352 88472 37380
rect 85669 37315 85727 37321
rect 84120 37284 85620 37312
rect 81529 37275 81587 37281
rect 79836 37216 81112 37244
rect 85592 37244 85620 37284
rect 85669 37281 85681 37315
rect 85715 37312 85727 37315
rect 85850 37312 85856 37324
rect 85715 37284 85856 37312
rect 85715 37281 85727 37284
rect 85669 37275 85727 37281
rect 85850 37272 85856 37284
rect 85908 37272 85914 37324
rect 85942 37272 85948 37324
rect 86000 37312 86006 37324
rect 86000 37284 86093 37312
rect 86000 37272 86006 37284
rect 85758 37244 85764 37256
rect 85592 37216 85764 37244
rect 79836 37204 79842 37216
rect 85758 37204 85764 37216
rect 85816 37244 85822 37256
rect 86512 37253 86540 37352
rect 87322 37272 87328 37324
rect 87380 37312 87386 37324
rect 88444 37321 88472 37352
rect 88245 37315 88303 37321
rect 88245 37312 88257 37315
rect 87380 37284 88257 37312
rect 87380 37272 87386 37284
rect 88245 37281 88257 37284
rect 88291 37281 88303 37315
rect 88245 37275 88303 37281
rect 88429 37315 88487 37321
rect 88429 37281 88441 37315
rect 88475 37312 88487 37315
rect 88889 37315 88947 37321
rect 88889 37312 88901 37315
rect 88475 37284 88901 37312
rect 88475 37281 88487 37284
rect 88429 37275 88487 37281
rect 88889 37281 88901 37284
rect 88935 37281 88947 37315
rect 88889 37275 88947 37281
rect 86497 37247 86555 37253
rect 86497 37244 86509 37247
rect 85816 37216 86509 37244
rect 85816 37204 85822 37216
rect 86497 37213 86509 37216
rect 86543 37213 86555 37247
rect 86497 37207 86555 37213
rect 64874 37136 64880 37188
rect 64932 37176 64938 37188
rect 65889 37179 65947 37185
rect 65889 37176 65901 37179
rect 64932 37148 65901 37176
rect 64932 37136 64938 37148
rect 65889 37145 65901 37148
rect 65935 37145 65947 37179
rect 65889 37139 65947 37145
rect 78950 37136 78956 37188
rect 79008 37176 79014 37188
rect 79597 37179 79655 37185
rect 79597 37176 79609 37179
rect 79008 37148 79609 37176
rect 79008 37136 79014 37148
rect 79597 37145 79609 37148
rect 79643 37145 79655 37179
rect 79597 37139 79655 37145
rect 65242 37108 65248 37120
rect 63543 37080 64184 37108
rect 65203 37080 65248 37108
rect 63543 37077 63555 37080
rect 63497 37071 63555 37077
rect 65242 37068 65248 37080
rect 65300 37068 65306 37120
rect 79962 37108 79968 37120
rect 79923 37080 79968 37108
rect 79962 37068 79968 37080
rect 80020 37068 80026 37120
rect 80422 37068 80428 37120
rect 80480 37108 80486 37120
rect 81161 37111 81219 37117
rect 81161 37108 81173 37111
rect 80480 37080 81173 37108
rect 80480 37068 80486 37080
rect 81161 37077 81173 37080
rect 81207 37077 81219 37111
rect 81161 37071 81219 37077
rect 88426 37068 88432 37120
rect 88484 37108 88490 37120
rect 88521 37111 88579 37117
rect 88521 37108 88533 37111
rect 88484 37080 88533 37108
rect 88484 37068 88490 37080
rect 88521 37077 88533 37080
rect 88567 37077 88579 37111
rect 88521 37071 88579 37077
rect 1104 37018 108008 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 65686 37018
rect 65738 36966 65750 37018
rect 65802 36966 65814 37018
rect 65866 36966 65878 37018
rect 65930 36966 96406 37018
rect 96458 36966 96470 37018
rect 96522 36966 96534 37018
rect 96586 36966 96598 37018
rect 96650 36966 108008 37018
rect 1104 36944 108008 36966
rect 5445 36907 5503 36913
rect 5445 36873 5457 36907
rect 5491 36904 5503 36907
rect 5718 36904 5724 36916
rect 5491 36876 5724 36904
rect 5491 36873 5503 36876
rect 5445 36867 5503 36873
rect 4798 36796 4804 36848
rect 4856 36836 4862 36848
rect 4985 36839 5043 36845
rect 4985 36836 4997 36839
rect 4856 36808 4997 36836
rect 4856 36796 4862 36808
rect 4985 36805 4997 36808
rect 5031 36805 5043 36839
rect 4985 36799 5043 36805
rect 3786 36700 3792 36712
rect 3699 36672 3792 36700
rect 3326 36524 3332 36576
rect 3384 36564 3390 36576
rect 3712 36573 3740 36672
rect 3786 36660 3792 36672
rect 3844 36700 3850 36712
rect 3881 36703 3939 36709
rect 3881 36700 3893 36703
rect 3844 36672 3893 36700
rect 3844 36660 3850 36672
rect 3881 36669 3893 36672
rect 3927 36669 3939 36703
rect 3881 36663 3939 36669
rect 4065 36703 4123 36709
rect 4065 36669 4077 36703
rect 4111 36700 4123 36703
rect 4617 36703 4675 36709
rect 4617 36700 4629 36703
rect 4111 36672 4629 36700
rect 4111 36669 4123 36672
rect 4065 36663 4123 36669
rect 4617 36669 4629 36672
rect 4663 36669 4675 36703
rect 4617 36663 4675 36669
rect 4801 36703 4859 36709
rect 4801 36669 4813 36703
rect 4847 36700 4859 36703
rect 5460 36700 5488 36867
rect 5718 36864 5724 36876
rect 5776 36864 5782 36916
rect 9769 36907 9827 36913
rect 9769 36873 9781 36907
rect 9815 36904 9827 36907
rect 9858 36904 9864 36916
rect 9815 36876 9864 36904
rect 9815 36873 9827 36876
rect 9769 36867 9827 36873
rect 9858 36864 9864 36876
rect 9916 36864 9922 36916
rect 9950 36864 9956 36916
rect 10008 36904 10014 36916
rect 11054 36904 11060 36916
rect 10008 36876 11060 36904
rect 10008 36864 10014 36876
rect 11054 36864 11060 36876
rect 11112 36864 11118 36916
rect 19242 36864 19248 36916
rect 19300 36904 19306 36916
rect 33137 36907 33195 36913
rect 19300 36876 33088 36904
rect 19300 36864 19306 36876
rect 5534 36796 5540 36848
rect 5592 36836 5598 36848
rect 16390 36836 16396 36848
rect 5592 36808 16396 36836
rect 5592 36796 5598 36808
rect 16390 36796 16396 36808
rect 16448 36796 16454 36848
rect 16666 36836 16672 36848
rect 16627 36808 16672 36836
rect 16666 36796 16672 36808
rect 16724 36796 16730 36848
rect 22281 36839 22339 36845
rect 22281 36836 22293 36839
rect 21560 36808 22293 36836
rect 8297 36771 8355 36777
rect 8297 36737 8309 36771
rect 8343 36768 8355 36771
rect 9122 36768 9128 36780
rect 8343 36740 9128 36768
rect 8343 36737 8355 36740
rect 8297 36731 8355 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 9950 36768 9956 36780
rect 9416 36740 9956 36768
rect 9416 36709 9444 36740
rect 9950 36728 9956 36740
rect 10008 36728 10014 36780
rect 16574 36728 16580 36780
rect 16632 36768 16638 36780
rect 21560 36777 21588 36808
rect 22281 36805 22293 36808
rect 22327 36836 22339 36839
rect 25498 36836 25504 36848
rect 22327 36808 25504 36836
rect 22327 36805 22339 36808
rect 22281 36799 22339 36805
rect 25498 36796 25504 36808
rect 25556 36796 25562 36848
rect 26234 36836 26240 36848
rect 25608 36808 26240 36836
rect 20809 36771 20867 36777
rect 20809 36768 20821 36771
rect 16632 36740 20821 36768
rect 16632 36728 16638 36740
rect 20809 36737 20821 36740
rect 20855 36737 20867 36771
rect 20809 36731 20867 36737
rect 21545 36771 21603 36777
rect 21545 36737 21557 36771
rect 21591 36737 21603 36771
rect 21545 36731 21603 36737
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36768 22247 36771
rect 25608 36768 25636 36808
rect 26234 36796 26240 36808
rect 26292 36796 26298 36848
rect 26326 36796 26332 36848
rect 26384 36836 26390 36848
rect 33060 36836 33088 36876
rect 33137 36873 33149 36907
rect 33183 36904 33195 36907
rect 33318 36904 33324 36916
rect 33183 36876 33324 36904
rect 33183 36873 33195 36876
rect 33137 36867 33195 36873
rect 33318 36864 33324 36876
rect 33376 36864 33382 36916
rect 38657 36907 38715 36913
rect 38657 36873 38669 36907
rect 38703 36904 38715 36907
rect 38746 36904 38752 36916
rect 38703 36876 38752 36904
rect 38703 36873 38715 36876
rect 38657 36867 38715 36873
rect 38746 36864 38752 36876
rect 38804 36864 38810 36916
rect 43533 36907 43591 36913
rect 42996 36876 43208 36904
rect 42996 36836 43024 36876
rect 26384 36808 26429 36836
rect 33060 36808 43024 36836
rect 43180 36836 43208 36876
rect 43533 36873 43545 36907
rect 43579 36904 43591 36907
rect 47854 36904 47860 36916
rect 43579 36876 47860 36904
rect 43579 36873 43591 36876
rect 43533 36867 43591 36873
rect 43548 36836 43576 36867
rect 47854 36864 47860 36876
rect 47912 36864 47918 36916
rect 50706 36904 50712 36916
rect 50667 36876 50712 36904
rect 50706 36864 50712 36876
rect 50764 36864 50770 36916
rect 50816 36876 52776 36904
rect 43180 36808 43576 36836
rect 26384 36796 26390 36808
rect 26421 36771 26479 36777
rect 26421 36768 26433 36771
rect 22235 36740 25636 36768
rect 25700 36740 26433 36768
rect 22235 36737 22247 36740
rect 22189 36731 22247 36737
rect 4847 36672 5488 36700
rect 9033 36703 9091 36709
rect 4847 36669 4859 36672
rect 4801 36663 4859 36669
rect 9033 36669 9045 36703
rect 9079 36669 9091 36703
rect 9033 36663 9091 36669
rect 9401 36703 9459 36709
rect 9401 36669 9413 36703
rect 9447 36669 9459 36703
rect 9401 36663 9459 36669
rect 9585 36703 9643 36709
rect 9585 36669 9597 36703
rect 9631 36700 9643 36703
rect 9858 36700 9864 36712
rect 9631 36672 9864 36700
rect 9631 36669 9643 36672
rect 9585 36663 9643 36669
rect 4632 36632 4660 36663
rect 4632 36604 5120 36632
rect 5092 36576 5120 36604
rect 6914 36592 6920 36644
rect 6972 36632 6978 36644
rect 8389 36635 8447 36641
rect 8389 36632 8401 36635
rect 6972 36604 8401 36632
rect 6972 36592 6978 36604
rect 8389 36601 8401 36604
rect 8435 36601 8447 36635
rect 9048 36632 9076 36663
rect 9858 36660 9864 36672
rect 9916 36660 9922 36712
rect 13538 36700 13544 36712
rect 13499 36672 13544 36700
rect 13538 36660 13544 36672
rect 13596 36660 13602 36712
rect 14274 36700 14280 36712
rect 14235 36672 14280 36700
rect 14274 36660 14280 36672
rect 14332 36660 14338 36712
rect 14553 36703 14611 36709
rect 14553 36669 14565 36703
rect 14599 36700 14611 36703
rect 15286 36700 15292 36712
rect 14599 36672 15292 36700
rect 14599 36669 14611 36672
rect 14553 36663 14611 36669
rect 15286 36660 15292 36672
rect 15344 36660 15350 36712
rect 15933 36703 15991 36709
rect 15933 36669 15945 36703
rect 15979 36700 15991 36703
rect 16485 36703 16543 36709
rect 16485 36700 16497 36703
rect 15979 36672 16497 36700
rect 15979 36669 15991 36672
rect 15933 36663 15991 36669
rect 16485 36669 16497 36672
rect 16531 36700 16543 36703
rect 19242 36700 19248 36712
rect 16531 36672 19248 36700
rect 16531 36669 16543 36672
rect 16485 36663 16543 36669
rect 19242 36660 19248 36672
rect 19300 36660 19306 36712
rect 21450 36700 21456 36712
rect 21411 36672 21456 36700
rect 21450 36660 21456 36672
rect 21508 36660 21514 36712
rect 21818 36700 21824 36712
rect 21779 36672 21824 36700
rect 21818 36660 21824 36672
rect 21876 36660 21882 36712
rect 22005 36703 22063 36709
rect 22005 36669 22017 36703
rect 22051 36700 22063 36703
rect 22204 36700 22232 36731
rect 22051 36672 22232 36700
rect 22051 36669 22063 36672
rect 22005 36663 22063 36669
rect 9766 36632 9772 36644
rect 9048 36604 9772 36632
rect 8389 36595 8447 36601
rect 9766 36592 9772 36604
rect 9824 36592 9830 36644
rect 15749 36635 15807 36641
rect 15749 36601 15761 36635
rect 15795 36632 15807 36635
rect 16666 36632 16672 36644
rect 15795 36604 16672 36632
rect 15795 36601 15807 36604
rect 15749 36595 15807 36601
rect 16666 36592 16672 36604
rect 16724 36592 16730 36644
rect 21836 36632 21864 36660
rect 22465 36635 22523 36641
rect 22465 36632 22477 36635
rect 21836 36604 22477 36632
rect 22465 36601 22477 36604
rect 22511 36601 22523 36635
rect 22465 36595 22523 36601
rect 3697 36567 3755 36573
rect 3697 36564 3709 36567
rect 3384 36536 3709 36564
rect 3384 36524 3390 36536
rect 3697 36533 3709 36536
rect 3743 36533 3755 36567
rect 3697 36527 3755 36533
rect 5074 36524 5080 36576
rect 5132 36564 5138 36576
rect 5537 36567 5595 36573
rect 5537 36564 5549 36567
rect 5132 36536 5549 36564
rect 5132 36524 5138 36536
rect 5537 36533 5549 36536
rect 5583 36564 5595 36567
rect 5721 36567 5779 36573
rect 5721 36564 5733 36567
rect 5583 36536 5733 36564
rect 5583 36533 5595 36536
rect 5537 36527 5595 36533
rect 5721 36533 5733 36536
rect 5767 36533 5779 36567
rect 13630 36564 13636 36576
rect 13591 36536 13636 36564
rect 5721 36527 5779 36533
rect 13630 36524 13636 36536
rect 13688 36524 13694 36576
rect 16022 36564 16028 36576
rect 15983 36536 16028 36564
rect 16022 36524 16028 36536
rect 16080 36524 16086 36576
rect 24762 36524 24768 36576
rect 24820 36564 24826 36576
rect 25700 36573 25728 36740
rect 26421 36737 26433 36740
rect 26467 36737 26479 36771
rect 26421 36731 26479 36737
rect 37185 36771 37243 36777
rect 37185 36737 37197 36771
rect 37231 36768 37243 36771
rect 37231 36740 37688 36768
rect 37231 36737 37243 36740
rect 37185 36731 37243 36737
rect 37660 36712 37688 36740
rect 26200 36703 26258 36709
rect 26200 36669 26212 36703
rect 26246 36700 26258 36703
rect 26602 36700 26608 36712
rect 26246 36672 26608 36700
rect 26246 36669 26258 36672
rect 26200 36663 26258 36669
rect 26602 36660 26608 36672
rect 26660 36660 26666 36712
rect 31941 36703 31999 36709
rect 31941 36669 31953 36703
rect 31987 36669 31999 36703
rect 31941 36663 31999 36669
rect 32125 36703 32183 36709
rect 32125 36669 32137 36703
rect 32171 36700 32183 36703
rect 32674 36700 32680 36712
rect 32171 36672 32680 36700
rect 32171 36669 32183 36672
rect 32125 36663 32183 36669
rect 26050 36632 26056 36644
rect 26011 36604 26056 36632
rect 26050 36592 26056 36604
rect 26108 36592 26114 36644
rect 26326 36592 26332 36644
rect 26384 36632 26390 36644
rect 30374 36632 30380 36644
rect 26384 36604 30380 36632
rect 26384 36592 26390 36604
rect 30374 36592 30380 36604
rect 30432 36592 30438 36644
rect 31849 36635 31907 36641
rect 31849 36601 31861 36635
rect 31895 36632 31907 36635
rect 31956 36632 31984 36663
rect 32674 36660 32680 36672
rect 32732 36660 32738 36712
rect 32861 36703 32919 36709
rect 32861 36669 32873 36703
rect 32907 36700 32919 36703
rect 33226 36700 33232 36712
rect 32907 36672 33232 36700
rect 32907 36669 32919 36672
rect 32861 36663 32919 36669
rect 33226 36660 33232 36672
rect 33284 36700 33290 36712
rect 33686 36700 33692 36712
rect 33284 36672 33692 36700
rect 33284 36660 33290 36672
rect 33686 36660 33692 36672
rect 33744 36660 33750 36712
rect 37461 36703 37519 36709
rect 37461 36700 37473 36703
rect 37384 36672 37473 36700
rect 32214 36632 32220 36644
rect 31895 36604 32220 36632
rect 31895 36601 31907 36604
rect 31849 36595 31907 36601
rect 32214 36592 32220 36604
rect 32272 36592 32278 36644
rect 32582 36592 32588 36644
rect 32640 36632 32646 36644
rect 37090 36632 37096 36644
rect 32640 36604 37096 36632
rect 32640 36592 32646 36604
rect 37090 36592 37096 36604
rect 37148 36592 37154 36644
rect 37384 36576 37412 36672
rect 37461 36669 37473 36672
rect 37507 36669 37519 36703
rect 37642 36700 37648 36712
rect 37603 36672 37648 36700
rect 37461 36663 37519 36669
rect 37642 36660 37648 36672
rect 37700 36660 37706 36712
rect 38102 36660 38108 36712
rect 38160 36700 38166 36712
rect 38243 36703 38301 36709
rect 38243 36700 38255 36703
rect 38160 36672 38255 36700
rect 38160 36660 38166 36672
rect 38243 36669 38255 36672
rect 38289 36669 38301 36703
rect 38243 36663 38301 36669
rect 38378 36660 38384 36712
rect 38436 36700 38442 36712
rect 41785 36703 41843 36709
rect 41785 36700 41797 36703
rect 38436 36672 38481 36700
rect 38580 36672 41797 36700
rect 38436 36660 38442 36672
rect 37734 36592 37740 36644
rect 37792 36632 37798 36644
rect 38580 36632 38608 36672
rect 41785 36669 41797 36672
rect 41831 36700 41843 36703
rect 41969 36703 42027 36709
rect 41969 36700 41981 36703
rect 41831 36672 41981 36700
rect 41831 36669 41843 36672
rect 41785 36663 41843 36669
rect 41969 36669 41981 36672
rect 42015 36669 42027 36703
rect 42150 36700 42156 36712
rect 42111 36672 42156 36700
rect 41969 36663 42027 36669
rect 42150 36660 42156 36672
rect 42208 36700 42214 36712
rect 42705 36703 42763 36709
rect 42705 36700 42717 36703
rect 42208 36672 42717 36700
rect 42208 36660 42214 36672
rect 42705 36669 42717 36672
rect 42751 36669 42763 36703
rect 42705 36663 42763 36669
rect 42889 36703 42947 36709
rect 42889 36669 42901 36703
rect 42935 36700 42947 36703
rect 43180 36700 43208 36808
rect 48130 36796 48136 36848
rect 48188 36836 48194 36848
rect 48225 36839 48283 36845
rect 48225 36836 48237 36839
rect 48188 36808 48237 36836
rect 48188 36796 48194 36808
rect 48225 36805 48237 36808
rect 48271 36836 48283 36839
rect 50816 36836 50844 36876
rect 48271 36808 50844 36836
rect 48271 36805 48283 36808
rect 48225 36799 48283 36805
rect 51350 36796 51356 36848
rect 51408 36836 51414 36848
rect 51445 36839 51503 36845
rect 51445 36836 51457 36839
rect 51408 36808 51457 36836
rect 51408 36796 51414 36808
rect 51445 36805 51457 36808
rect 51491 36836 51503 36839
rect 51718 36836 51724 36848
rect 51491 36808 51724 36836
rect 51491 36805 51503 36808
rect 51445 36799 51503 36805
rect 51718 36796 51724 36808
rect 51776 36796 51782 36848
rect 43257 36771 43315 36777
rect 43257 36737 43269 36771
rect 43303 36768 43315 36771
rect 46937 36771 46995 36777
rect 46937 36768 46949 36771
rect 43303 36740 46949 36768
rect 43303 36737 43315 36740
rect 43257 36731 43315 36737
rect 46937 36737 46949 36740
rect 46983 36737 46995 36771
rect 46937 36731 46995 36737
rect 50798 36728 50804 36780
rect 50856 36768 50862 36780
rect 51997 36771 52055 36777
rect 51997 36768 52009 36771
rect 50856 36740 52009 36768
rect 50856 36728 50862 36740
rect 51997 36737 52009 36740
rect 52043 36737 52055 36771
rect 52748 36768 52776 36876
rect 59906 36864 59912 36916
rect 59964 36904 59970 36916
rect 60918 36904 60924 36916
rect 59964 36876 60924 36904
rect 59964 36864 59970 36876
rect 60918 36864 60924 36876
rect 60976 36864 60982 36916
rect 64233 36907 64291 36913
rect 64233 36873 64245 36907
rect 64279 36904 64291 36907
rect 64874 36904 64880 36916
rect 64279 36876 64880 36904
rect 64279 36873 64291 36876
rect 64233 36867 64291 36873
rect 64874 36864 64880 36876
rect 64932 36864 64938 36916
rect 65242 36864 65248 36916
rect 65300 36904 65306 36916
rect 65521 36907 65579 36913
rect 65521 36904 65533 36907
rect 65300 36876 65533 36904
rect 65300 36864 65306 36876
rect 65521 36873 65533 36876
rect 65567 36904 65579 36907
rect 65567 36876 78720 36904
rect 65567 36873 65579 36876
rect 65521 36867 65579 36873
rect 65334 36836 65340 36848
rect 65295 36808 65340 36836
rect 65334 36796 65340 36808
rect 65392 36796 65398 36848
rect 66070 36836 66076 36848
rect 66031 36808 66076 36836
rect 66070 36796 66076 36808
rect 66128 36796 66134 36848
rect 78692 36836 78720 36876
rect 78766 36864 78772 36916
rect 78824 36904 78830 36916
rect 78824 36876 78869 36904
rect 78824 36864 78830 36876
rect 79134 36864 79140 36916
rect 79192 36904 79198 36916
rect 79870 36904 79876 36916
rect 79192 36876 79876 36904
rect 79192 36864 79198 36876
rect 79870 36864 79876 36876
rect 79928 36904 79934 36916
rect 80057 36907 80115 36913
rect 80057 36904 80069 36907
rect 79928 36876 80069 36904
rect 79928 36864 79934 36876
rect 80057 36873 80069 36876
rect 80103 36873 80115 36907
rect 80057 36867 80115 36873
rect 83902 36907 83960 36913
rect 83902 36873 83914 36907
rect 83948 36904 83960 36907
rect 84746 36904 84752 36916
rect 83948 36876 84752 36904
rect 83948 36873 83960 36876
rect 83902 36867 83960 36873
rect 84746 36864 84752 36876
rect 84804 36864 84810 36916
rect 85390 36864 85396 36916
rect 85448 36904 85454 36916
rect 85761 36907 85819 36913
rect 85761 36904 85773 36907
rect 85448 36876 85773 36904
rect 85448 36864 85454 36876
rect 85761 36873 85773 36876
rect 85807 36873 85819 36907
rect 85942 36904 85948 36916
rect 85903 36876 85948 36904
rect 85761 36867 85819 36873
rect 78953 36839 79011 36845
rect 78953 36836 78965 36839
rect 78692 36808 78965 36836
rect 52748 36740 61976 36768
rect 51997 36731 52055 36737
rect 42935 36672 43208 36700
rect 46661 36703 46719 36709
rect 42935 36669 42947 36672
rect 42889 36663 42947 36669
rect 46661 36669 46673 36703
rect 46707 36700 46719 36703
rect 46750 36700 46756 36712
rect 46707 36672 46756 36700
rect 46707 36669 46719 36672
rect 46661 36663 46719 36669
rect 37792 36604 38608 36632
rect 42720 36632 42748 36663
rect 46750 36660 46756 36672
rect 46808 36700 46814 36712
rect 50617 36703 50675 36709
rect 46808 36672 48544 36700
rect 46808 36660 46814 36672
rect 43714 36632 43720 36644
rect 42720 36604 43720 36632
rect 37792 36592 37798 36604
rect 43714 36592 43720 36604
rect 43772 36592 43778 36644
rect 48516 36576 48544 36672
rect 50617 36669 50629 36703
rect 50663 36669 50675 36703
rect 51718 36700 51724 36712
rect 51679 36672 51724 36700
rect 50617 36663 50675 36669
rect 50632 36632 50660 36663
rect 51718 36660 51724 36672
rect 51776 36660 51782 36712
rect 58161 36703 58219 36709
rect 58161 36669 58173 36703
rect 58207 36669 58219 36703
rect 58434 36700 58440 36712
rect 58395 36672 58440 36700
rect 58161 36663 58219 36669
rect 50632 36604 51120 36632
rect 25685 36567 25743 36573
rect 25685 36564 25697 36567
rect 24820 36536 25697 36564
rect 24820 36524 24826 36536
rect 25685 36533 25697 36536
rect 25731 36533 25743 36567
rect 25866 36564 25872 36576
rect 25827 36536 25872 36564
rect 25685 36527 25743 36533
rect 25866 36524 25872 36536
rect 25924 36524 25930 36576
rect 26697 36567 26755 36573
rect 26697 36533 26709 36567
rect 26743 36564 26755 36567
rect 36630 36564 36636 36576
rect 26743 36536 36636 36564
rect 26743 36533 26755 36536
rect 26697 36527 26755 36533
rect 36630 36524 36636 36536
rect 36688 36524 36694 36576
rect 37366 36564 37372 36576
rect 37327 36536 37372 36564
rect 37366 36524 37372 36536
rect 37424 36524 37430 36576
rect 48498 36564 48504 36576
rect 48459 36536 48504 36564
rect 48498 36524 48504 36536
rect 48556 36524 48562 36576
rect 51092 36564 51120 36604
rect 52362 36564 52368 36576
rect 51092 36536 52368 36564
rect 52362 36524 52368 36536
rect 52420 36524 52426 36576
rect 53098 36564 53104 36576
rect 53059 36536 53104 36564
rect 53098 36524 53104 36536
rect 53156 36524 53162 36576
rect 58176 36564 58204 36663
rect 58434 36660 58440 36672
rect 58492 36660 58498 36712
rect 61948 36700 61976 36740
rect 62022 36728 62028 36780
rect 62080 36768 62086 36780
rect 64877 36771 64935 36777
rect 64877 36768 64889 36771
rect 62080 36740 64889 36768
rect 62080 36728 62086 36740
rect 64877 36737 64889 36740
rect 64923 36737 64935 36771
rect 64877 36731 64935 36737
rect 64414 36700 64420 36712
rect 61948 36672 63264 36700
rect 64375 36672 64420 36700
rect 59817 36635 59875 36641
rect 59817 36601 59829 36635
rect 59863 36632 59875 36635
rect 63126 36632 63132 36644
rect 59863 36604 63132 36632
rect 59863 36601 59875 36604
rect 59817 36595 59875 36601
rect 63126 36592 63132 36604
rect 63184 36592 63190 36644
rect 59906 36564 59912 36576
rect 58176 36536 59912 36564
rect 59906 36524 59912 36536
rect 59964 36524 59970 36576
rect 63236 36564 63264 36672
rect 64414 36660 64420 36672
rect 64472 36660 64478 36712
rect 64598 36700 64604 36712
rect 64511 36672 64604 36700
rect 64598 36660 64604 36672
rect 64656 36660 64662 36712
rect 64969 36703 65027 36709
rect 64969 36669 64981 36703
rect 65015 36700 65027 36703
rect 65242 36700 65248 36712
rect 65015 36672 65248 36700
rect 65015 36669 65027 36672
rect 64969 36663 65027 36669
rect 65242 36660 65248 36672
rect 65300 36660 65306 36712
rect 64616 36632 64644 36660
rect 65352 36632 65380 36796
rect 66438 36768 66444 36780
rect 66399 36740 66444 36768
rect 66438 36728 66444 36740
rect 66496 36728 66502 36780
rect 71130 36768 71136 36780
rect 71091 36740 71136 36768
rect 71130 36728 71136 36740
rect 71188 36728 71194 36780
rect 65978 36700 65984 36712
rect 65939 36672 65984 36700
rect 65978 36660 65984 36672
rect 66036 36660 66042 36712
rect 66162 36660 66168 36712
rect 66220 36700 66226 36712
rect 66257 36703 66315 36709
rect 66257 36700 66269 36703
rect 66220 36672 66269 36700
rect 66220 36660 66226 36672
rect 66257 36669 66269 36672
rect 66303 36669 66315 36703
rect 66257 36663 66315 36669
rect 70857 36703 70915 36709
rect 70857 36669 70869 36703
rect 70903 36700 70915 36703
rect 75914 36700 75920 36712
rect 70903 36672 72740 36700
rect 75875 36672 75920 36700
rect 70903 36669 70915 36672
rect 70857 36663 70915 36669
rect 64616 36604 65380 36632
rect 65426 36592 65432 36644
rect 65484 36632 65490 36644
rect 68646 36632 68652 36644
rect 65484 36604 68652 36632
rect 65484 36592 65490 36604
rect 68646 36592 68652 36604
rect 68704 36592 68710 36644
rect 68094 36564 68100 36576
rect 63236 36536 68100 36564
rect 68094 36524 68100 36536
rect 68152 36524 68158 36576
rect 72418 36564 72424 36576
rect 72379 36536 72424 36564
rect 72418 36524 72424 36536
rect 72476 36524 72482 36576
rect 72712 36573 72740 36672
rect 75914 36660 75920 36672
rect 75972 36660 75978 36712
rect 78692 36709 78720 36808
rect 78953 36805 78965 36808
rect 78999 36836 79011 36839
rect 79778 36836 79784 36848
rect 78999 36808 79784 36836
rect 78999 36805 79011 36808
rect 78953 36799 79011 36805
rect 79778 36796 79784 36808
rect 79836 36796 79842 36848
rect 79962 36796 79968 36848
rect 80020 36836 80026 36848
rect 81529 36839 81587 36845
rect 81529 36836 81541 36839
rect 80020 36808 81541 36836
rect 80020 36796 80026 36808
rect 81529 36805 81541 36808
rect 81575 36805 81587 36839
rect 81529 36799 81587 36805
rect 84013 36839 84071 36845
rect 84013 36805 84025 36839
rect 84059 36836 84071 36839
rect 85482 36836 85488 36848
rect 84059 36808 85488 36836
rect 84059 36805 84071 36808
rect 84013 36799 84071 36805
rect 85482 36796 85488 36808
rect 85540 36796 85546 36848
rect 80330 36768 80336 36780
rect 79796 36740 80336 36768
rect 79796 36709 79824 36740
rect 80330 36728 80336 36740
rect 80388 36728 80394 36780
rect 85776 36768 85804 36867
rect 85942 36864 85948 36876
rect 86000 36864 86006 36916
rect 86221 36907 86279 36913
rect 86221 36873 86233 36907
rect 86267 36904 86279 36907
rect 86586 36904 86592 36916
rect 86267 36876 86592 36904
rect 86267 36873 86279 36876
rect 86221 36867 86279 36873
rect 86586 36864 86592 36876
rect 86644 36864 86650 36916
rect 86770 36864 86776 36916
rect 86828 36904 86834 36916
rect 86828 36876 87000 36904
rect 86828 36864 86834 36876
rect 86681 36771 86739 36777
rect 86681 36768 86693 36771
rect 85776 36740 86693 36768
rect 86681 36737 86693 36740
rect 86727 36737 86739 36771
rect 86972 36768 87000 36876
rect 87233 36771 87291 36777
rect 87233 36768 87245 36771
rect 86972 36740 87245 36768
rect 86681 36731 86739 36737
rect 87233 36737 87245 36740
rect 87279 36737 87291 36771
rect 87233 36731 87291 36737
rect 78677 36703 78735 36709
rect 78677 36669 78689 36703
rect 78723 36669 78735 36703
rect 78677 36663 78735 36669
rect 79781 36703 79839 36709
rect 79781 36669 79793 36703
rect 79827 36669 79839 36703
rect 79781 36663 79839 36669
rect 79965 36703 80023 36709
rect 79965 36669 79977 36703
rect 80011 36700 80023 36703
rect 80425 36703 80483 36709
rect 80425 36700 80437 36703
rect 80011 36672 80437 36700
rect 80011 36669 80023 36672
rect 79965 36663 80023 36669
rect 80425 36669 80437 36672
rect 80471 36669 80483 36703
rect 81434 36700 81440 36712
rect 81395 36672 81440 36700
rect 80425 36663 80483 36669
rect 72786 36592 72792 36644
rect 72844 36632 72850 36644
rect 72844 36604 76236 36632
rect 72844 36592 72850 36604
rect 72697 36567 72755 36573
rect 72697 36533 72709 36567
rect 72743 36564 72755 36567
rect 73338 36564 73344 36576
rect 72743 36536 73344 36564
rect 72743 36533 72755 36536
rect 72697 36527 72755 36533
rect 73338 36524 73344 36536
rect 73396 36524 73402 36576
rect 74994 36524 75000 36576
rect 75052 36564 75058 36576
rect 76101 36567 76159 36573
rect 76101 36564 76113 36567
rect 75052 36536 76113 36564
rect 75052 36524 75058 36536
rect 76101 36533 76113 36536
rect 76147 36533 76159 36567
rect 76208 36564 76236 36604
rect 79686 36592 79692 36644
rect 79744 36632 79750 36644
rect 79980 36632 80008 36663
rect 81434 36660 81440 36672
rect 81492 36660 81498 36712
rect 81713 36703 81771 36709
rect 81713 36669 81725 36703
rect 81759 36700 81771 36703
rect 84076 36703 84134 36709
rect 81759 36672 83872 36700
rect 81759 36669 81771 36672
rect 81713 36663 81771 36669
rect 79744 36604 80008 36632
rect 83737 36635 83795 36641
rect 79744 36592 79750 36604
rect 83737 36601 83749 36635
rect 83783 36601 83795 36635
rect 83844 36632 83872 36672
rect 84076 36669 84088 36703
rect 84122 36700 84134 36703
rect 86773 36703 86831 36709
rect 84122 36672 85068 36700
rect 84122 36669 84134 36672
rect 84076 36663 84134 36669
rect 84473 36635 84531 36641
rect 84473 36632 84485 36635
rect 83844 36604 84485 36632
rect 83737 36595 83795 36601
rect 84473 36601 84485 36604
rect 84519 36601 84531 36635
rect 84473 36595 84531 36601
rect 81897 36567 81955 36573
rect 81897 36564 81909 36567
rect 76208 36536 81909 36564
rect 76101 36527 76159 36533
rect 81897 36533 81909 36536
rect 81943 36533 81955 36567
rect 83752 36564 83780 36595
rect 84102 36564 84108 36576
rect 83752 36536 84108 36564
rect 81897 36527 81955 36533
rect 84102 36524 84108 36536
rect 84160 36564 84166 36576
rect 85040 36573 85068 36672
rect 86773 36669 86785 36703
rect 86819 36669 86831 36703
rect 86773 36663 86831 36669
rect 86788 36632 86816 36663
rect 86954 36660 86960 36712
rect 87012 36700 87018 36712
rect 87141 36703 87199 36709
rect 87141 36700 87153 36703
rect 87012 36672 87153 36700
rect 87012 36660 87018 36672
rect 87141 36669 87153 36672
rect 87187 36669 87199 36703
rect 88153 36703 88211 36709
rect 88153 36700 88165 36703
rect 87141 36663 87199 36669
rect 87984 36672 88165 36700
rect 87874 36632 87880 36644
rect 86788 36604 87880 36632
rect 87874 36592 87880 36604
rect 87932 36592 87938 36644
rect 87984 36576 88012 36672
rect 88153 36669 88165 36672
rect 88199 36669 88211 36703
rect 88426 36700 88432 36712
rect 88387 36672 88432 36700
rect 88153 36663 88211 36669
rect 88426 36660 88432 36672
rect 88484 36660 88490 36712
rect 88334 36632 88340 36644
rect 88295 36604 88340 36632
rect 88334 36592 88340 36604
rect 88392 36592 88398 36644
rect 88702 36592 88708 36644
rect 88760 36632 88766 36644
rect 88889 36635 88947 36641
rect 88889 36632 88901 36635
rect 88760 36604 88901 36632
rect 88760 36592 88766 36604
rect 88889 36601 88901 36604
rect 88935 36601 88947 36635
rect 88889 36595 88947 36601
rect 84565 36567 84623 36573
rect 84565 36564 84577 36567
rect 84160 36536 84577 36564
rect 84160 36524 84166 36536
rect 84565 36533 84577 36536
rect 84611 36533 84623 36567
rect 84565 36527 84623 36533
rect 85025 36567 85083 36573
rect 85025 36533 85037 36567
rect 85071 36564 85083 36567
rect 85298 36564 85304 36576
rect 85071 36536 85304 36564
rect 85071 36533 85083 36536
rect 85025 36527 85083 36533
rect 85298 36524 85304 36536
rect 85356 36524 85362 36576
rect 87966 36564 87972 36576
rect 87927 36536 87972 36564
rect 87966 36524 87972 36536
rect 88024 36524 88030 36576
rect 1104 36474 108008 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 81046 36474
rect 81098 36422 81110 36474
rect 81162 36422 81174 36474
rect 81226 36422 81238 36474
rect 81290 36422 108008 36474
rect 1104 36400 108008 36422
rect 4798 36320 4804 36372
rect 4856 36360 4862 36372
rect 5353 36363 5411 36369
rect 5353 36360 5365 36363
rect 4856 36332 5365 36360
rect 4856 36320 4862 36332
rect 5353 36329 5365 36332
rect 5399 36329 5411 36363
rect 5353 36323 5411 36329
rect 16485 36363 16543 36369
rect 16485 36329 16497 36363
rect 16531 36360 16543 36363
rect 16666 36360 16672 36372
rect 16531 36332 16672 36360
rect 16531 36329 16543 36332
rect 16485 36323 16543 36329
rect 16666 36320 16672 36332
rect 16724 36320 16730 36372
rect 17126 36360 17132 36372
rect 17087 36332 17132 36360
rect 17126 36320 17132 36332
rect 17184 36320 17190 36372
rect 18414 36320 18420 36372
rect 18472 36360 18478 36372
rect 24486 36360 24492 36372
rect 18472 36332 24492 36360
rect 18472 36320 18478 36332
rect 24486 36320 24492 36332
rect 24544 36320 24550 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 26804 36332 37473 36360
rect 3234 36252 3240 36304
rect 3292 36292 3298 36304
rect 26804 36292 26832 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 3292 36264 26832 36292
rect 3292 36252 3298 36264
rect 26878 36252 26884 36304
rect 26936 36252 26942 36304
rect 33873 36295 33931 36301
rect 32784 36264 33364 36292
rect 5258 36224 5264 36236
rect 5219 36196 5264 36224
rect 5258 36184 5264 36196
rect 5316 36184 5322 36236
rect 5813 36227 5871 36233
rect 5813 36193 5825 36227
rect 5859 36224 5871 36227
rect 9674 36224 9680 36236
rect 5859 36196 9680 36224
rect 5859 36193 5871 36196
rect 5813 36187 5871 36193
rect 9674 36184 9680 36196
rect 9732 36184 9738 36236
rect 15286 36224 15292 36236
rect 15247 36196 15292 36224
rect 15286 36184 15292 36196
rect 15344 36184 15350 36236
rect 16117 36227 16175 36233
rect 16117 36193 16129 36227
rect 16163 36193 16175 36227
rect 16117 36187 16175 36193
rect 15194 36116 15200 36168
rect 15252 36156 15258 36168
rect 15841 36159 15899 36165
rect 15841 36156 15853 36159
rect 15252 36128 15853 36156
rect 15252 36116 15258 36128
rect 15841 36125 15853 36128
rect 15887 36125 15899 36159
rect 16132 36156 16160 36187
rect 16206 36184 16212 36236
rect 16264 36224 16270 36236
rect 16301 36227 16359 36233
rect 16301 36224 16313 36227
rect 16264 36196 16313 36224
rect 16264 36184 16270 36196
rect 16301 36193 16313 36196
rect 16347 36193 16359 36227
rect 16301 36187 16359 36193
rect 17313 36227 17371 36233
rect 17313 36193 17325 36227
rect 17359 36224 17371 36227
rect 17494 36224 17500 36236
rect 17359 36196 17500 36224
rect 17359 36193 17371 36196
rect 17313 36187 17371 36193
rect 17494 36184 17500 36196
rect 17552 36184 17558 36236
rect 19705 36227 19763 36233
rect 19705 36193 19717 36227
rect 19751 36224 19763 36227
rect 19886 36224 19892 36236
rect 19751 36196 19892 36224
rect 19751 36193 19763 36196
rect 19705 36187 19763 36193
rect 19886 36184 19892 36196
rect 19944 36184 19950 36236
rect 21450 36184 21456 36236
rect 21508 36224 21514 36236
rect 21545 36227 21603 36233
rect 21545 36224 21557 36227
rect 21508 36196 21557 36224
rect 21508 36184 21514 36196
rect 21545 36193 21557 36196
rect 21591 36193 21603 36227
rect 21910 36224 21916 36236
rect 21871 36196 21916 36224
rect 21545 36187 21603 36193
rect 16666 36156 16672 36168
rect 16132 36128 16672 36156
rect 15841 36119 15899 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 20901 36159 20959 36165
rect 20901 36156 20913 36159
rect 19392 36128 20913 36156
rect 19392 36116 19398 36128
rect 20901 36125 20913 36128
rect 20947 36125 20959 36159
rect 20901 36119 20959 36125
rect 9766 36048 9772 36100
rect 9824 36088 9830 36100
rect 10318 36088 10324 36100
rect 9824 36060 10324 36088
rect 9824 36048 9830 36060
rect 10318 36048 10324 36060
rect 10376 36088 10382 36100
rect 19889 36091 19947 36097
rect 19889 36088 19901 36091
rect 10376 36060 19901 36088
rect 10376 36048 10382 36060
rect 19889 36057 19901 36060
rect 19935 36088 19947 36091
rect 21560 36088 21588 36187
rect 21910 36184 21916 36196
rect 21968 36224 21974 36236
rect 22189 36227 22247 36233
rect 22189 36224 22201 36227
rect 21968 36196 22201 36224
rect 21968 36184 21974 36196
rect 22189 36193 22201 36196
rect 22235 36193 22247 36227
rect 22189 36187 22247 36193
rect 22278 36184 22284 36236
rect 22336 36224 22342 36236
rect 22465 36227 22523 36233
rect 22465 36224 22477 36227
rect 22336 36196 22477 36224
rect 22336 36184 22342 36196
rect 22465 36193 22477 36196
rect 22511 36224 22523 36227
rect 26326 36224 26332 36236
rect 22511 36196 26332 36224
rect 22511 36193 22523 36196
rect 22465 36187 22523 36193
rect 26326 36184 26332 36196
rect 26384 36184 26390 36236
rect 26510 36224 26516 36236
rect 26471 36196 26516 36224
rect 26510 36184 26516 36196
rect 26568 36184 26574 36236
rect 26660 36227 26718 36233
rect 26660 36193 26672 36227
rect 26706 36224 26718 36227
rect 26896 36224 26924 36252
rect 32784 36233 32812 36264
rect 26706 36196 26924 36224
rect 32769 36227 32827 36233
rect 26706 36193 26718 36196
rect 26660 36187 26718 36193
rect 32769 36193 32781 36227
rect 32815 36193 32827 36227
rect 32769 36187 32827 36193
rect 32861 36227 32919 36233
rect 32861 36193 32873 36227
rect 32907 36224 32919 36227
rect 33134 36224 33140 36236
rect 32907 36196 33140 36224
rect 32907 36193 32919 36196
rect 32861 36187 32919 36193
rect 33134 36184 33140 36196
rect 33192 36224 33198 36236
rect 33336 36233 33364 36264
rect 33873 36261 33885 36295
rect 33919 36292 33931 36295
rect 37274 36292 37280 36304
rect 33919 36264 37280 36292
rect 33919 36261 33931 36264
rect 33873 36255 33931 36261
rect 37274 36252 37280 36264
rect 37332 36252 37338 36304
rect 33229 36227 33287 36233
rect 33229 36224 33241 36227
rect 33192 36196 33241 36224
rect 33192 36184 33198 36196
rect 33229 36193 33241 36196
rect 33275 36193 33287 36227
rect 33229 36187 33287 36193
rect 33321 36227 33379 36233
rect 33321 36193 33333 36227
rect 33367 36224 33379 36227
rect 34146 36224 34152 36236
rect 33367 36196 34152 36224
rect 33367 36193 33379 36196
rect 33321 36187 33379 36193
rect 34146 36184 34152 36196
rect 34204 36184 34210 36236
rect 37476 36224 37504 36323
rect 37642 36320 37648 36372
rect 37700 36360 37706 36372
rect 56321 36363 56379 36369
rect 56321 36360 56333 36363
rect 37700 36332 56333 36360
rect 37700 36320 37706 36332
rect 56321 36329 56333 36332
rect 56367 36360 56379 36363
rect 56505 36363 56563 36369
rect 56505 36360 56517 36363
rect 56367 36332 56517 36360
rect 56367 36329 56379 36332
rect 56321 36323 56379 36329
rect 56505 36329 56517 36332
rect 56551 36360 56563 36363
rect 68554 36360 68560 36372
rect 56551 36332 57100 36360
rect 68515 36332 68560 36360
rect 56551 36329 56563 36332
rect 56505 36323 56563 36329
rect 39025 36295 39083 36301
rect 39025 36261 39037 36295
rect 39071 36261 39083 36295
rect 47854 36292 47860 36304
rect 47815 36264 47860 36292
rect 39025 36255 39083 36261
rect 37734 36224 37740 36236
rect 37476 36196 37740 36224
rect 37734 36184 37740 36196
rect 37792 36184 37798 36236
rect 37921 36227 37979 36233
rect 37921 36193 37933 36227
rect 37967 36224 37979 36227
rect 38102 36224 38108 36236
rect 37967 36196 38108 36224
rect 37967 36193 37979 36196
rect 37921 36187 37979 36193
rect 21637 36159 21695 36165
rect 21637 36125 21649 36159
rect 21683 36125 21695 36159
rect 21637 36119 21695 36125
rect 21821 36159 21879 36165
rect 21821 36125 21833 36159
rect 21867 36125 21879 36159
rect 21821 36119 21879 36125
rect 19935 36060 21588 36088
rect 19935 36057 19947 36060
rect 19889 36051 19947 36057
rect 15105 36023 15163 36029
rect 15105 35989 15117 36023
rect 15151 36020 15163 36023
rect 15194 36020 15200 36032
rect 15151 35992 15200 36020
rect 15151 35989 15163 35992
rect 15105 35983 15163 35989
rect 15194 35980 15200 35992
rect 15252 35980 15258 36032
rect 17494 36020 17500 36032
rect 17455 35992 17500 36020
rect 17494 35980 17500 35992
rect 17552 35980 17558 36032
rect 21652 36020 21680 36119
rect 21836 36088 21864 36119
rect 24486 36116 24492 36168
rect 24544 36156 24550 36168
rect 26881 36159 26939 36165
rect 26881 36156 26893 36159
rect 24544 36128 26893 36156
rect 24544 36116 24550 36128
rect 26881 36125 26893 36128
rect 26927 36125 26939 36159
rect 37936 36156 37964 36187
rect 38102 36184 38108 36196
rect 38160 36224 38166 36236
rect 38473 36227 38531 36233
rect 38473 36224 38485 36227
rect 38160 36196 38485 36224
rect 38160 36184 38166 36196
rect 38473 36193 38485 36196
rect 38519 36193 38531 36227
rect 38473 36187 38531 36193
rect 38657 36227 38715 36233
rect 38657 36193 38669 36227
rect 38703 36224 38715 36227
rect 39040 36224 39068 36255
rect 47854 36252 47860 36264
rect 47912 36252 47918 36304
rect 48130 36292 48136 36304
rect 48091 36264 48136 36292
rect 48130 36252 48136 36264
rect 48188 36252 48194 36304
rect 52362 36252 52368 36304
rect 52420 36292 52426 36304
rect 52457 36295 52515 36301
rect 52457 36292 52469 36295
rect 52420 36264 52469 36292
rect 52420 36252 52426 36264
rect 52457 36261 52469 36264
rect 52503 36261 52515 36295
rect 52457 36255 52515 36261
rect 45465 36227 45523 36233
rect 45465 36224 45477 36227
rect 38703 36196 38884 36224
rect 39040 36196 45477 36224
rect 38703 36193 38715 36196
rect 38657 36187 38715 36193
rect 26881 36119 26939 36125
rect 26988 36128 32720 36156
rect 26988 36088 27016 36128
rect 21836 36060 27016 36088
rect 27157 36091 27215 36097
rect 27157 36057 27169 36091
rect 27203 36088 27215 36091
rect 32582 36088 32588 36100
rect 27203 36060 32588 36088
rect 27203 36057 27215 36060
rect 27157 36051 27215 36057
rect 32582 36048 32588 36060
rect 32640 36048 32646 36100
rect 32692 36088 32720 36128
rect 33980 36128 37964 36156
rect 33226 36088 33232 36100
rect 32692 36060 33232 36088
rect 33226 36048 33232 36060
rect 33284 36048 33290 36100
rect 22278 36020 22284 36032
rect 21652 35992 22284 36020
rect 22278 35980 22284 35992
rect 22336 35980 22342 36032
rect 25498 35980 25504 36032
rect 25556 36020 25562 36032
rect 25866 36020 25872 36032
rect 25556 35992 25872 36020
rect 25556 35980 25562 35992
rect 25866 35980 25872 35992
rect 25924 36020 25930 36032
rect 26237 36023 26295 36029
rect 26237 36020 26249 36023
rect 25924 35992 26249 36020
rect 25924 35980 25930 35992
rect 26237 35989 26249 35992
rect 26283 36020 26295 36023
rect 26418 36020 26424 36032
rect 26283 35992 26424 36020
rect 26283 35989 26295 35992
rect 26237 35983 26295 35989
rect 26418 35980 26424 35992
rect 26476 36020 26482 36032
rect 26789 36023 26847 36029
rect 26789 36020 26801 36023
rect 26476 35992 26801 36020
rect 26476 35980 26482 35992
rect 26789 35989 26801 35992
rect 26835 35989 26847 36023
rect 26789 35983 26847 35989
rect 32674 35980 32680 36032
rect 32732 36020 32738 36032
rect 33980 36020 34008 36128
rect 38286 36048 38292 36100
rect 38344 36088 38350 36100
rect 38856 36088 38884 36196
rect 45465 36193 45477 36196
rect 45511 36193 45523 36227
rect 45465 36187 45523 36193
rect 47765 36227 47823 36233
rect 47765 36193 47777 36227
rect 47811 36224 47823 36227
rect 48148 36224 48176 36252
rect 51350 36224 51356 36236
rect 47811 36196 48176 36224
rect 50816 36196 51356 36224
rect 47811 36193 47823 36196
rect 47765 36187 47823 36193
rect 44910 36116 44916 36168
rect 44968 36156 44974 36168
rect 50816 36165 50844 36196
rect 51350 36184 51356 36196
rect 51408 36184 51414 36236
rect 57072 36233 57100 36332
rect 68554 36320 68560 36332
rect 68612 36320 68618 36372
rect 68646 36320 68652 36372
rect 68704 36360 68710 36372
rect 74537 36363 74595 36369
rect 74537 36360 74549 36363
rect 68704 36332 74549 36360
rect 68704 36320 68710 36332
rect 74537 36329 74549 36332
rect 74583 36329 74595 36363
rect 74537 36323 74595 36329
rect 74629 36363 74687 36369
rect 74629 36329 74641 36363
rect 74675 36360 74687 36363
rect 76006 36360 76012 36372
rect 74675 36332 76012 36360
rect 74675 36329 74687 36332
rect 74629 36323 74687 36329
rect 63221 36295 63279 36301
rect 63221 36292 63233 36295
rect 61856 36264 63233 36292
rect 57057 36227 57115 36233
rect 57057 36193 57069 36227
rect 57103 36224 57115 36227
rect 57609 36227 57667 36233
rect 57609 36224 57621 36227
rect 57103 36196 57621 36224
rect 57103 36193 57115 36196
rect 57057 36187 57115 36193
rect 57609 36193 57621 36196
rect 57655 36193 57667 36227
rect 57609 36187 57667 36193
rect 57698 36184 57704 36236
rect 57756 36224 57762 36236
rect 57793 36227 57851 36233
rect 57793 36224 57805 36227
rect 57756 36196 57805 36224
rect 57756 36184 57762 36196
rect 57793 36193 57805 36196
rect 57839 36224 57851 36227
rect 61856 36224 61884 36264
rect 63221 36261 63233 36264
rect 63267 36292 63279 36295
rect 64414 36292 64420 36304
rect 63267 36264 64420 36292
rect 63267 36261 63279 36264
rect 63221 36255 63279 36261
rect 64414 36252 64420 36264
rect 64472 36252 64478 36304
rect 66990 36292 66996 36304
rect 66951 36264 66996 36292
rect 66990 36252 66996 36264
rect 67048 36252 67054 36304
rect 68572 36292 68600 36320
rect 67652 36264 68600 36292
rect 67652 36236 67680 36264
rect 57839 36196 61884 36224
rect 57839 36193 57851 36196
rect 57793 36187 57851 36193
rect 62022 36184 62028 36236
rect 62080 36224 62086 36236
rect 63129 36227 63187 36233
rect 63129 36224 63141 36227
rect 62080 36196 63141 36224
rect 62080 36184 62086 36196
rect 63129 36193 63141 36196
rect 63175 36193 63187 36227
rect 67634 36224 67640 36236
rect 67547 36196 67640 36224
rect 63129 36187 63187 36193
rect 67634 36184 67640 36196
rect 67692 36184 67698 36236
rect 68002 36224 68008 36236
rect 67915 36196 68008 36224
rect 68002 36184 68008 36196
rect 68060 36224 68066 36236
rect 71501 36227 71559 36233
rect 68060 36196 68784 36224
rect 68060 36184 68066 36196
rect 45189 36159 45247 36165
rect 45189 36156 45201 36159
rect 44968 36128 45201 36156
rect 44968 36116 44974 36128
rect 45189 36125 45201 36128
rect 45235 36156 45247 36159
rect 50801 36159 50859 36165
rect 50801 36156 50813 36159
rect 45235 36128 47164 36156
rect 45235 36125 45247 36128
rect 45189 36119 45247 36125
rect 39209 36091 39267 36097
rect 39209 36088 39221 36091
rect 38344 36060 39221 36088
rect 38344 36048 38350 36060
rect 39209 36057 39221 36060
rect 39255 36057 39267 36091
rect 47026 36088 47032 36100
rect 39209 36051 39267 36057
rect 46584 36060 47032 36088
rect 34146 36020 34152 36032
rect 32732 35992 34008 36020
rect 34059 35992 34152 36020
rect 32732 35980 32738 35992
rect 34146 35980 34152 35992
rect 34204 36020 34210 36032
rect 34241 36023 34299 36029
rect 34241 36020 34253 36023
rect 34204 35992 34253 36020
rect 34204 35980 34210 35992
rect 34241 35989 34253 35992
rect 34287 36020 34299 36023
rect 38378 36020 38384 36032
rect 34287 35992 38384 36020
rect 34287 35989 34299 35992
rect 34241 35983 34299 35989
rect 38378 35980 38384 35992
rect 38436 35980 38442 36032
rect 39224 36020 39252 36051
rect 46584 36020 46612 36060
rect 47026 36048 47032 36060
rect 47084 36048 47090 36100
rect 46750 36020 46756 36032
rect 39224 35992 46612 36020
rect 46711 35992 46756 36020
rect 46750 35980 46756 35992
rect 46808 35980 46814 36032
rect 46937 36023 46995 36029
rect 46937 35989 46949 36023
rect 46983 36020 46995 36023
rect 47136 36020 47164 36128
rect 50632 36128 50813 36156
rect 48498 36020 48504 36032
rect 46983 35992 48504 36020
rect 46983 35989 46995 35992
rect 46937 35983 46995 35989
rect 48498 35980 48504 35992
rect 48556 36020 48562 36032
rect 50632 36029 50660 36128
rect 50801 36125 50813 36128
rect 50847 36125 50859 36159
rect 50801 36119 50859 36125
rect 50982 36116 50988 36168
rect 51040 36156 51046 36168
rect 51077 36159 51135 36165
rect 51077 36156 51089 36159
rect 51040 36128 51089 36156
rect 51040 36116 51046 36128
rect 51077 36125 51089 36128
rect 51123 36125 51135 36159
rect 51077 36119 51135 36125
rect 56781 36159 56839 36165
rect 56781 36125 56793 36159
rect 56827 36156 56839 36159
rect 56873 36159 56931 36165
rect 56873 36156 56885 36159
rect 56827 36128 56885 36156
rect 56827 36125 56839 36128
rect 56781 36119 56839 36125
rect 56873 36125 56885 36128
rect 56919 36156 56931 36159
rect 56962 36156 56968 36168
rect 56919 36128 56968 36156
rect 56919 36125 56931 36128
rect 56873 36119 56931 36125
rect 56962 36116 56968 36128
rect 57020 36116 57026 36168
rect 67726 36156 67732 36168
rect 67687 36128 67732 36156
rect 67726 36116 67732 36128
rect 67784 36116 67790 36168
rect 67910 36156 67916 36168
rect 67871 36128 67916 36156
rect 67910 36116 67916 36128
rect 67968 36116 67974 36168
rect 67744 36088 67772 36116
rect 68281 36091 68339 36097
rect 68281 36088 68293 36091
rect 67744 36060 68293 36088
rect 68281 36057 68293 36060
rect 68327 36057 68339 36091
rect 68281 36051 68339 36057
rect 50617 36023 50675 36029
rect 50617 36020 50629 36023
rect 48556 35992 50629 36020
rect 48556 35980 48562 35992
rect 50617 35989 50629 35992
rect 50663 35989 50675 36023
rect 58066 36020 58072 36032
rect 58027 35992 58072 36020
rect 50617 35983 50675 35989
rect 58066 35980 58072 35992
rect 58124 35980 58130 36032
rect 62758 35980 62764 36032
rect 62816 36020 62822 36032
rect 68646 36020 68652 36032
rect 62816 35992 68652 36020
rect 62816 35980 62822 35992
rect 68646 35980 68652 35992
rect 68704 35980 68710 36032
rect 68756 36029 68784 36196
rect 71501 36193 71513 36227
rect 71547 36224 71559 36227
rect 73338 36224 73344 36236
rect 71547 36196 73344 36224
rect 71547 36193 71559 36196
rect 71501 36187 71559 36193
rect 73338 36184 73344 36196
rect 73396 36184 73402 36236
rect 74552 36224 74580 36323
rect 76006 36320 76012 36332
rect 76064 36320 76070 36372
rect 85942 36320 85948 36372
rect 86000 36360 86006 36372
rect 86589 36363 86647 36369
rect 86589 36360 86601 36363
rect 86000 36332 86601 36360
rect 86000 36320 86006 36332
rect 86589 36329 86601 36332
rect 86635 36360 86647 36363
rect 86862 36360 86868 36372
rect 86635 36332 86868 36360
rect 86635 36329 86647 36332
rect 86589 36323 86647 36329
rect 86862 36320 86868 36332
rect 86920 36360 86926 36372
rect 86920 36332 87000 36360
rect 86920 36320 86926 36332
rect 74920 36264 85804 36292
rect 74813 36227 74871 36233
rect 74813 36224 74825 36227
rect 74552 36196 74825 36224
rect 74813 36193 74825 36196
rect 74859 36193 74871 36227
rect 74813 36187 74871 36193
rect 71777 36159 71835 36165
rect 71777 36125 71789 36159
rect 71823 36156 71835 36159
rect 71958 36156 71964 36168
rect 71823 36128 71964 36156
rect 71823 36125 71835 36128
rect 71777 36119 71835 36125
rect 71958 36116 71964 36128
rect 72016 36116 72022 36168
rect 74920 36088 74948 36264
rect 75178 36184 75184 36236
rect 75236 36224 75242 36236
rect 75273 36227 75331 36233
rect 75273 36224 75285 36227
rect 75236 36196 75285 36224
rect 75236 36184 75242 36196
rect 75273 36193 75285 36196
rect 75319 36193 75331 36227
rect 75273 36187 75331 36193
rect 75362 36184 75368 36236
rect 75420 36224 75426 36236
rect 75420 36196 75465 36224
rect 75420 36184 75426 36196
rect 79870 36184 79876 36236
rect 79928 36224 79934 36236
rect 79965 36227 80023 36233
rect 79965 36224 79977 36227
rect 79928 36196 79977 36224
rect 79928 36184 79934 36196
rect 79965 36193 79977 36196
rect 80011 36193 80023 36227
rect 79965 36187 80023 36193
rect 80057 36227 80115 36233
rect 80057 36193 80069 36227
rect 80103 36224 80115 36227
rect 80422 36224 80428 36236
rect 80103 36196 80428 36224
rect 80103 36193 80115 36196
rect 80057 36187 80115 36193
rect 80422 36184 80428 36196
rect 80480 36184 80486 36236
rect 85776 36233 85804 36264
rect 85850 36252 85856 36304
rect 85908 36292 85914 36304
rect 86770 36292 86776 36304
rect 85908 36264 86776 36292
rect 85908 36252 85914 36264
rect 86770 36252 86776 36264
rect 86828 36252 86834 36304
rect 86972 36233 87000 36332
rect 87322 36292 87328 36304
rect 87283 36264 87328 36292
rect 87322 36252 87328 36264
rect 87380 36252 87386 36304
rect 85761 36227 85819 36233
rect 85761 36193 85773 36227
rect 85807 36224 85819 36227
rect 86037 36227 86095 36233
rect 86037 36224 86049 36227
rect 85807 36196 86049 36224
rect 85807 36193 85819 36196
rect 85761 36187 85819 36193
rect 86037 36193 86049 36196
rect 86083 36193 86095 36227
rect 86037 36187 86095 36193
rect 86957 36227 87015 36233
rect 86957 36193 86969 36227
rect 87003 36193 87015 36227
rect 88702 36224 88708 36236
rect 86957 36187 87015 36193
rect 88076 36196 88564 36224
rect 88663 36196 88708 36224
rect 75822 36156 75828 36168
rect 75783 36128 75828 36156
rect 75822 36116 75828 36128
rect 75880 36116 75886 36168
rect 86052 36156 86080 36187
rect 88076 36168 88104 36196
rect 88058 36156 88064 36168
rect 86052 36128 88064 36156
rect 88058 36116 88064 36128
rect 88116 36116 88122 36168
rect 88429 36159 88487 36165
rect 88429 36156 88441 36159
rect 88260 36128 88441 36156
rect 72436 36060 74948 36088
rect 75089 36091 75147 36097
rect 68741 36023 68799 36029
rect 68741 35989 68753 36023
rect 68787 36020 68799 36023
rect 72436 36020 72464 36060
rect 75089 36057 75101 36091
rect 75135 36088 75147 36091
rect 77202 36088 77208 36100
rect 75135 36060 77208 36088
rect 75135 36057 75147 36060
rect 75089 36051 75147 36057
rect 77202 36048 77208 36060
rect 77260 36048 77266 36100
rect 79796 36060 85712 36088
rect 72878 36020 72884 36032
rect 68787 35992 72464 36020
rect 72839 35992 72884 36020
rect 68787 35989 68799 35992
rect 68741 35983 68799 35989
rect 72878 35980 72884 35992
rect 72936 35980 72942 36032
rect 73338 36020 73344 36032
rect 73251 35992 73344 36020
rect 73338 35980 73344 35992
rect 73396 36020 73402 36032
rect 76650 36020 76656 36032
rect 73396 35992 76656 36020
rect 73396 35980 73402 35992
rect 76650 35980 76656 35992
rect 76708 35980 76714 36032
rect 79502 35980 79508 36032
rect 79560 36020 79566 36032
rect 79796 36029 79824 36060
rect 79597 36023 79655 36029
rect 79597 36020 79609 36023
rect 79560 35992 79609 36020
rect 79560 35980 79566 35992
rect 79597 35989 79609 35992
rect 79643 36020 79655 36023
rect 79781 36023 79839 36029
rect 79781 36020 79793 36023
rect 79643 35992 79793 36020
rect 79643 35989 79655 35992
rect 79597 35983 79655 35989
rect 79781 35989 79793 35992
rect 79827 35989 79839 36023
rect 80238 36020 80244 36032
rect 80199 35992 80244 36020
rect 79781 35983 79839 35989
rect 80238 35980 80244 35992
rect 80296 35980 80302 36032
rect 85684 36020 85712 36060
rect 85758 36048 85764 36100
rect 85816 36088 85822 36100
rect 85853 36091 85911 36097
rect 85853 36088 85865 36091
rect 85816 36060 85865 36088
rect 85816 36048 85822 36060
rect 85853 36057 85865 36060
rect 85899 36057 85911 36091
rect 87966 36088 87972 36100
rect 85853 36051 85911 36057
rect 86236 36060 87972 36088
rect 86236 36020 86264 36060
rect 87966 36048 87972 36060
rect 88024 36048 88030 36100
rect 85684 35992 86264 36020
rect 86310 35980 86316 36032
rect 86368 36020 86374 36032
rect 88260 36029 88288 36128
rect 88429 36125 88441 36128
rect 88475 36125 88487 36159
rect 88536 36156 88564 36196
rect 88702 36184 88708 36196
rect 88760 36184 88766 36236
rect 88536 36128 89392 36156
rect 88429 36119 88487 36125
rect 88245 36023 88303 36029
rect 88245 36020 88257 36023
rect 86368 35992 88257 36020
rect 86368 35980 86374 35992
rect 88245 35989 88257 35992
rect 88291 35989 88303 36023
rect 89364 36020 89392 36128
rect 89809 36023 89867 36029
rect 89809 36020 89821 36023
rect 89364 35992 89821 36020
rect 88245 35983 88303 35989
rect 89809 35989 89821 35992
rect 89855 35989 89867 36023
rect 89809 35983 89867 35989
rect 1104 35930 108008 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 65686 35930
rect 65738 35878 65750 35930
rect 65802 35878 65814 35930
rect 65866 35878 65878 35930
rect 65930 35878 96406 35930
rect 96458 35878 96470 35930
rect 96522 35878 96534 35930
rect 96586 35878 96598 35930
rect 96650 35878 108008 35930
rect 1104 35856 108008 35878
rect 4062 35776 4068 35828
rect 4120 35816 4126 35828
rect 17770 35816 17776 35828
rect 4120 35788 17776 35816
rect 4120 35776 4126 35788
rect 17770 35776 17776 35788
rect 17828 35776 17834 35828
rect 17862 35776 17868 35828
rect 17920 35816 17926 35828
rect 20622 35816 20628 35828
rect 17920 35788 20628 35816
rect 17920 35776 17926 35788
rect 20622 35776 20628 35788
rect 20680 35776 20686 35828
rect 21637 35819 21695 35825
rect 21637 35785 21649 35819
rect 21683 35816 21695 35819
rect 21910 35816 21916 35828
rect 21683 35788 21916 35816
rect 21683 35785 21695 35788
rect 21637 35779 21695 35785
rect 21910 35776 21916 35788
rect 21968 35776 21974 35828
rect 26050 35776 26056 35828
rect 26108 35816 26114 35828
rect 26145 35819 26203 35825
rect 26145 35816 26157 35819
rect 26108 35788 26157 35816
rect 26108 35776 26114 35788
rect 26145 35785 26157 35788
rect 26191 35785 26203 35819
rect 26145 35779 26203 35785
rect 26694 35776 26700 35828
rect 26752 35816 26758 35828
rect 38286 35816 38292 35828
rect 26752 35788 38292 35816
rect 26752 35776 26758 35788
rect 38286 35776 38292 35788
rect 38344 35776 38350 35828
rect 38378 35776 38384 35828
rect 38436 35816 38442 35828
rect 62758 35816 62764 35828
rect 38436 35788 62764 35816
rect 38436 35776 38442 35788
rect 62758 35776 62764 35788
rect 62816 35776 62822 35828
rect 65978 35776 65984 35828
rect 66036 35816 66042 35828
rect 66073 35819 66131 35825
rect 66073 35816 66085 35819
rect 66036 35788 66085 35816
rect 66036 35776 66042 35788
rect 66073 35785 66085 35788
rect 66119 35785 66131 35819
rect 66073 35779 66131 35785
rect 66806 35776 66812 35828
rect 66864 35816 66870 35828
rect 67361 35819 67419 35825
rect 67361 35816 67373 35819
rect 66864 35788 67373 35816
rect 66864 35776 66870 35788
rect 67361 35785 67373 35788
rect 67407 35816 67419 35819
rect 68002 35816 68008 35828
rect 67407 35788 68008 35816
rect 67407 35785 67419 35788
rect 67361 35779 67419 35785
rect 68002 35776 68008 35788
rect 68060 35776 68066 35828
rect 71682 35776 71688 35828
rect 71740 35816 71746 35828
rect 72237 35819 72295 35825
rect 72237 35816 72249 35819
rect 71740 35788 72249 35816
rect 71740 35776 71746 35788
rect 72237 35785 72249 35788
rect 72283 35785 72295 35819
rect 72237 35779 72295 35785
rect 75914 35776 75920 35828
rect 75972 35816 75978 35828
rect 76929 35819 76987 35825
rect 76929 35816 76941 35819
rect 75972 35788 76941 35816
rect 75972 35776 75978 35788
rect 76929 35785 76941 35788
rect 76975 35816 76987 35819
rect 77018 35816 77024 35828
rect 76975 35788 77024 35816
rect 76975 35785 76987 35788
rect 76929 35779 76987 35785
rect 77018 35776 77024 35788
rect 77076 35776 77082 35828
rect 81342 35816 81348 35828
rect 81303 35788 81348 35816
rect 81342 35776 81348 35788
rect 81400 35776 81406 35828
rect 5994 35748 6000 35760
rect 5955 35720 6000 35748
rect 5994 35708 6000 35720
rect 6052 35708 6058 35760
rect 9398 35708 9404 35760
rect 9456 35748 9462 35760
rect 27614 35748 27620 35760
rect 9456 35720 27620 35748
rect 9456 35708 9462 35720
rect 27614 35708 27620 35720
rect 27672 35708 27678 35760
rect 29362 35708 29368 35760
rect 29420 35748 29426 35760
rect 29457 35751 29515 35757
rect 29457 35748 29469 35751
rect 29420 35720 29469 35748
rect 29420 35708 29426 35720
rect 29457 35717 29469 35720
rect 29503 35717 29515 35751
rect 29457 35711 29515 35717
rect 32232 35720 33180 35748
rect 2590 35680 2596 35692
rect 2551 35652 2596 35680
rect 2590 35640 2596 35652
rect 2648 35640 2654 35692
rect 2869 35683 2927 35689
rect 2869 35649 2881 35683
rect 2915 35680 2927 35683
rect 3050 35680 3056 35692
rect 2915 35652 3056 35680
rect 2915 35649 2927 35652
rect 2869 35643 2927 35649
rect 3050 35640 3056 35652
rect 3108 35640 3114 35692
rect 4890 35640 4896 35692
rect 4948 35680 4954 35692
rect 5258 35680 5264 35692
rect 4948 35652 5264 35680
rect 4948 35640 4954 35652
rect 5258 35640 5264 35652
rect 5316 35680 5322 35692
rect 5316 35652 5396 35680
rect 5316 35640 5322 35652
rect 2608 35612 2636 35640
rect 4341 35615 4399 35621
rect 4341 35612 4353 35615
rect 2608 35584 4353 35612
rect 4341 35581 4353 35584
rect 4387 35612 4399 35615
rect 4706 35612 4712 35624
rect 4387 35584 4712 35612
rect 4387 35581 4399 35584
rect 4341 35575 4399 35581
rect 4706 35572 4712 35584
rect 4764 35612 4770 35624
rect 5368 35621 5396 35652
rect 5353 35615 5411 35621
rect 4764 35584 5304 35612
rect 4764 35572 4770 35584
rect 5276 35544 5304 35584
rect 5353 35581 5365 35615
rect 5399 35581 5411 35615
rect 5353 35575 5411 35581
rect 5629 35615 5687 35621
rect 5629 35581 5641 35615
rect 5675 35612 5687 35615
rect 6012 35612 6040 35708
rect 8665 35683 8723 35689
rect 8665 35649 8677 35683
rect 8711 35680 8723 35683
rect 13630 35680 13636 35692
rect 8711 35652 13636 35680
rect 8711 35649 8723 35652
rect 8665 35643 8723 35649
rect 13630 35640 13636 35652
rect 13688 35640 13694 35692
rect 16022 35680 16028 35692
rect 14108 35652 16028 35680
rect 5675 35584 6040 35612
rect 8389 35615 8447 35621
rect 5675 35581 5687 35584
rect 5629 35575 5687 35581
rect 8389 35581 8401 35615
rect 8435 35612 8447 35615
rect 9306 35612 9312 35624
rect 8435 35584 9312 35612
rect 8435 35581 8447 35584
rect 8389 35575 8447 35581
rect 8404 35544 8432 35575
rect 9306 35572 9312 35584
rect 9364 35612 9370 35624
rect 10137 35615 10195 35621
rect 10137 35612 10149 35615
rect 9364 35584 10149 35612
rect 9364 35572 9370 35584
rect 10137 35581 10149 35584
rect 10183 35581 10195 35615
rect 13357 35615 13415 35621
rect 13357 35612 13369 35615
rect 10137 35575 10195 35581
rect 12360 35584 13369 35612
rect 12360 35544 12388 35584
rect 13357 35581 13369 35584
rect 13403 35612 13415 35615
rect 13538 35612 13544 35624
rect 13403 35584 13544 35612
rect 13403 35581 13415 35584
rect 13357 35575 13415 35581
rect 13538 35572 13544 35584
rect 13596 35572 13602 35624
rect 14108 35621 14136 35652
rect 16022 35640 16028 35652
rect 16080 35640 16086 35692
rect 16577 35683 16635 35689
rect 16577 35680 16589 35683
rect 16132 35652 16589 35680
rect 16132 35624 16160 35652
rect 16577 35649 16589 35652
rect 16623 35680 16635 35683
rect 21082 35680 21088 35692
rect 16623 35652 21088 35680
rect 16623 35649 16635 35652
rect 16577 35643 16635 35649
rect 21082 35640 21088 35652
rect 21140 35640 21146 35692
rect 21818 35640 21824 35692
rect 21876 35680 21882 35692
rect 31938 35680 31944 35692
rect 21876 35652 31944 35680
rect 21876 35640 21882 35652
rect 31938 35640 31944 35652
rect 31996 35640 32002 35692
rect 14093 35615 14151 35621
rect 14093 35581 14105 35615
rect 14139 35581 14151 35615
rect 14093 35575 14151 35581
rect 14369 35615 14427 35621
rect 14369 35581 14381 35615
rect 14415 35612 14427 35615
rect 15289 35615 15347 35621
rect 15289 35612 15301 35615
rect 14415 35584 15301 35612
rect 14415 35581 14427 35584
rect 14369 35575 14427 35581
rect 15289 35581 15301 35584
rect 15335 35581 15347 35615
rect 15289 35575 15347 35581
rect 15841 35615 15899 35621
rect 15841 35581 15853 35615
rect 15887 35581 15899 35615
rect 16114 35612 16120 35624
rect 16075 35584 16120 35612
rect 15841 35575 15899 35581
rect 3528 35516 5212 35544
rect 5276 35516 8432 35544
rect 9692 35516 12388 35544
rect 3142 35436 3148 35488
rect 3200 35476 3206 35488
rect 3528 35476 3556 35516
rect 4154 35476 4160 35488
rect 3200 35448 3556 35476
rect 4115 35448 4160 35476
rect 3200 35436 3206 35448
rect 4154 35436 4160 35448
rect 4212 35436 4218 35488
rect 5184 35485 5212 35516
rect 5169 35479 5227 35485
rect 5169 35445 5181 35479
rect 5215 35445 5227 35479
rect 5169 35439 5227 35445
rect 7282 35436 7288 35488
rect 7340 35476 7346 35488
rect 9692 35476 9720 35516
rect 12710 35504 12716 35556
rect 12768 35544 12774 35556
rect 15194 35544 15200 35556
rect 12768 35516 15200 35544
rect 12768 35504 12774 35516
rect 15194 35504 15200 35516
rect 15252 35544 15258 35556
rect 15856 35544 15884 35575
rect 16114 35572 16120 35584
rect 16172 35572 16178 35624
rect 16301 35615 16359 35621
rect 16301 35581 16313 35615
rect 16347 35612 16359 35615
rect 16347 35584 16528 35612
rect 16347 35581 16359 35584
rect 16301 35575 16359 35581
rect 15252 35516 15884 35544
rect 15252 35504 15258 35516
rect 16500 35488 16528 35584
rect 19886 35572 19892 35624
rect 19944 35612 19950 35624
rect 20349 35615 20407 35621
rect 20349 35612 20361 35615
rect 19944 35584 20361 35612
rect 19944 35572 19950 35584
rect 20349 35581 20361 35584
rect 20395 35581 20407 35615
rect 20349 35575 20407 35581
rect 21358 35572 21364 35624
rect 21416 35612 21422 35624
rect 21453 35615 21511 35621
rect 21453 35612 21465 35615
rect 21416 35584 21465 35612
rect 21416 35572 21422 35584
rect 21453 35581 21465 35584
rect 21499 35612 21511 35615
rect 21913 35615 21971 35621
rect 21913 35612 21925 35615
rect 21499 35584 21925 35612
rect 21499 35581 21511 35584
rect 21453 35575 21511 35581
rect 21913 35581 21925 35584
rect 21959 35581 21971 35615
rect 26326 35612 26332 35624
rect 26287 35584 26332 35612
rect 21913 35575 21971 35581
rect 26326 35572 26332 35584
rect 26384 35572 26390 35624
rect 26513 35615 26571 35621
rect 26513 35581 26525 35615
rect 26559 35612 26571 35615
rect 26602 35612 26608 35624
rect 26559 35584 26608 35612
rect 26559 35581 26571 35584
rect 26513 35575 26571 35581
rect 26602 35572 26608 35584
rect 26660 35572 26666 35624
rect 26878 35612 26884 35624
rect 26839 35584 26884 35612
rect 26878 35572 26884 35584
rect 26936 35572 26942 35624
rect 26973 35615 27031 35621
rect 26973 35581 26985 35615
rect 27019 35581 27031 35615
rect 26973 35575 27031 35581
rect 16666 35504 16672 35556
rect 16724 35544 16730 35556
rect 24762 35544 24768 35556
rect 16724 35516 24768 35544
rect 16724 35504 16730 35516
rect 24762 35504 24768 35516
rect 24820 35504 24826 35556
rect 26234 35504 26240 35556
rect 26292 35544 26298 35556
rect 26988 35544 27016 35575
rect 27062 35572 27068 35624
rect 27120 35612 27126 35624
rect 29273 35615 29331 35621
rect 29273 35612 29285 35615
rect 27120 35584 29285 35612
rect 27120 35572 27126 35584
rect 29273 35581 29285 35584
rect 29319 35581 29331 35615
rect 32030 35612 32036 35624
rect 31991 35584 32036 35612
rect 29273 35575 29331 35581
rect 26292 35516 27016 35544
rect 26292 35504 26298 35516
rect 27246 35504 27252 35556
rect 27304 35544 27310 35556
rect 29288 35544 29316 35575
rect 32030 35572 32036 35584
rect 32088 35572 32094 35624
rect 32232 35621 32260 35720
rect 32217 35615 32275 35621
rect 32217 35581 32229 35615
rect 32263 35581 32275 35615
rect 32217 35575 32275 35581
rect 32582 35572 32588 35624
rect 32640 35612 32646 35624
rect 32677 35615 32735 35621
rect 32677 35612 32689 35615
rect 32640 35584 32689 35612
rect 32640 35572 32646 35584
rect 32677 35581 32689 35584
rect 32723 35581 32735 35615
rect 32677 35575 32735 35581
rect 32769 35615 32827 35621
rect 32769 35581 32781 35615
rect 32815 35612 32827 35615
rect 33152 35612 33180 35720
rect 38838 35708 38844 35760
rect 38896 35748 38902 35760
rect 47026 35748 47032 35760
rect 38896 35720 44128 35748
rect 46987 35720 47032 35748
rect 38896 35708 38902 35720
rect 33321 35683 33379 35689
rect 33321 35649 33333 35683
rect 33367 35680 33379 35683
rect 41230 35680 41236 35692
rect 33367 35652 41236 35680
rect 33367 35649 33379 35652
rect 33321 35643 33379 35649
rect 41230 35640 41236 35652
rect 41288 35640 41294 35692
rect 33965 35615 34023 35621
rect 33965 35612 33977 35615
rect 32815 35584 33977 35612
rect 32815 35581 32827 35584
rect 32769 35575 32827 35581
rect 33965 35581 33977 35584
rect 34011 35612 34023 35615
rect 34146 35612 34152 35624
rect 34011 35584 34152 35612
rect 34011 35581 34023 35584
rect 33965 35575 34023 35581
rect 34146 35572 34152 35584
rect 34204 35572 34210 35624
rect 37366 35572 37372 35624
rect 37424 35612 37430 35624
rect 42797 35615 42855 35621
rect 42797 35612 42809 35615
rect 37424 35584 42809 35612
rect 37424 35572 37430 35584
rect 42797 35581 42809 35584
rect 42843 35612 42855 35615
rect 42981 35615 43039 35621
rect 42981 35612 42993 35615
rect 42843 35584 42993 35612
rect 42843 35581 42855 35584
rect 42797 35575 42855 35581
rect 42981 35581 42993 35584
rect 43027 35581 43039 35615
rect 42981 35575 43039 35581
rect 43165 35615 43223 35621
rect 43165 35581 43177 35615
rect 43211 35581 43223 35615
rect 43714 35612 43720 35624
rect 43675 35584 43720 35612
rect 43165 35575 43223 35581
rect 29733 35547 29791 35553
rect 29733 35544 29745 35547
rect 27304 35516 27476 35544
rect 29288 35516 29745 35544
rect 27304 35504 27310 35516
rect 7340 35448 9720 35476
rect 9769 35479 9827 35485
rect 7340 35436 7346 35448
rect 9769 35445 9781 35479
rect 9815 35476 9827 35479
rect 9858 35476 9864 35488
rect 9815 35448 9864 35476
rect 9815 35445 9827 35448
rect 9769 35439 9827 35445
rect 9858 35436 9864 35448
rect 9916 35436 9922 35488
rect 13446 35476 13452 35488
rect 13407 35448 13452 35476
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 16482 35476 16488 35488
rect 16443 35448 16488 35476
rect 16482 35436 16488 35448
rect 16540 35436 16546 35488
rect 16758 35436 16764 35488
rect 16816 35476 16822 35488
rect 20530 35476 20536 35488
rect 16816 35448 20536 35476
rect 16816 35436 16822 35448
rect 20530 35436 20536 35448
rect 20588 35436 20594 35488
rect 20622 35436 20628 35488
rect 20680 35476 20686 35488
rect 27062 35476 27068 35488
rect 20680 35448 27068 35476
rect 20680 35436 20686 35448
rect 27062 35436 27068 35448
rect 27120 35436 27126 35488
rect 27154 35436 27160 35488
rect 27212 35476 27218 35488
rect 27448 35485 27476 35516
rect 29733 35513 29745 35516
rect 29779 35544 29791 35547
rect 42426 35544 42432 35556
rect 29779 35516 42432 35544
rect 29779 35513 29791 35516
rect 29733 35507 29791 35513
rect 42426 35504 42432 35516
rect 42484 35504 42490 35556
rect 27433 35479 27491 35485
rect 27212 35448 27257 35476
rect 27212 35436 27218 35448
rect 27433 35445 27445 35479
rect 27479 35476 27491 35479
rect 28074 35476 28080 35488
rect 27479 35448 28080 35476
rect 27479 35445 27491 35448
rect 27433 35439 27491 35445
rect 28074 35436 28080 35448
rect 28132 35436 28138 35488
rect 33502 35476 33508 35488
rect 33463 35448 33508 35476
rect 33502 35436 33508 35448
rect 33560 35476 33566 35488
rect 33689 35479 33747 35485
rect 33689 35476 33701 35479
rect 33560 35448 33701 35476
rect 33560 35436 33566 35448
rect 33689 35445 33701 35448
rect 33735 35445 33747 35479
rect 33689 35439 33747 35445
rect 33778 35436 33784 35488
rect 33836 35476 33842 35488
rect 39758 35476 39764 35488
rect 33836 35448 39764 35476
rect 33836 35436 33842 35448
rect 39758 35436 39764 35448
rect 39816 35436 39822 35488
rect 43180 35476 43208 35575
rect 43714 35572 43720 35584
rect 43772 35572 43778 35624
rect 43901 35615 43959 35621
rect 43901 35581 43913 35615
rect 43947 35612 43959 35615
rect 44100 35612 44128 35720
rect 47026 35708 47032 35720
rect 47084 35708 47090 35760
rect 51166 35708 51172 35760
rect 51224 35748 51230 35760
rect 51902 35748 51908 35760
rect 51224 35720 51908 35748
rect 51224 35708 51230 35720
rect 51902 35708 51908 35720
rect 51960 35748 51966 35760
rect 51997 35751 52055 35757
rect 51997 35748 52009 35751
rect 51960 35720 52009 35748
rect 51960 35708 51966 35720
rect 51997 35717 52009 35720
rect 52043 35717 52055 35751
rect 51997 35711 52055 35717
rect 44269 35683 44327 35689
rect 44269 35649 44281 35683
rect 44315 35680 44327 35683
rect 45186 35680 45192 35692
rect 44315 35652 45192 35680
rect 44315 35649 44327 35652
rect 44269 35643 44327 35649
rect 45186 35640 45192 35652
rect 45244 35640 45250 35692
rect 46750 35640 46756 35692
rect 46808 35680 46814 35692
rect 46845 35683 46903 35689
rect 46845 35680 46857 35683
rect 46808 35652 46857 35680
rect 46808 35640 46814 35652
rect 46845 35649 46857 35652
rect 46891 35680 46903 35683
rect 57054 35680 57060 35692
rect 46891 35652 57060 35680
rect 46891 35649 46903 35652
rect 46845 35643 46903 35649
rect 46198 35612 46204 35624
rect 43947 35584 46204 35612
rect 43947 35581 43959 35584
rect 43901 35575 43959 35581
rect 46198 35572 46204 35584
rect 46256 35572 46262 35624
rect 46952 35621 46980 35652
rect 57054 35640 57060 35652
rect 57112 35640 57118 35692
rect 58066 35640 58072 35692
rect 58124 35680 58130 35692
rect 58713 35683 58771 35689
rect 58713 35680 58725 35683
rect 58124 35652 58725 35680
rect 58124 35640 58130 35652
rect 58713 35649 58725 35652
rect 58759 35649 58771 35683
rect 58713 35643 58771 35649
rect 60093 35683 60151 35689
rect 60093 35649 60105 35683
rect 60139 35680 60151 35683
rect 62022 35680 62028 35692
rect 60139 35652 62028 35680
rect 60139 35649 60151 35652
rect 60093 35643 60151 35649
rect 62022 35640 62028 35652
rect 62080 35640 62086 35692
rect 67177 35683 67235 35689
rect 67177 35680 67189 35683
rect 66456 35652 67189 35680
rect 46937 35615 46995 35621
rect 46937 35581 46949 35615
rect 46983 35581 46995 35615
rect 46937 35575 46995 35581
rect 51905 35615 51963 35621
rect 51905 35581 51917 35615
rect 51951 35612 51963 35615
rect 53098 35612 53104 35624
rect 51951 35584 53104 35612
rect 51951 35581 51963 35584
rect 51905 35575 51963 35581
rect 53098 35572 53104 35584
rect 53156 35572 53162 35624
rect 58437 35615 58495 35621
rect 58437 35581 58449 35615
rect 58483 35581 58495 35615
rect 63126 35612 63132 35624
rect 63087 35584 63132 35612
rect 58437 35575 58495 35581
rect 43530 35504 43536 35556
rect 43588 35544 43594 35556
rect 49694 35544 49700 35556
rect 43588 35516 49700 35544
rect 43588 35504 43594 35516
rect 49694 35504 49700 35516
rect 49752 35504 49758 35556
rect 56594 35504 56600 35556
rect 56652 35544 56658 35556
rect 56870 35544 56876 35556
rect 56652 35516 56876 35544
rect 56652 35504 56658 35516
rect 56870 35504 56876 35516
rect 56928 35504 56934 35556
rect 43254 35476 43260 35488
rect 43180 35448 43260 35476
rect 43254 35436 43260 35448
rect 43312 35436 43318 35488
rect 44358 35436 44364 35488
rect 44416 35476 44422 35488
rect 44453 35479 44511 35485
rect 44453 35476 44465 35479
rect 44416 35448 44465 35476
rect 44416 35436 44422 35448
rect 44453 35445 44465 35448
rect 44499 35445 44511 35479
rect 58452 35476 58480 35575
rect 63126 35572 63132 35584
rect 63184 35572 63190 35624
rect 66456 35621 66484 35652
rect 67177 35649 67189 35652
rect 67223 35680 67235 35683
rect 67634 35680 67640 35692
rect 67223 35652 67640 35680
rect 67223 35649 67235 35652
rect 67177 35643 67235 35649
rect 67634 35640 67640 35652
rect 67692 35640 67698 35692
rect 71409 35683 71467 35689
rect 71409 35649 71421 35683
rect 71455 35680 71467 35683
rect 71700 35680 71728 35776
rect 85482 35748 85488 35760
rect 85443 35720 85488 35748
rect 85482 35708 85488 35720
rect 85540 35708 85546 35760
rect 71958 35680 71964 35692
rect 71455 35652 71728 35680
rect 71919 35652 71964 35680
rect 71455 35649 71467 35652
rect 71409 35643 71467 35649
rect 71958 35640 71964 35652
rect 72016 35640 72022 35692
rect 74721 35683 74779 35689
rect 74721 35649 74733 35683
rect 74767 35680 74779 35683
rect 75362 35680 75368 35692
rect 74767 35652 75368 35680
rect 74767 35649 74779 35652
rect 74721 35643 74779 35649
rect 75362 35640 75368 35652
rect 75420 35640 75426 35692
rect 75822 35680 75828 35692
rect 75783 35652 75828 35680
rect 75822 35640 75828 35652
rect 75880 35640 75886 35692
rect 80057 35683 80115 35689
rect 80057 35649 80069 35683
rect 80103 35680 80115 35683
rect 80238 35680 80244 35692
rect 80103 35652 80244 35680
rect 80103 35649 80115 35652
rect 80057 35643 80115 35649
rect 80238 35640 80244 35652
rect 80296 35640 80302 35692
rect 85298 35640 85304 35692
rect 85356 35680 85362 35692
rect 85850 35680 85856 35692
rect 85356 35652 85712 35680
rect 85811 35652 85856 35680
rect 85356 35640 85362 35652
rect 66257 35615 66315 35621
rect 66257 35612 66269 35615
rect 65628 35584 66269 35612
rect 59446 35476 59452 35488
rect 58452 35448 59452 35476
rect 44453 35439 44511 35445
rect 59446 35436 59452 35448
rect 59504 35476 59510 35488
rect 60185 35479 60243 35485
rect 60185 35476 60197 35479
rect 59504 35448 60197 35476
rect 59504 35436 59510 35448
rect 60185 35445 60197 35448
rect 60231 35476 60243 35479
rect 60918 35476 60924 35488
rect 60231 35448 60924 35476
rect 60231 35445 60243 35448
rect 60185 35439 60243 35445
rect 60918 35436 60924 35448
rect 60976 35436 60982 35488
rect 63218 35476 63224 35488
rect 63179 35448 63224 35476
rect 63218 35436 63224 35448
rect 63276 35436 63282 35488
rect 65518 35436 65524 35488
rect 65576 35476 65582 35488
rect 65628 35485 65656 35584
rect 66257 35581 66269 35584
rect 66303 35581 66315 35615
rect 66257 35575 66315 35581
rect 66441 35615 66499 35621
rect 66441 35581 66453 35615
rect 66487 35581 66499 35615
rect 66806 35612 66812 35624
rect 66767 35584 66812 35612
rect 66441 35575 66499 35581
rect 66806 35572 66812 35584
rect 66864 35572 66870 35624
rect 66901 35615 66959 35621
rect 66901 35581 66913 35615
rect 66947 35581 66959 35615
rect 66901 35575 66959 35581
rect 71501 35615 71559 35621
rect 71501 35581 71513 35615
rect 71547 35612 71559 35615
rect 72142 35612 72148 35624
rect 71547 35584 72148 35612
rect 71547 35581 71559 35584
rect 71501 35575 71559 35581
rect 65978 35504 65984 35556
rect 66036 35544 66042 35556
rect 66916 35544 66944 35575
rect 72142 35572 72148 35584
rect 72200 35572 72206 35624
rect 72878 35572 72884 35624
rect 72936 35612 72942 35624
rect 74353 35615 74411 35621
rect 74353 35612 74365 35615
rect 72936 35584 74365 35612
rect 72936 35572 72942 35584
rect 74353 35581 74365 35584
rect 74399 35612 74411 35615
rect 74813 35615 74871 35621
rect 74813 35612 74825 35615
rect 74399 35584 74825 35612
rect 74399 35581 74411 35584
rect 74353 35575 74411 35581
rect 74813 35581 74825 35584
rect 74859 35581 74871 35615
rect 74813 35575 74871 35581
rect 75549 35615 75607 35621
rect 75549 35581 75561 35615
rect 75595 35581 75607 35615
rect 79781 35615 79839 35621
rect 79781 35612 79793 35615
rect 75549 35575 75607 35581
rect 79520 35584 79793 35612
rect 66036 35516 66944 35544
rect 66036 35504 66042 35516
rect 74166 35504 74172 35556
rect 74224 35544 74230 35556
rect 74224 35516 74266 35544
rect 74224 35504 74230 35516
rect 65613 35479 65671 35485
rect 65613 35476 65625 35479
rect 65576 35448 65625 35476
rect 65576 35436 65582 35448
rect 65613 35445 65625 35448
rect 65659 35445 65671 35479
rect 72142 35476 72148 35488
rect 72103 35448 72148 35476
rect 65613 35439 65671 35445
rect 72142 35436 72148 35448
rect 72200 35436 72206 35488
rect 74184 35476 74212 35504
rect 74994 35476 75000 35488
rect 74184 35448 75000 35476
rect 74994 35436 75000 35448
rect 75052 35436 75058 35488
rect 75564 35476 75592 35575
rect 77294 35476 77300 35488
rect 75564 35448 77300 35476
rect 77294 35436 77300 35448
rect 77352 35476 77358 35488
rect 79520 35485 79548 35584
rect 79781 35581 79793 35584
rect 79827 35581 79839 35615
rect 79781 35575 79839 35581
rect 81434 35572 81440 35624
rect 81492 35612 81498 35624
rect 85684 35621 85712 35652
rect 85850 35640 85856 35652
rect 85908 35640 85914 35692
rect 88334 35680 88340 35692
rect 88295 35652 88340 35680
rect 88334 35640 88340 35652
rect 88392 35640 88398 35692
rect 85393 35615 85451 35621
rect 85393 35612 85405 35615
rect 81492 35584 85405 35612
rect 81492 35572 81498 35584
rect 85393 35581 85405 35584
rect 85439 35581 85451 35615
rect 85393 35575 85451 35581
rect 85669 35615 85727 35621
rect 85669 35581 85681 35615
rect 85715 35612 85727 35615
rect 86221 35615 86279 35621
rect 86221 35612 86233 35615
rect 85715 35584 86233 35612
rect 85715 35581 85727 35584
rect 85669 35575 85727 35581
rect 86221 35581 86233 35584
rect 86267 35581 86279 35615
rect 87874 35612 87880 35624
rect 87835 35584 87880 35612
rect 86221 35575 86279 35581
rect 85408 35544 85436 35575
rect 87874 35572 87880 35584
rect 87932 35572 87938 35624
rect 88058 35612 88064 35624
rect 88019 35584 88064 35612
rect 88058 35572 88064 35584
rect 88116 35612 88122 35624
rect 88521 35615 88579 35621
rect 88521 35612 88533 35615
rect 88116 35584 88533 35612
rect 88116 35572 88122 35584
rect 88521 35581 88533 35584
rect 88567 35581 88579 35615
rect 88521 35575 88579 35581
rect 86770 35544 86776 35556
rect 85408 35516 86776 35544
rect 86770 35504 86776 35516
rect 86828 35504 86834 35556
rect 79505 35479 79563 35485
rect 79505 35476 79517 35479
rect 77352 35448 79517 35476
rect 77352 35436 77358 35448
rect 79505 35445 79517 35448
rect 79551 35445 79563 35479
rect 79505 35439 79563 35445
rect 1104 35386 108008 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 81046 35386
rect 81098 35334 81110 35386
rect 81162 35334 81174 35386
rect 81226 35334 81238 35386
rect 81290 35334 108008 35386
rect 1104 35312 108008 35334
rect 3142 35232 3148 35284
rect 3200 35272 3206 35284
rect 4617 35275 4675 35281
rect 4617 35272 4629 35275
rect 3200 35244 4629 35272
rect 3200 35232 3206 35244
rect 4617 35241 4629 35244
rect 4663 35241 4675 35275
rect 4617 35235 4675 35241
rect 5445 35275 5503 35281
rect 5445 35241 5457 35275
rect 5491 35272 5503 35275
rect 5534 35272 5540 35284
rect 5491 35244 5540 35272
rect 5491 35241 5503 35244
rect 5445 35235 5503 35241
rect 5534 35232 5540 35244
rect 5592 35232 5598 35284
rect 6181 35275 6239 35281
rect 6181 35241 6193 35275
rect 6227 35241 6239 35275
rect 6181 35235 6239 35241
rect 16945 35275 17003 35281
rect 16945 35241 16957 35275
rect 16991 35272 17003 35275
rect 17310 35272 17316 35284
rect 16991 35244 17316 35272
rect 16991 35241 17003 35244
rect 16945 35235 17003 35241
rect 3510 35164 3516 35216
rect 3568 35204 3574 35216
rect 6196 35204 6224 35235
rect 17310 35232 17316 35244
rect 17368 35272 17374 35284
rect 17497 35275 17555 35281
rect 17497 35272 17509 35275
rect 17368 35244 17509 35272
rect 17368 35232 17374 35244
rect 17497 35241 17509 35244
rect 17543 35272 17555 35275
rect 18138 35272 18144 35284
rect 17543 35244 18144 35272
rect 17543 35241 17555 35244
rect 17497 35235 17555 35241
rect 18138 35232 18144 35244
rect 18196 35232 18202 35284
rect 21082 35272 21088 35284
rect 21043 35244 21088 35272
rect 21082 35232 21088 35244
rect 21140 35232 21146 35284
rect 21358 35272 21364 35284
rect 21319 35244 21364 35272
rect 21358 35232 21364 35244
rect 21416 35232 21422 35284
rect 32490 35272 32496 35284
rect 24136 35244 32496 35272
rect 24136 35204 24164 35244
rect 32490 35232 32496 35244
rect 32548 35232 32554 35284
rect 32674 35272 32680 35284
rect 32635 35244 32680 35272
rect 32674 35232 32680 35244
rect 32732 35232 32738 35284
rect 32950 35272 32956 35284
rect 32911 35244 32956 35272
rect 32950 35232 32956 35244
rect 33008 35232 33014 35284
rect 48777 35275 48835 35281
rect 48777 35272 48789 35275
rect 35084 35244 48789 35272
rect 26510 35204 26516 35216
rect 3568 35176 6224 35204
rect 14476 35176 24164 35204
rect 26471 35176 26516 35204
rect 3568 35164 3574 35176
rect 4801 35139 4859 35145
rect 4801 35105 4813 35139
rect 4847 35136 4859 35139
rect 4890 35136 4896 35148
rect 4847 35108 4896 35136
rect 4847 35105 4859 35108
rect 4801 35099 4859 35105
rect 4890 35096 4896 35108
rect 4948 35096 4954 35148
rect 5077 35139 5135 35145
rect 5077 35105 5089 35139
rect 5123 35136 5135 35139
rect 5534 35136 5540 35148
rect 5123 35108 5540 35136
rect 5123 35105 5135 35108
rect 5077 35099 5135 35105
rect 5534 35096 5540 35108
rect 5592 35096 5598 35148
rect 6086 35136 6092 35148
rect 6047 35108 6092 35136
rect 6086 35096 6092 35108
rect 6144 35096 6150 35148
rect 6641 35139 6699 35145
rect 6641 35105 6653 35139
rect 6687 35136 6699 35139
rect 6914 35136 6920 35148
rect 6687 35108 6920 35136
rect 6687 35105 6699 35108
rect 6641 35099 6699 35105
rect 6914 35096 6920 35108
rect 6972 35096 6978 35148
rect 13906 35096 13912 35148
rect 13964 35136 13970 35148
rect 14093 35139 14151 35145
rect 14093 35136 14105 35139
rect 13964 35108 14105 35136
rect 13964 35096 13970 35108
rect 14093 35105 14105 35108
rect 14139 35105 14151 35139
rect 14093 35099 14151 35105
rect 14476 35068 14504 35176
rect 26510 35164 26516 35176
rect 26568 35164 26574 35216
rect 26878 35164 26884 35216
rect 26936 35204 26942 35216
rect 35084 35204 35112 35244
rect 48777 35241 48789 35244
rect 48823 35241 48835 35275
rect 48777 35235 48835 35241
rect 55309 35275 55367 35281
rect 55309 35241 55321 35275
rect 55355 35272 55367 35275
rect 56594 35272 56600 35284
rect 55355 35244 56600 35272
rect 55355 35241 55367 35244
rect 55309 35235 55367 35241
rect 56594 35232 56600 35244
rect 56652 35232 56658 35284
rect 57241 35275 57299 35281
rect 57241 35241 57253 35275
rect 57287 35272 57299 35275
rect 58434 35272 58440 35284
rect 57287 35244 58440 35272
rect 57287 35241 57299 35244
rect 57241 35235 57299 35241
rect 58434 35232 58440 35244
rect 58492 35232 58498 35284
rect 79502 35272 79508 35284
rect 79463 35244 79508 35272
rect 79502 35232 79508 35244
rect 79560 35232 79566 35284
rect 87874 35232 87880 35284
rect 87932 35272 87938 35284
rect 88337 35275 88395 35281
rect 88337 35272 88349 35275
rect 87932 35244 88349 35272
rect 87932 35232 87938 35244
rect 88337 35241 88349 35244
rect 88383 35241 88395 35275
rect 88337 35235 88395 35241
rect 26936 35176 35112 35204
rect 26936 35164 26942 35176
rect 36262 35164 36268 35216
rect 36320 35204 36326 35216
rect 36357 35207 36415 35213
rect 36357 35204 36369 35207
rect 36320 35176 36369 35204
rect 36320 35164 36326 35176
rect 36357 35173 36369 35176
rect 36403 35204 36415 35207
rect 38381 35207 38439 35213
rect 36403 35176 36584 35204
rect 36403 35173 36415 35176
rect 36357 35167 36415 35173
rect 16945 35139 17003 35145
rect 16945 35105 16957 35139
rect 16991 35136 17003 35139
rect 17037 35139 17095 35145
rect 17037 35136 17049 35139
rect 16991 35108 17049 35136
rect 16991 35105 17003 35108
rect 16945 35099 17003 35105
rect 17037 35105 17049 35108
rect 17083 35105 17095 35139
rect 17037 35099 17095 35105
rect 20901 35139 20959 35145
rect 20901 35105 20913 35139
rect 20947 35136 20959 35139
rect 21358 35136 21364 35148
rect 20947 35108 21364 35136
rect 20947 35105 20959 35108
rect 20901 35099 20959 35105
rect 21358 35096 21364 35108
rect 21416 35096 21422 35148
rect 26602 35096 26608 35148
rect 26660 35136 26666 35148
rect 27154 35136 27160 35148
rect 26660 35108 27160 35136
rect 26660 35096 26666 35108
rect 27154 35096 27160 35108
rect 27212 35096 27218 35148
rect 27525 35139 27583 35145
rect 27525 35105 27537 35139
rect 27571 35136 27583 35139
rect 28074 35136 28080 35148
rect 27571 35108 28080 35136
rect 27571 35105 27583 35108
rect 27525 35099 27583 35105
rect 28074 35096 28080 35108
rect 28132 35136 28138 35148
rect 31662 35136 31668 35148
rect 28132 35108 31668 35136
rect 28132 35096 28138 35108
rect 31662 35096 31668 35108
rect 31720 35096 31726 35148
rect 32398 35096 32404 35148
rect 32456 35136 32462 35148
rect 36556 35145 36584 35176
rect 38381 35173 38393 35207
rect 38427 35204 38439 35207
rect 38470 35204 38476 35216
rect 38427 35176 38476 35204
rect 38427 35173 38439 35176
rect 38381 35167 38439 35173
rect 38470 35164 38476 35176
rect 38528 35164 38534 35216
rect 39574 35204 39580 35216
rect 39408 35176 39580 35204
rect 32493 35139 32551 35145
rect 32493 35136 32505 35139
rect 32456 35108 32505 35136
rect 32456 35096 32462 35108
rect 32493 35105 32505 35108
rect 32539 35105 32551 35139
rect 32493 35099 32551 35105
rect 36541 35139 36599 35145
rect 36541 35105 36553 35139
rect 36587 35105 36599 35139
rect 39408 35136 39436 35176
rect 39574 35164 39580 35176
rect 39632 35164 39638 35216
rect 39666 35164 39672 35216
rect 39724 35204 39730 35216
rect 40129 35207 40187 35213
rect 40129 35204 40141 35207
rect 39724 35176 40141 35204
rect 39724 35164 39730 35176
rect 40129 35173 40141 35176
rect 40175 35204 40187 35207
rect 42610 35204 42616 35216
rect 40175 35176 42616 35204
rect 40175 35173 40187 35176
rect 40129 35167 40187 35173
rect 42610 35164 42616 35176
rect 42668 35164 42674 35216
rect 43806 35164 43812 35216
rect 43864 35204 43870 35216
rect 44545 35207 44603 35213
rect 44545 35204 44557 35207
rect 43864 35176 44557 35204
rect 43864 35164 43870 35176
rect 44545 35173 44557 35176
rect 44591 35173 44603 35207
rect 44545 35167 44603 35173
rect 44821 35207 44879 35213
rect 44821 35173 44833 35207
rect 44867 35204 44879 35207
rect 45554 35204 45560 35216
rect 44867 35176 45560 35204
rect 44867 35173 44879 35176
rect 44821 35167 44879 35173
rect 36541 35099 36599 35105
rect 36648 35108 39436 35136
rect 5092 35040 14504 35068
rect 5092 35012 5120 35040
rect 16482 35028 16488 35080
rect 16540 35068 16546 35080
rect 26694 35068 26700 35080
rect 16540 35040 26700 35068
rect 16540 35028 16546 35040
rect 26694 35028 26700 35040
rect 26752 35028 26758 35080
rect 5074 34960 5080 35012
rect 5132 34960 5138 35012
rect 26878 35000 26884 35012
rect 13740 34972 26884 35000
rect 3786 34892 3792 34944
rect 3844 34932 3850 34944
rect 13740 34932 13768 34972
rect 26878 34960 26884 34972
rect 26936 34960 26942 35012
rect 27172 35000 27200 35096
rect 27246 35028 27252 35080
rect 27304 35068 27310 35080
rect 27430 35068 27436 35080
rect 27304 35040 27349 35068
rect 27391 35040 27436 35068
rect 27304 35028 27310 35040
rect 27430 35028 27436 35040
rect 27488 35028 27494 35080
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35068 27951 35071
rect 36648 35068 36676 35108
rect 42426 35096 42432 35148
rect 42484 35136 42490 35148
rect 42978 35136 42984 35148
rect 42484 35108 42984 35136
rect 42484 35096 42490 35108
rect 42978 35096 42984 35108
rect 43036 35136 43042 35148
rect 43349 35139 43407 35145
rect 43349 35136 43361 35139
rect 43036 35108 43361 35136
rect 43036 35096 43042 35108
rect 43349 35105 43361 35108
rect 43395 35136 43407 35139
rect 43717 35139 43775 35145
rect 43717 35136 43729 35139
rect 43395 35108 43729 35136
rect 43395 35105 43407 35108
rect 43349 35099 43407 35105
rect 43717 35105 43729 35108
rect 43763 35105 43775 35139
rect 43717 35099 43775 35105
rect 44453 35139 44511 35145
rect 44453 35105 44465 35139
rect 44499 35136 44511 35139
rect 44836 35136 44864 35167
rect 45554 35164 45560 35176
rect 45612 35164 45618 35216
rect 55214 35204 55220 35216
rect 51736 35176 55220 35204
rect 44499 35108 44864 35136
rect 44499 35105 44511 35108
rect 44453 35099 44511 35105
rect 38470 35068 38476 35080
rect 27939 35040 36676 35068
rect 38431 35040 38476 35068
rect 27939 35037 27951 35040
rect 27893 35031 27951 35037
rect 27908 35000 27936 35031
rect 38470 35028 38476 35040
rect 38528 35028 38534 35080
rect 38746 35068 38752 35080
rect 38707 35040 38752 35068
rect 38746 35028 38752 35040
rect 38804 35028 38810 35080
rect 43165 35071 43223 35077
rect 43165 35037 43177 35071
rect 43211 35068 43223 35071
rect 51736 35068 51764 35176
rect 55214 35164 55220 35176
rect 55272 35164 55278 35216
rect 64782 35164 64788 35216
rect 64840 35204 64846 35216
rect 64840 35176 71912 35204
rect 64840 35164 64846 35176
rect 52546 35096 52552 35148
rect 52604 35136 52610 35148
rect 55493 35139 55551 35145
rect 55493 35136 55505 35139
rect 52604 35108 55505 35136
rect 52604 35096 52610 35108
rect 55493 35105 55505 35108
rect 55539 35136 55551 35139
rect 55677 35139 55735 35145
rect 55677 35136 55689 35139
rect 55539 35108 55689 35136
rect 55539 35105 55551 35108
rect 55493 35099 55551 35105
rect 55677 35105 55689 35108
rect 55723 35136 55735 35139
rect 56229 35139 56287 35145
rect 56229 35136 56241 35139
rect 55723 35108 56241 35136
rect 55723 35105 55735 35108
rect 55677 35099 55735 35105
rect 56229 35105 56241 35108
rect 56275 35136 56287 35139
rect 56781 35139 56839 35145
rect 56781 35136 56793 35139
rect 56275 35108 56793 35136
rect 56275 35105 56287 35108
rect 56229 35099 56287 35105
rect 56781 35105 56793 35108
rect 56827 35105 56839 35139
rect 56962 35136 56968 35148
rect 56875 35108 56968 35136
rect 56781 35099 56839 35105
rect 56962 35096 56968 35108
rect 57020 35136 57026 35148
rect 57609 35139 57667 35145
rect 57609 35136 57621 35139
rect 57020 35108 57621 35136
rect 57020 35096 57026 35108
rect 57609 35105 57621 35108
rect 57655 35136 57667 35139
rect 63218 35136 63224 35148
rect 57655 35108 63224 35136
rect 57655 35105 57667 35108
rect 57609 35099 57667 35105
rect 63218 35096 63224 35108
rect 63276 35096 63282 35148
rect 67910 35136 67916 35148
rect 67823 35108 67916 35136
rect 67910 35096 67916 35108
rect 67968 35136 67974 35148
rect 68554 35136 68560 35148
rect 67968 35108 68560 35136
rect 67968 35096 67974 35108
rect 68554 35096 68560 35108
rect 68612 35096 68618 35148
rect 71884 35136 71912 35176
rect 72053 35139 72111 35145
rect 72053 35136 72065 35139
rect 71884 35108 72065 35136
rect 72053 35105 72065 35108
rect 72099 35136 72111 35139
rect 72329 35139 72387 35145
rect 72329 35136 72341 35139
rect 72099 35108 72341 35136
rect 72099 35105 72111 35108
rect 72053 35099 72111 35105
rect 72329 35105 72341 35108
rect 72375 35136 72387 35139
rect 72878 35136 72884 35148
rect 72375 35108 72884 35136
rect 72375 35105 72387 35108
rect 72329 35099 72387 35105
rect 72878 35096 72884 35108
rect 72936 35096 72942 35148
rect 74994 35136 75000 35148
rect 74955 35108 75000 35136
rect 74994 35096 75000 35108
rect 75052 35096 75058 35148
rect 75181 35139 75239 35145
rect 75181 35105 75193 35139
rect 75227 35136 75239 35139
rect 77018 35136 77024 35148
rect 75227 35108 75776 35136
rect 76979 35108 77024 35136
rect 75227 35105 75239 35108
rect 75181 35099 75239 35105
rect 43211 35040 51764 35068
rect 55309 35071 55367 35077
rect 43211 35037 43223 35040
rect 43165 35031 43223 35037
rect 55309 35037 55321 35071
rect 55355 35068 55367 35071
rect 55861 35071 55919 35077
rect 55861 35068 55873 35071
rect 55355 35040 55873 35068
rect 55355 35037 55367 35040
rect 55309 35031 55367 35037
rect 55861 35037 55873 35040
rect 55907 35068 55919 35071
rect 56045 35071 56103 35077
rect 56045 35068 56057 35071
rect 55907 35040 56057 35068
rect 55907 35037 55919 35040
rect 55861 35031 55919 35037
rect 56045 35037 56057 35040
rect 56091 35037 56103 35071
rect 75546 35068 75552 35080
rect 75507 35040 75552 35068
rect 56045 35031 56103 35037
rect 75546 35028 75552 35040
rect 75604 35028 75610 35080
rect 28074 35000 28080 35012
rect 27172 34972 27936 35000
rect 28035 34972 28080 35000
rect 28074 34960 28080 34972
rect 28132 34960 28138 35012
rect 36725 35003 36783 35009
rect 36725 34969 36737 35003
rect 36771 35000 36783 35003
rect 37182 35000 37188 35012
rect 36771 34972 37188 35000
rect 36771 34969 36783 34972
rect 36725 34963 36783 34969
rect 37182 34960 37188 34972
rect 37240 35000 37246 35012
rect 37642 35000 37648 35012
rect 37240 34972 37648 35000
rect 37240 34960 37246 34972
rect 37642 34960 37648 34972
rect 37700 34960 37706 35012
rect 39574 34960 39580 35012
rect 39632 35000 39638 35012
rect 72142 35000 72148 35012
rect 39632 34972 72148 35000
rect 39632 34960 39638 34972
rect 72142 34960 72148 34972
rect 72200 35000 72206 35012
rect 75178 35000 75184 35012
rect 72200 34972 75184 35000
rect 72200 34960 72206 34972
rect 75178 34960 75184 34972
rect 75236 34960 75242 35012
rect 13906 34932 13912 34944
rect 3844 34904 13768 34932
rect 13867 34904 13912 34932
rect 3844 34892 3850 34904
rect 13906 34892 13912 34904
rect 13964 34892 13970 34944
rect 14182 34932 14188 34944
rect 14143 34904 14188 34932
rect 14182 34892 14188 34904
rect 14240 34892 14246 34944
rect 17218 34932 17224 34944
rect 17179 34904 17224 34932
rect 17218 34892 17224 34904
rect 17276 34892 17282 34944
rect 20530 34892 20536 34944
rect 20588 34932 20594 34944
rect 21910 34932 21916 34944
rect 20588 34904 21916 34932
rect 20588 34892 20594 34904
rect 21910 34892 21916 34904
rect 21968 34892 21974 34944
rect 32490 34892 32496 34944
rect 32548 34932 32554 34944
rect 37366 34932 37372 34944
rect 32548 34904 37372 34932
rect 32548 34892 32554 34904
rect 37366 34892 37372 34904
rect 37424 34892 37430 34944
rect 37458 34892 37464 34944
rect 37516 34932 37522 34944
rect 43165 34935 43223 34941
rect 43165 34932 43177 34935
rect 37516 34904 43177 34932
rect 37516 34892 37522 34904
rect 43165 34901 43177 34904
rect 43211 34901 43223 34935
rect 43165 34895 43223 34901
rect 43254 34892 43260 34944
rect 43312 34932 43318 34944
rect 43533 34935 43591 34941
rect 43533 34932 43545 34935
rect 43312 34904 43545 34932
rect 43312 34892 43318 34904
rect 43533 34901 43545 34904
rect 43579 34932 43591 34935
rect 43806 34932 43812 34944
rect 43579 34904 43812 34932
rect 43579 34901 43591 34904
rect 43533 34895 43591 34901
rect 43806 34892 43812 34904
rect 43864 34892 43870 34944
rect 48777 34935 48835 34941
rect 48777 34901 48789 34935
rect 48823 34932 48835 34935
rect 55309 34935 55367 34941
rect 55309 34932 55321 34935
rect 48823 34904 55321 34932
rect 48823 34901 48835 34904
rect 48777 34895 48835 34901
rect 55309 34901 55321 34904
rect 55355 34901 55367 34935
rect 55309 34895 55367 34901
rect 67726 34892 67732 34944
rect 67784 34932 67790 34944
rect 68002 34932 68008 34944
rect 67784 34904 68008 34932
rect 67784 34892 67790 34904
rect 68002 34892 68008 34904
rect 68060 34892 68066 34944
rect 75748 34941 75776 35108
rect 77018 35096 77024 35108
rect 77076 35096 77082 35148
rect 77202 35096 77208 35148
rect 77260 35136 77266 35148
rect 79321 35139 79379 35145
rect 79321 35136 79333 35139
rect 77260 35108 79333 35136
rect 77260 35096 77266 35108
rect 79321 35105 79333 35108
rect 79367 35105 79379 35139
rect 79321 35099 79379 35105
rect 87322 35096 87328 35148
rect 87380 35136 87386 35148
rect 88245 35139 88303 35145
rect 88245 35136 88257 35139
rect 87380 35108 88257 35136
rect 87380 35096 87386 35108
rect 88245 35105 88257 35108
rect 88291 35105 88303 35139
rect 88245 35099 88303 35105
rect 75733 34935 75791 34941
rect 75733 34901 75745 34935
rect 75779 34932 75791 34935
rect 75822 34932 75828 34944
rect 75779 34904 75828 34932
rect 75779 34901 75791 34904
rect 75733 34895 75791 34901
rect 75822 34892 75828 34904
rect 75880 34892 75886 34944
rect 76834 34892 76840 34944
rect 76892 34932 76898 34944
rect 77113 34935 77171 34941
rect 77113 34932 77125 34935
rect 76892 34904 77125 34932
rect 76892 34892 76898 34904
rect 77113 34901 77125 34904
rect 77159 34901 77171 34935
rect 77113 34895 77171 34901
rect 1104 34842 108008 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 65686 34842
rect 65738 34790 65750 34842
rect 65802 34790 65814 34842
rect 65866 34790 65878 34842
rect 65930 34790 96406 34842
rect 96458 34790 96470 34842
rect 96522 34790 96534 34842
rect 96586 34790 96598 34842
rect 96650 34790 108008 34842
rect 1104 34768 108008 34790
rect 5537 34731 5595 34737
rect 5537 34697 5549 34731
rect 5583 34728 5595 34731
rect 19334 34728 19340 34740
rect 5583 34700 19340 34728
rect 5583 34697 5595 34700
rect 5537 34691 5595 34697
rect 4890 34524 4896 34536
rect 4851 34496 4896 34524
rect 4890 34484 4896 34496
rect 4948 34484 4954 34536
rect 5169 34527 5227 34533
rect 5169 34493 5181 34527
rect 5215 34524 5227 34527
rect 5552 34524 5580 34691
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 21818 34728 21824 34740
rect 21008 34700 21824 34728
rect 7282 34660 7288 34672
rect 7243 34632 7288 34660
rect 7282 34620 7288 34632
rect 7340 34620 7346 34672
rect 14182 34620 14188 34672
rect 14240 34660 14246 34672
rect 15105 34663 15163 34669
rect 15105 34660 15117 34663
rect 14240 34632 15117 34660
rect 14240 34620 14246 34632
rect 15105 34629 15117 34632
rect 15151 34660 15163 34663
rect 15746 34660 15752 34672
rect 15151 34632 15752 34660
rect 15151 34629 15163 34632
rect 15105 34623 15163 34629
rect 15746 34620 15752 34632
rect 15804 34660 15810 34672
rect 16666 34660 16672 34672
rect 15804 34632 16672 34660
rect 15804 34620 15810 34632
rect 16666 34620 16672 34632
rect 16724 34620 16730 34672
rect 7098 34524 7104 34536
rect 5215 34496 5580 34524
rect 7059 34496 7104 34524
rect 5215 34493 5227 34496
rect 5169 34487 5227 34493
rect 7098 34484 7104 34496
rect 7156 34484 7162 34536
rect 7300 34524 7328 34620
rect 21008 34601 21036 34700
rect 21818 34688 21824 34700
rect 21876 34688 21882 34740
rect 22002 34688 22008 34740
rect 22060 34728 22066 34740
rect 22097 34731 22155 34737
rect 22097 34728 22109 34731
rect 22060 34700 22109 34728
rect 22060 34688 22066 34700
rect 22097 34697 22109 34700
rect 22143 34697 22155 34731
rect 27341 34731 27399 34737
rect 22097 34691 22155 34697
rect 25792 34700 27292 34728
rect 21082 34620 21088 34672
rect 21140 34660 21146 34672
rect 21913 34663 21971 34669
rect 21913 34660 21925 34663
rect 21140 34632 21925 34660
rect 21140 34620 21146 34632
rect 21913 34629 21925 34632
rect 21959 34629 21971 34663
rect 21913 34623 21971 34629
rect 20257 34595 20315 34601
rect 20257 34592 20269 34595
rect 9876 34564 20269 34592
rect 8205 34527 8263 34533
rect 8205 34524 8217 34527
rect 7300 34496 8217 34524
rect 8205 34493 8217 34496
rect 8251 34493 8263 34527
rect 8205 34487 8263 34493
rect 8757 34527 8815 34533
rect 8757 34493 8769 34527
rect 8803 34524 8815 34527
rect 9876 34524 9904 34564
rect 20257 34561 20269 34564
rect 20303 34561 20315 34595
rect 20257 34555 20315 34561
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34561 21051 34595
rect 21637 34595 21695 34601
rect 21637 34592 21649 34595
rect 20993 34555 21051 34561
rect 21468 34564 21649 34592
rect 8803 34496 9904 34524
rect 13081 34527 13139 34533
rect 8803 34493 8815 34496
rect 8757 34487 8815 34493
rect 13081 34493 13093 34527
rect 13127 34524 13139 34527
rect 13814 34524 13820 34536
rect 13127 34496 13820 34524
rect 13127 34493 13139 34496
rect 13081 34487 13139 34493
rect 13814 34484 13820 34496
rect 13872 34484 13878 34536
rect 15746 34524 15752 34536
rect 15707 34496 15752 34524
rect 15746 34484 15752 34496
rect 15804 34484 15810 34536
rect 15838 34484 15844 34536
rect 15896 34524 15902 34536
rect 16025 34527 16083 34533
rect 16025 34524 16037 34527
rect 15896 34496 16037 34524
rect 15896 34484 15902 34496
rect 16025 34493 16037 34496
rect 16071 34524 16083 34527
rect 16114 34524 16120 34536
rect 16071 34496 16120 34524
rect 16071 34493 16083 34496
rect 16025 34487 16083 34493
rect 16114 34484 16120 34496
rect 16172 34484 16178 34536
rect 16206 34484 16212 34536
rect 16264 34524 16270 34536
rect 16264 34496 16309 34524
rect 16264 34484 16270 34496
rect 16574 34484 16580 34536
rect 16632 34524 16638 34536
rect 19886 34524 19892 34536
rect 16632 34496 19892 34524
rect 16632 34484 16638 34496
rect 19886 34484 19892 34496
rect 19944 34484 19950 34536
rect 20530 34484 20536 34536
rect 20588 34524 20594 34536
rect 20901 34527 20959 34533
rect 20901 34524 20913 34527
rect 20588 34496 20913 34524
rect 20588 34484 20594 34496
rect 20901 34493 20913 34496
rect 20947 34493 20959 34527
rect 20901 34487 20959 34493
rect 21082 34484 21088 34536
rect 21140 34524 21146 34536
rect 21468 34533 21496 34564
rect 21637 34561 21649 34564
rect 21683 34592 21695 34595
rect 25590 34592 25596 34604
rect 21683 34564 25596 34592
rect 21683 34561 21695 34564
rect 21637 34555 21695 34561
rect 25590 34552 25596 34564
rect 25648 34552 25654 34604
rect 25792 34592 25820 34700
rect 27264 34660 27292 34700
rect 27341 34697 27353 34731
rect 27387 34728 27399 34731
rect 27430 34728 27436 34740
rect 27387 34700 27436 34728
rect 27387 34697 27399 34700
rect 27341 34691 27399 34697
rect 27430 34688 27436 34700
rect 27488 34688 27494 34740
rect 27614 34688 27620 34740
rect 27672 34728 27678 34740
rect 37001 34731 37059 34737
rect 37001 34728 37013 34731
rect 27672 34700 37013 34728
rect 27672 34688 27678 34700
rect 37001 34697 37013 34700
rect 37047 34697 37059 34731
rect 37001 34691 37059 34697
rect 37274 34688 37280 34740
rect 37332 34728 37338 34740
rect 38838 34728 38844 34740
rect 37332 34700 38844 34728
rect 37332 34688 37338 34700
rect 38838 34688 38844 34700
rect 38896 34688 38902 34740
rect 39666 34728 39672 34740
rect 39627 34700 39672 34728
rect 39666 34688 39672 34700
rect 39724 34688 39730 34740
rect 40313 34731 40371 34737
rect 40313 34697 40325 34731
rect 40359 34728 40371 34731
rect 49142 34728 49148 34740
rect 40359 34700 49148 34728
rect 40359 34697 40371 34700
rect 40313 34691 40371 34697
rect 49142 34688 49148 34700
rect 49200 34688 49206 34740
rect 51442 34728 51448 34740
rect 51403 34700 51448 34728
rect 51442 34688 51448 34700
rect 51500 34688 51506 34740
rect 53285 34731 53343 34737
rect 53285 34697 53297 34731
rect 53331 34728 53343 34731
rect 56962 34728 56968 34740
rect 53331 34700 56968 34728
rect 53331 34697 53343 34700
rect 53285 34691 53343 34697
rect 27706 34660 27712 34672
rect 27264 34632 27712 34660
rect 27706 34620 27712 34632
rect 27764 34620 27770 34672
rect 41598 34660 41604 34672
rect 32324 34632 41604 34660
rect 25792 34564 25912 34592
rect 21269 34527 21327 34533
rect 21269 34524 21281 34527
rect 21140 34496 21281 34524
rect 21140 34484 21146 34496
rect 21269 34493 21281 34496
rect 21315 34493 21327 34527
rect 21269 34487 21327 34493
rect 21453 34527 21511 34533
rect 21453 34493 21465 34527
rect 21499 34493 21511 34527
rect 21453 34487 21511 34493
rect 25682 34484 25688 34536
rect 25740 34524 25746 34536
rect 25777 34527 25835 34533
rect 25777 34524 25789 34527
rect 25740 34496 25789 34524
rect 25740 34484 25746 34496
rect 25777 34493 25789 34496
rect 25823 34493 25835 34527
rect 25884 34524 25912 34564
rect 25958 34552 25964 34604
rect 26016 34592 26022 34604
rect 32324 34592 32352 34632
rect 41598 34620 41604 34632
rect 41656 34620 41662 34672
rect 44266 34660 44272 34672
rect 44227 34632 44272 34660
rect 44266 34620 44272 34632
rect 44324 34620 44330 34672
rect 44358 34620 44364 34672
rect 44416 34660 44422 34672
rect 44637 34663 44695 34669
rect 44637 34660 44649 34663
rect 44416 34632 44649 34660
rect 44416 34620 44422 34632
rect 44637 34629 44649 34632
rect 44683 34660 44695 34663
rect 44821 34663 44879 34669
rect 44821 34660 44833 34663
rect 44683 34632 44833 34660
rect 44683 34629 44695 34632
rect 44637 34623 44695 34629
rect 44821 34629 44833 34632
rect 44867 34660 44879 34663
rect 52546 34660 52552 34672
rect 44867 34632 52552 34660
rect 44867 34629 44879 34632
rect 44821 34623 44879 34629
rect 52546 34620 52552 34632
rect 52604 34620 52610 34672
rect 26016 34564 32352 34592
rect 26016 34552 26022 34564
rect 32398 34552 32404 34604
rect 32456 34592 32462 34604
rect 32950 34592 32956 34604
rect 32456 34564 32956 34592
rect 32456 34552 32462 34564
rect 32950 34552 32956 34564
rect 33008 34552 33014 34604
rect 36633 34595 36691 34601
rect 36633 34561 36645 34595
rect 36679 34592 36691 34595
rect 38286 34592 38292 34604
rect 36679 34564 38292 34592
rect 36679 34561 36691 34564
rect 36633 34555 36691 34561
rect 26053 34527 26111 34533
rect 26053 34524 26065 34527
rect 25884 34496 26065 34524
rect 25777 34487 25835 34493
rect 26053 34493 26065 34496
rect 26099 34493 26111 34527
rect 26053 34487 26111 34493
rect 26142 34484 26148 34536
rect 26200 34524 26206 34536
rect 37185 34527 37243 34533
rect 26200 34496 27752 34524
rect 26200 34484 26206 34496
rect 5258 34416 5264 34468
rect 5316 34456 5322 34468
rect 5353 34459 5411 34465
rect 5353 34456 5365 34459
rect 5316 34428 5365 34456
rect 5316 34416 5322 34428
rect 5353 34425 5365 34428
rect 5399 34425 5411 34459
rect 5353 34419 5411 34425
rect 8941 34459 8999 34465
rect 8941 34425 8953 34459
rect 8987 34456 8999 34459
rect 9030 34456 9036 34468
rect 8987 34428 9036 34456
rect 8987 34425 8999 34428
rect 8941 34419 8999 34425
rect 9030 34416 9036 34428
rect 9088 34416 9094 34468
rect 15197 34459 15255 34465
rect 12544 34428 13308 34456
rect 6362 34348 6368 34400
rect 6420 34388 6426 34400
rect 12544 34388 12572 34428
rect 13170 34388 13176 34400
rect 6420 34360 12572 34388
rect 13131 34360 13176 34388
rect 6420 34348 6426 34360
rect 13170 34348 13176 34360
rect 13228 34348 13234 34400
rect 13280 34388 13308 34428
rect 15197 34425 15209 34459
rect 15243 34456 15255 34459
rect 15562 34456 15568 34468
rect 15243 34428 15568 34456
rect 15243 34425 15255 34428
rect 15197 34419 15255 34425
rect 15562 34416 15568 34428
rect 15620 34416 15626 34468
rect 27724 34456 27752 34496
rect 37185 34493 37197 34527
rect 37231 34524 37243 34527
rect 37274 34524 37280 34536
rect 37231 34496 37280 34524
rect 37231 34493 37243 34496
rect 37185 34487 37243 34493
rect 37274 34484 37280 34496
rect 37332 34484 37338 34536
rect 37366 34484 37372 34536
rect 37424 34524 37430 34536
rect 37752 34533 37780 34564
rect 38286 34552 38292 34564
rect 38344 34592 38350 34604
rect 40313 34595 40371 34601
rect 40313 34592 40325 34595
rect 38344 34564 40325 34592
rect 38344 34552 38350 34564
rect 40313 34561 40325 34564
rect 40359 34561 40371 34595
rect 40313 34555 40371 34561
rect 46934 34552 46940 34604
rect 46992 34592 46998 34604
rect 51905 34595 51963 34601
rect 51905 34592 51917 34595
rect 46992 34564 51917 34592
rect 46992 34552 46998 34564
rect 51905 34561 51917 34564
rect 51951 34561 51963 34595
rect 51905 34555 51963 34561
rect 52641 34595 52699 34601
rect 52641 34561 52653 34595
rect 52687 34592 52699 34595
rect 53300 34592 53328 34691
rect 56962 34688 56968 34700
rect 57020 34688 57026 34740
rect 57054 34688 57060 34740
rect 57112 34728 57118 34740
rect 62669 34731 62727 34737
rect 62669 34728 62681 34731
rect 57112 34700 62681 34728
rect 57112 34688 57118 34700
rect 60829 34663 60887 34669
rect 60829 34660 60841 34663
rect 60384 34632 60841 34660
rect 59446 34592 59452 34604
rect 52687 34564 53328 34592
rect 59407 34564 59452 34592
rect 52687 34561 52699 34564
rect 52641 34555 52699 34561
rect 59446 34552 59452 34564
rect 59504 34552 59510 34604
rect 59722 34592 59728 34604
rect 59683 34564 59728 34592
rect 59722 34552 59728 34564
rect 59780 34552 59786 34604
rect 59906 34552 59912 34604
rect 59964 34592 59970 34604
rect 60384 34592 60412 34632
rect 60829 34629 60841 34632
rect 60875 34629 60887 34663
rect 60829 34623 60887 34629
rect 60918 34620 60924 34672
rect 60976 34660 60982 34672
rect 61197 34663 61255 34669
rect 61197 34660 61209 34663
rect 60976 34632 61209 34660
rect 60976 34620 60982 34632
rect 61197 34629 61209 34632
rect 61243 34629 61255 34663
rect 61197 34623 61255 34629
rect 59964 34564 60412 34592
rect 62500 34592 62528 34700
rect 62669 34697 62681 34700
rect 62715 34697 62727 34731
rect 62669 34691 62727 34697
rect 63034 34688 63040 34740
rect 63092 34728 63098 34740
rect 64417 34731 64475 34737
rect 64417 34728 64429 34731
rect 63092 34700 64429 34728
rect 63092 34688 63098 34700
rect 64417 34697 64429 34700
rect 64463 34728 64475 34731
rect 67729 34731 67787 34737
rect 67729 34728 67741 34731
rect 64463 34700 67741 34728
rect 64463 34697 64475 34700
rect 64417 34691 64475 34697
rect 67729 34697 67741 34700
rect 67775 34697 67787 34731
rect 68094 34728 68100 34740
rect 68055 34700 68100 34728
rect 67729 34691 67787 34697
rect 68094 34688 68100 34700
rect 68152 34728 68158 34740
rect 68922 34728 68928 34740
rect 68152 34700 68928 34728
rect 68152 34688 68158 34700
rect 68922 34688 68928 34700
rect 68980 34688 68986 34740
rect 75730 34688 75736 34740
rect 75788 34728 75794 34740
rect 76653 34731 76711 34737
rect 76653 34728 76665 34731
rect 75788 34700 76665 34728
rect 75788 34688 75794 34700
rect 76653 34697 76665 34700
rect 76699 34728 76711 34731
rect 77018 34728 77024 34740
rect 76699 34700 77024 34728
rect 76699 34697 76711 34700
rect 76653 34691 76711 34697
rect 77018 34688 77024 34700
rect 77076 34688 77082 34740
rect 77113 34731 77171 34737
rect 77113 34697 77125 34731
rect 77159 34697 77171 34731
rect 77113 34691 77171 34697
rect 62574 34620 62580 34672
rect 62632 34660 62638 34672
rect 64049 34663 64107 34669
rect 64049 34660 64061 34663
rect 62632 34632 64061 34660
rect 62632 34620 62638 34632
rect 64049 34629 64061 34632
rect 64095 34629 64107 34663
rect 64049 34623 64107 34629
rect 64693 34663 64751 34669
rect 64693 34629 64705 34663
rect 64739 34660 64751 34663
rect 68278 34660 68284 34672
rect 64739 34632 68284 34660
rect 64739 34629 64751 34632
rect 64693 34623 64751 34629
rect 62500 34564 63356 34592
rect 59964 34552 59970 34564
rect 37737 34527 37795 34533
rect 37424 34496 37469 34524
rect 37424 34484 37430 34496
rect 37737 34493 37749 34527
rect 37783 34493 37795 34527
rect 37737 34487 37795 34493
rect 37921 34527 37979 34533
rect 37921 34493 37933 34527
rect 37967 34524 37979 34527
rect 38102 34524 38108 34536
rect 37967 34496 38108 34524
rect 37967 34493 37979 34496
rect 37921 34487 37979 34493
rect 38102 34484 38108 34496
rect 38160 34484 38166 34536
rect 38194 34484 38200 34536
rect 38252 34524 38258 34536
rect 39206 34524 39212 34536
rect 38252 34496 39212 34524
rect 38252 34484 38258 34496
rect 39206 34484 39212 34496
rect 39264 34484 39270 34536
rect 39301 34527 39359 34533
rect 39301 34493 39313 34527
rect 39347 34524 39359 34527
rect 39666 34524 39672 34536
rect 39347 34496 39672 34524
rect 39347 34493 39359 34496
rect 39301 34487 39359 34493
rect 39666 34484 39672 34496
rect 39724 34484 39730 34536
rect 39758 34484 39764 34536
rect 39816 34524 39822 34536
rect 41506 34524 41512 34536
rect 39816 34496 41512 34524
rect 39816 34484 39822 34496
rect 41506 34484 41512 34496
rect 41564 34484 41570 34536
rect 42886 34524 42892 34536
rect 42847 34496 42892 34524
rect 42886 34484 42892 34496
rect 42944 34524 42950 34536
rect 43073 34527 43131 34533
rect 43073 34524 43085 34527
rect 42944 34496 43085 34524
rect 42944 34484 42950 34496
rect 43073 34493 43085 34496
rect 43119 34493 43131 34527
rect 43254 34524 43260 34536
rect 43215 34496 43260 34524
rect 43073 34487 43131 34493
rect 43254 34484 43260 34496
rect 43312 34484 43318 34536
rect 43714 34524 43720 34536
rect 43675 34496 43720 34524
rect 43714 34484 43720 34496
rect 43772 34484 43778 34536
rect 43806 34484 43812 34536
rect 43864 34524 43870 34536
rect 43990 34524 43996 34536
rect 43864 34496 43996 34524
rect 43864 34484 43870 34496
rect 43990 34484 43996 34496
rect 44048 34484 44054 34536
rect 49694 34484 49700 34536
rect 49752 34524 49758 34536
rect 51721 34527 51779 34533
rect 51721 34524 51733 34527
rect 49752 34496 51733 34524
rect 49752 34484 49758 34496
rect 51721 34493 51733 34496
rect 51767 34524 51779 34527
rect 52549 34527 52607 34533
rect 52549 34524 52561 34527
rect 51767 34496 52561 34524
rect 51767 34493 51779 34496
rect 51721 34487 51779 34493
rect 52549 34493 52561 34496
rect 52595 34493 52607 34527
rect 52549 34487 52607 34493
rect 52822 34484 52828 34536
rect 52880 34524 52886 34536
rect 52917 34527 52975 34533
rect 52917 34524 52929 34527
rect 52880 34496 52929 34524
rect 52880 34484 52886 34496
rect 52917 34493 52929 34496
rect 52963 34493 52975 34527
rect 52917 34487 52975 34493
rect 53101 34527 53159 34533
rect 53101 34493 53113 34527
rect 53147 34524 53159 34527
rect 57698 34524 57704 34536
rect 53147 34496 57704 34524
rect 53147 34493 53159 34496
rect 53101 34487 53159 34493
rect 57698 34484 57704 34496
rect 57756 34484 57762 34536
rect 62390 34484 62396 34536
rect 62448 34524 62454 34536
rect 62945 34527 63003 34533
rect 62945 34524 62957 34527
rect 62448 34496 62957 34524
rect 62448 34484 62454 34496
rect 62945 34493 62957 34496
rect 62991 34493 63003 34527
rect 62945 34487 63003 34493
rect 63034 34484 63040 34536
rect 63092 34524 63098 34536
rect 63129 34527 63187 34533
rect 63129 34524 63141 34527
rect 63092 34496 63141 34524
rect 63092 34484 63098 34496
rect 63129 34493 63141 34496
rect 63175 34493 63187 34527
rect 63328 34524 63356 34564
rect 63589 34527 63647 34533
rect 63589 34524 63601 34527
rect 63328 34496 63601 34524
rect 63129 34487 63187 34493
rect 63589 34493 63601 34496
rect 63635 34493 63647 34527
rect 63589 34487 63647 34493
rect 63681 34527 63739 34533
rect 63681 34493 63693 34527
rect 63727 34524 63739 34527
rect 64708 34524 64736 34623
rect 68278 34620 68284 34632
rect 68336 34660 68342 34672
rect 68646 34660 68652 34672
rect 68336 34632 68652 34660
rect 68336 34620 68342 34632
rect 68646 34620 68652 34632
rect 68704 34620 68710 34672
rect 74994 34620 75000 34672
rect 75052 34660 75058 34672
rect 77128 34660 77156 34691
rect 75052 34632 77156 34660
rect 75052 34620 75058 34632
rect 67913 34595 67971 34601
rect 67913 34561 67925 34595
rect 67959 34592 67971 34595
rect 68094 34592 68100 34604
rect 67959 34564 68100 34592
rect 67959 34561 67971 34564
rect 67913 34555 67971 34561
rect 68094 34552 68100 34564
rect 68152 34592 68158 34604
rect 68557 34595 68615 34601
rect 68557 34592 68569 34595
rect 68152 34564 68569 34592
rect 68152 34552 68158 34564
rect 68557 34561 68569 34564
rect 68603 34561 68615 34595
rect 68557 34555 68615 34561
rect 63727 34496 64736 34524
rect 65613 34527 65671 34533
rect 63727 34493 63739 34496
rect 63681 34487 63739 34493
rect 65613 34493 65625 34527
rect 65659 34524 65671 34527
rect 65978 34524 65984 34536
rect 65659 34496 65984 34524
rect 65659 34493 65671 34496
rect 65613 34487 65671 34493
rect 65978 34484 65984 34496
rect 66036 34484 66042 34536
rect 67729 34527 67787 34533
rect 67729 34493 67741 34527
rect 67775 34524 67787 34527
rect 68741 34527 68799 34533
rect 68741 34524 68753 34527
rect 67775 34496 68753 34524
rect 67775 34493 67787 34496
rect 67729 34487 67787 34493
rect 68741 34493 68753 34496
rect 68787 34493 68799 34527
rect 68741 34487 68799 34493
rect 59538 34456 59544 34468
rect 15672 34428 25912 34456
rect 15672 34388 15700 34428
rect 13280 34360 15700 34388
rect 16666 34348 16672 34400
rect 16724 34388 16730 34400
rect 25774 34388 25780 34400
rect 16724 34360 25780 34388
rect 16724 34348 16730 34360
rect 25774 34348 25780 34360
rect 25832 34348 25838 34400
rect 25884 34388 25912 34428
rect 26712 34428 27660 34456
rect 27724 34428 59544 34456
rect 26712 34388 26740 34428
rect 27522 34388 27528 34400
rect 25884 34360 26740 34388
rect 27483 34360 27528 34388
rect 27522 34348 27528 34360
rect 27580 34348 27586 34400
rect 27632 34388 27660 34428
rect 59538 34416 59544 34428
rect 59596 34416 59602 34468
rect 65518 34456 65524 34468
rect 60568 34428 65524 34456
rect 36262 34388 36268 34400
rect 27632 34360 36268 34388
rect 36262 34348 36268 34360
rect 36320 34348 36326 34400
rect 36446 34388 36452 34400
rect 36359 34360 36452 34388
rect 36446 34348 36452 34360
rect 36504 34388 36510 34400
rect 37366 34388 37372 34400
rect 36504 34360 37372 34388
rect 36504 34348 36510 34360
rect 37366 34348 37372 34360
rect 37424 34388 37430 34400
rect 38194 34388 38200 34400
rect 37424 34360 38200 34388
rect 37424 34348 37430 34360
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 39390 34388 39396 34400
rect 39351 34360 39396 34388
rect 39390 34348 39396 34360
rect 39448 34348 39454 34400
rect 39482 34348 39488 34400
rect 39540 34388 39546 34400
rect 54389 34391 54447 34397
rect 54389 34388 54401 34391
rect 39540 34360 54401 34388
rect 39540 34348 39546 34360
rect 54389 34357 54401 34360
rect 54435 34388 54447 34391
rect 54570 34388 54576 34400
rect 54435 34360 54576 34388
rect 54435 34357 54447 34360
rect 54389 34351 54447 34357
rect 54570 34348 54576 34360
rect 54628 34348 54634 34400
rect 56042 34348 56048 34400
rect 56100 34388 56106 34400
rect 60568 34388 60596 34428
rect 65518 34416 65524 34428
rect 65576 34456 65582 34468
rect 65705 34459 65763 34465
rect 65705 34456 65717 34459
rect 65576 34428 65717 34456
rect 65576 34416 65582 34428
rect 65705 34425 65717 34428
rect 65751 34425 65763 34459
rect 65705 34419 65763 34425
rect 68756 34400 68784 34487
rect 68830 34484 68836 34536
rect 68888 34484 68894 34536
rect 68922 34484 68928 34536
rect 68980 34524 68986 34536
rect 75564 34533 75592 34632
rect 85390 34620 85396 34672
rect 85448 34660 85454 34672
rect 85485 34663 85543 34669
rect 85485 34660 85497 34663
rect 85448 34632 85497 34660
rect 85448 34620 85454 34632
rect 85485 34629 85497 34632
rect 85531 34629 85543 34663
rect 85485 34623 85543 34629
rect 75641 34595 75699 34601
rect 75641 34561 75653 34595
rect 75687 34592 75699 34595
rect 77110 34592 77116 34604
rect 75687 34564 77116 34592
rect 75687 34561 75699 34564
rect 75641 34555 75699 34561
rect 77110 34552 77116 34564
rect 77168 34552 77174 34604
rect 89441 34595 89499 34601
rect 89441 34592 89453 34595
rect 88168 34564 89453 34592
rect 69201 34527 69259 34533
rect 69201 34524 69213 34527
rect 68980 34496 69213 34524
rect 68980 34484 68986 34496
rect 69201 34493 69213 34496
rect 69247 34493 69259 34527
rect 69201 34487 69259 34493
rect 69293 34527 69351 34533
rect 69293 34493 69305 34527
rect 69339 34493 69351 34527
rect 69293 34487 69351 34493
rect 75549 34527 75607 34533
rect 75549 34493 75561 34527
rect 75595 34493 75607 34527
rect 75822 34524 75828 34536
rect 75783 34496 75828 34524
rect 75549 34487 75607 34493
rect 68848 34456 68876 34484
rect 69308 34456 69336 34487
rect 75822 34484 75828 34496
rect 75880 34484 75886 34536
rect 77018 34524 77024 34536
rect 76979 34496 77024 34524
rect 77018 34484 77024 34496
rect 77076 34484 77082 34536
rect 85022 34484 85028 34536
rect 85080 34524 85086 34536
rect 85393 34527 85451 34533
rect 85393 34524 85405 34527
rect 85080 34496 85405 34524
rect 85080 34484 85086 34496
rect 85393 34493 85405 34496
rect 85439 34493 85451 34527
rect 85393 34487 85451 34493
rect 85482 34484 85488 34536
rect 85540 34524 85546 34536
rect 88168 34533 88196 34564
rect 89441 34561 89453 34564
rect 89487 34561 89499 34595
rect 89441 34555 89499 34561
rect 88153 34527 88211 34533
rect 88153 34524 88165 34527
rect 85540 34496 88165 34524
rect 85540 34484 85546 34496
rect 88153 34493 88165 34496
rect 88199 34493 88211 34527
rect 88153 34487 88211 34493
rect 89349 34527 89407 34533
rect 89349 34493 89361 34527
rect 89395 34524 89407 34527
rect 89806 34524 89812 34536
rect 89395 34496 89812 34524
rect 89395 34493 89407 34496
rect 89349 34487 89407 34493
rect 89806 34484 89812 34496
rect 89864 34484 89870 34536
rect 68848 34428 69336 34456
rect 69400 34428 70164 34456
rect 62390 34388 62396 34400
rect 56100 34360 60596 34388
rect 62351 34360 62396 34388
rect 56100 34348 56106 34360
rect 62390 34348 62396 34360
rect 62448 34348 62454 34400
rect 68738 34388 68744 34400
rect 68651 34360 68744 34388
rect 68738 34348 68744 34360
rect 68796 34388 68802 34400
rect 69400 34388 69428 34428
rect 70136 34400 70164 34428
rect 76834 34416 76840 34468
rect 76892 34456 76898 34468
rect 76892 34428 76937 34456
rect 76892 34416 76898 34428
rect 87138 34416 87144 34468
rect 87196 34456 87202 34468
rect 87969 34459 88027 34465
rect 87969 34456 87981 34459
rect 87196 34428 87981 34456
rect 87196 34416 87202 34428
rect 87969 34425 87981 34428
rect 88015 34425 88027 34459
rect 88518 34456 88524 34468
rect 88479 34428 88524 34456
rect 87969 34419 88027 34425
rect 88518 34416 88524 34428
rect 88576 34416 88582 34468
rect 69750 34388 69756 34400
rect 68796 34360 69428 34388
rect 69711 34360 69756 34388
rect 68796 34348 68802 34360
rect 69750 34348 69756 34360
rect 69808 34348 69814 34400
rect 70118 34388 70124 34400
rect 70079 34360 70124 34388
rect 70118 34348 70124 34360
rect 70176 34348 70182 34400
rect 75822 34348 75828 34400
rect 75880 34388 75886 34400
rect 76101 34391 76159 34397
rect 76101 34388 76113 34391
rect 75880 34360 76113 34388
rect 75880 34348 75886 34360
rect 76101 34357 76113 34360
rect 76147 34357 76159 34391
rect 76101 34351 76159 34357
rect 76282 34348 76288 34400
rect 76340 34388 76346 34400
rect 88334 34388 88340 34400
rect 76340 34360 88340 34388
rect 76340 34348 76346 34360
rect 88334 34348 88340 34360
rect 88392 34348 88398 34400
rect 1104 34298 108008 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 81046 34298
rect 81098 34246 81110 34298
rect 81162 34246 81174 34298
rect 81226 34246 81238 34298
rect 81290 34246 108008 34298
rect 1104 34224 108008 34246
rect 2774 34144 2780 34196
rect 2832 34184 2838 34196
rect 4341 34187 4399 34193
rect 4341 34184 4353 34187
rect 2832 34156 4353 34184
rect 2832 34144 2838 34156
rect 4341 34153 4353 34156
rect 4387 34153 4399 34187
rect 4341 34147 4399 34153
rect 4356 34048 4384 34147
rect 4890 34144 4896 34196
rect 4948 34184 4954 34196
rect 5721 34187 5779 34193
rect 5721 34184 5733 34187
rect 4948 34156 5733 34184
rect 4948 34144 4954 34156
rect 5721 34153 5733 34156
rect 5767 34184 5779 34187
rect 6086 34184 6092 34196
rect 5767 34156 6092 34184
rect 5767 34153 5779 34156
rect 5721 34147 5779 34153
rect 6086 34144 6092 34156
rect 6144 34144 6150 34196
rect 9306 34184 9312 34196
rect 9267 34156 9312 34184
rect 9306 34144 9312 34156
rect 9364 34184 9370 34196
rect 11517 34187 11575 34193
rect 11517 34184 11529 34187
rect 9364 34156 11529 34184
rect 9364 34144 9370 34156
rect 11517 34153 11529 34156
rect 11563 34184 11575 34187
rect 11698 34184 11704 34196
rect 11563 34156 11704 34184
rect 11563 34153 11575 34156
rect 11517 34147 11575 34153
rect 11698 34144 11704 34156
rect 11756 34144 11762 34196
rect 13814 34144 13820 34196
rect 13872 34184 13878 34196
rect 16025 34187 16083 34193
rect 16025 34184 16037 34187
rect 13872 34156 16037 34184
rect 13872 34144 13878 34156
rect 16025 34153 16037 34156
rect 16071 34153 16083 34187
rect 16025 34147 16083 34153
rect 18966 34144 18972 34196
rect 19024 34184 19030 34196
rect 72418 34184 72424 34196
rect 19024 34156 72424 34184
rect 19024 34144 19030 34156
rect 72418 34144 72424 34156
rect 72476 34184 72482 34196
rect 75178 34184 75184 34196
rect 72476 34156 74672 34184
rect 75139 34156 75184 34184
rect 72476 34144 72482 34156
rect 16666 34116 16672 34128
rect 15672 34088 16672 34116
rect 4522 34048 4528 34060
rect 4356 34020 4528 34048
rect 4522 34008 4528 34020
rect 4580 34008 4586 34060
rect 4617 34051 4675 34057
rect 4617 34017 4629 34051
rect 4663 34048 4675 34051
rect 5537 34051 5595 34057
rect 5537 34048 5549 34051
rect 4663 34020 5549 34048
rect 4663 34017 4675 34020
rect 4617 34011 4675 34017
rect 5537 34017 5549 34020
rect 5583 34048 5595 34051
rect 7098 34048 7104 34060
rect 5583 34020 7104 34048
rect 5583 34017 5595 34020
rect 5537 34011 5595 34017
rect 7098 34008 7104 34020
rect 7156 34008 7162 34060
rect 9493 34051 9551 34057
rect 9493 34017 9505 34051
rect 9539 34048 9551 34051
rect 9582 34048 9588 34060
rect 9539 34020 9588 34048
rect 9539 34017 9551 34020
rect 9493 34011 9551 34017
rect 9582 34008 9588 34020
rect 9640 34008 9646 34060
rect 11977 34051 12035 34057
rect 11532 34020 11836 34048
rect 4890 33940 4896 33992
rect 4948 33980 4954 33992
rect 11532 33980 11560 34020
rect 11698 33980 11704 33992
rect 4948 33952 11560 33980
rect 11659 33952 11704 33980
rect 4948 33940 4954 33952
rect 11698 33940 11704 33952
rect 11756 33940 11762 33992
rect 11808 33980 11836 34020
rect 11977 34017 11989 34051
rect 12023 34048 12035 34051
rect 13170 34048 13176 34060
rect 12023 34020 13176 34048
rect 12023 34017 12035 34020
rect 11977 34011 12035 34017
rect 13170 34008 13176 34020
rect 13228 34008 13234 34060
rect 15562 34048 15568 34060
rect 15523 34020 15568 34048
rect 15562 34008 15568 34020
rect 15620 34008 15626 34060
rect 15672 34057 15700 34088
rect 16666 34076 16672 34088
rect 16724 34076 16730 34128
rect 27062 34116 27068 34128
rect 16776 34088 27068 34116
rect 15657 34051 15715 34057
rect 15657 34017 15669 34051
rect 15703 34017 15715 34051
rect 15657 34011 15715 34017
rect 15841 34051 15899 34057
rect 15841 34017 15853 34051
rect 15887 34048 15899 34051
rect 16482 34048 16488 34060
rect 15887 34020 16488 34048
rect 15887 34017 15899 34020
rect 15841 34011 15899 34017
rect 16482 34008 16488 34020
rect 16540 34008 16546 34060
rect 16776 33980 16804 34088
rect 27062 34076 27068 34088
rect 27120 34076 27126 34128
rect 27264 34088 27568 34116
rect 16850 34008 16856 34060
rect 16908 34048 16914 34060
rect 18414 34048 18420 34060
rect 16908 34020 18184 34048
rect 18375 34020 18420 34048
rect 16908 34008 16914 34020
rect 11808 33952 16804 33980
rect 17865 33983 17923 33989
rect 17865 33949 17877 33983
rect 17911 33980 17923 33983
rect 18046 33980 18052 33992
rect 17911 33952 18052 33980
rect 17911 33949 17923 33952
rect 17865 33943 17923 33949
rect 18046 33940 18052 33952
rect 18104 33940 18110 33992
rect 18156 33980 18184 34020
rect 18414 34008 18420 34020
rect 18472 34008 18478 34060
rect 18693 34051 18751 34057
rect 18693 34017 18705 34051
rect 18739 34048 18751 34051
rect 19061 34051 19119 34057
rect 19061 34048 19073 34051
rect 18739 34020 19073 34048
rect 18739 34017 18751 34020
rect 18693 34011 18751 34017
rect 19061 34017 19073 34020
rect 19107 34048 19119 34051
rect 21358 34048 21364 34060
rect 19107 34020 21364 34048
rect 19107 34017 19119 34020
rect 19061 34011 19119 34017
rect 21358 34008 21364 34020
rect 21416 34008 21422 34060
rect 21637 34051 21695 34057
rect 21637 34017 21649 34051
rect 21683 34048 21695 34051
rect 21729 34051 21787 34057
rect 21729 34048 21741 34051
rect 21683 34020 21741 34048
rect 21683 34017 21695 34020
rect 21637 34011 21695 34017
rect 21729 34017 21741 34020
rect 21775 34017 21787 34051
rect 25406 34048 25412 34060
rect 25367 34020 25412 34048
rect 21729 34011 21787 34017
rect 25406 34008 25412 34020
rect 25464 34008 25470 34060
rect 25501 34051 25559 34057
rect 25501 34017 25513 34051
rect 25547 34048 25559 34051
rect 26326 34048 26332 34060
rect 25547 34020 26332 34048
rect 25547 34017 25559 34020
rect 25501 34011 25559 34017
rect 26326 34008 26332 34020
rect 26384 34008 26390 34060
rect 26697 34051 26755 34057
rect 26697 34017 26709 34051
rect 26743 34048 26755 34051
rect 27154 34048 27160 34060
rect 26743 34020 27160 34048
rect 26743 34017 26755 34020
rect 26697 34011 26755 34017
rect 27154 34008 27160 34020
rect 27212 34048 27218 34060
rect 27264 34057 27292 34088
rect 27249 34051 27307 34057
rect 27249 34048 27261 34051
rect 27212 34020 27261 34048
rect 27212 34008 27218 34020
rect 27249 34017 27261 34020
rect 27295 34017 27307 34051
rect 27249 34011 27307 34017
rect 27338 34008 27344 34060
rect 27396 34048 27402 34060
rect 27433 34051 27491 34057
rect 27433 34048 27445 34051
rect 27396 34020 27445 34048
rect 27396 34008 27402 34020
rect 27433 34017 27445 34020
rect 27479 34017 27491 34051
rect 27540 34048 27568 34088
rect 27614 34076 27620 34128
rect 27672 34116 27678 34128
rect 37182 34116 37188 34128
rect 27672 34088 36584 34116
rect 37143 34088 37188 34116
rect 27672 34076 27678 34088
rect 28077 34051 28135 34057
rect 28077 34048 28089 34051
rect 27540 34020 28089 34048
rect 27433 34011 27491 34017
rect 28077 34017 28089 34020
rect 28123 34048 28135 34051
rect 28261 34051 28319 34057
rect 28261 34048 28273 34051
rect 28123 34020 28273 34048
rect 28123 34017 28135 34020
rect 28077 34011 28135 34017
rect 28261 34017 28273 34020
rect 28307 34048 28319 34051
rect 29270 34048 29276 34060
rect 28307 34020 29276 34048
rect 28307 34017 28319 34020
rect 28261 34011 28319 34017
rect 29270 34008 29276 34020
rect 29328 34008 29334 34060
rect 32122 34048 32128 34060
rect 32083 34020 32128 34048
rect 32122 34008 32128 34020
rect 32180 34008 32186 34060
rect 18877 33983 18935 33989
rect 18877 33980 18889 33983
rect 18156 33952 18889 33980
rect 18877 33949 18889 33952
rect 18923 33949 18935 33983
rect 25424 33980 25452 34008
rect 26050 33980 26056 33992
rect 18877 33943 18935 33949
rect 19076 33952 23520 33980
rect 25424 33952 26056 33980
rect 16390 33872 16396 33924
rect 16448 33912 16454 33924
rect 19076 33912 19104 33952
rect 21910 33912 21916 33924
rect 16448 33884 19104 33912
rect 21871 33884 21916 33912
rect 16448 33872 16454 33884
rect 21910 33872 21916 33884
rect 21968 33872 21974 33924
rect 23492 33912 23520 33952
rect 26050 33940 26056 33952
rect 26108 33940 26114 33992
rect 26234 33940 26240 33992
rect 26292 33980 26298 33992
rect 26513 33983 26571 33989
rect 26513 33980 26525 33983
rect 26292 33952 26525 33980
rect 26292 33940 26298 33952
rect 26513 33949 26525 33952
rect 26559 33949 26571 33983
rect 35526 33980 35532 33992
rect 26513 33943 26571 33949
rect 27632 33952 35532 33980
rect 27632 33912 27660 33952
rect 35526 33940 35532 33952
rect 35584 33940 35590 33992
rect 23492 33884 27660 33912
rect 27798 33872 27804 33924
rect 27856 33912 27862 33924
rect 36446 33912 36452 33924
rect 27856 33884 36452 33912
rect 27856 33872 27862 33884
rect 36446 33872 36452 33884
rect 36504 33872 36510 33924
rect 36556 33912 36584 34088
rect 37182 34076 37188 34088
rect 37240 34116 37246 34128
rect 37369 34119 37427 34125
rect 37369 34116 37381 34119
rect 37240 34088 37381 34116
rect 37240 34076 37246 34088
rect 37369 34085 37381 34088
rect 37415 34116 37427 34119
rect 37415 34088 37964 34116
rect 37415 34085 37427 34088
rect 37369 34079 37427 34085
rect 37936 34057 37964 34088
rect 38746 34076 38752 34128
rect 38804 34116 38810 34128
rect 39025 34119 39083 34125
rect 39025 34116 39037 34119
rect 38804 34088 39037 34116
rect 38804 34076 38810 34088
rect 39025 34085 39037 34088
rect 39071 34085 39083 34119
rect 39025 34079 39083 34085
rect 50617 34119 50675 34125
rect 50617 34085 50629 34119
rect 50663 34116 50675 34119
rect 50982 34116 50988 34128
rect 50663 34088 50988 34116
rect 50663 34085 50675 34088
rect 50617 34079 50675 34085
rect 50982 34076 50988 34088
rect 51040 34076 51046 34128
rect 56778 34116 56784 34128
rect 56739 34088 56784 34116
rect 56778 34076 56784 34088
rect 56836 34116 56842 34128
rect 58253 34119 58311 34125
rect 56836 34088 57008 34116
rect 56836 34076 56842 34088
rect 37921 34051 37979 34057
rect 37921 34017 37933 34051
rect 37967 34048 37979 34051
rect 38473 34051 38531 34057
rect 38473 34048 38485 34051
rect 37967 34020 38485 34048
rect 37967 34017 37979 34020
rect 37921 34011 37979 34017
rect 38473 34017 38485 34020
rect 38519 34017 38531 34051
rect 38473 34011 38531 34017
rect 38657 34051 38715 34057
rect 38657 34017 38669 34051
rect 38703 34048 38715 34051
rect 38838 34048 38844 34060
rect 38703 34020 38844 34048
rect 38703 34017 38715 34020
rect 38657 34011 38715 34017
rect 38838 34008 38844 34020
rect 38896 34048 38902 34060
rect 39390 34048 39396 34060
rect 38896 34020 39396 34048
rect 38896 34008 38902 34020
rect 39390 34008 39396 34020
rect 39448 34008 39454 34060
rect 41340 34020 43484 34048
rect 37553 33983 37611 33989
rect 37553 33949 37565 33983
rect 37599 33980 37611 33983
rect 37737 33983 37795 33989
rect 37737 33980 37749 33983
rect 37599 33952 37749 33980
rect 37599 33949 37611 33952
rect 37553 33943 37611 33949
rect 37737 33949 37749 33952
rect 37783 33949 37795 33983
rect 37737 33943 37795 33949
rect 41340 33912 41368 34020
rect 36556 33884 41368 33912
rect 4982 33804 4988 33856
rect 5040 33844 5046 33856
rect 13081 33847 13139 33853
rect 13081 33844 13093 33847
rect 5040 33816 13093 33844
rect 5040 33804 5046 33816
rect 13081 33813 13093 33816
rect 13127 33844 13139 33847
rect 13906 33844 13912 33856
rect 13127 33816 13912 33844
rect 13127 33813 13139 33816
rect 13081 33807 13139 33813
rect 13906 33804 13912 33816
rect 13964 33804 13970 33856
rect 16482 33844 16488 33856
rect 16395 33816 16488 33844
rect 16482 33804 16488 33816
rect 16540 33844 16546 33856
rect 17218 33844 17224 33856
rect 16540 33816 17224 33844
rect 16540 33804 16546 33816
rect 17218 33804 17224 33816
rect 17276 33844 17282 33856
rect 17954 33844 17960 33856
rect 17276 33816 17960 33844
rect 17276 33804 17282 33816
rect 17954 33804 17960 33816
rect 18012 33804 18018 33856
rect 19886 33804 19892 33856
rect 19944 33844 19950 33856
rect 21637 33847 21695 33853
rect 21637 33844 21649 33847
rect 19944 33816 21649 33844
rect 19944 33804 19950 33816
rect 21637 33813 21649 33816
rect 21683 33813 21695 33847
rect 21637 33807 21695 33813
rect 27706 33804 27712 33856
rect 27764 33844 27770 33856
rect 27764 33816 27809 33844
rect 27764 33804 27770 33816
rect 31202 33804 31208 33856
rect 31260 33844 31266 33856
rect 32030 33844 32036 33856
rect 31260 33816 32036 33844
rect 31260 33804 31266 33816
rect 32030 33804 32036 33816
rect 32088 33844 32094 33856
rect 32217 33847 32275 33853
rect 32217 33844 32229 33847
rect 32088 33816 32229 33844
rect 32088 33804 32094 33816
rect 32217 33813 32229 33816
rect 32263 33813 32275 33847
rect 32217 33807 32275 33813
rect 32858 33804 32864 33856
rect 32916 33844 32922 33856
rect 37001 33847 37059 33853
rect 37001 33844 37013 33847
rect 32916 33816 37013 33844
rect 32916 33804 32922 33816
rect 37001 33813 37013 33816
rect 37047 33844 37059 33847
rect 37553 33847 37611 33853
rect 37553 33844 37565 33847
rect 37047 33816 37565 33844
rect 37047 33813 37059 33816
rect 37001 33807 37059 33813
rect 37553 33813 37565 33816
rect 37599 33844 37611 33847
rect 42886 33844 42892 33856
rect 37599 33816 42892 33844
rect 37599 33813 37611 33816
rect 37553 33807 37611 33813
rect 42886 33804 42892 33816
rect 42944 33804 42950 33856
rect 43456 33844 43484 34020
rect 44266 34008 44272 34060
rect 44324 34048 44330 34060
rect 44637 34051 44695 34057
rect 44637 34048 44649 34051
rect 44324 34020 44649 34048
rect 44324 34008 44330 34020
rect 44637 34017 44649 34020
rect 44683 34017 44695 34051
rect 49513 34051 49571 34057
rect 49513 34048 49525 34051
rect 44637 34011 44695 34017
rect 49436 34020 49525 34048
rect 43806 33940 43812 33992
rect 43864 33980 43870 33992
rect 44361 33983 44419 33989
rect 44361 33980 44373 33983
rect 43864 33952 44373 33980
rect 43864 33940 43870 33952
rect 44361 33949 44373 33952
rect 44407 33949 44419 33983
rect 44361 33943 44419 33949
rect 45554 33940 45560 33992
rect 45612 33980 45618 33992
rect 45741 33983 45799 33989
rect 45741 33980 45753 33983
rect 45612 33952 45753 33980
rect 45612 33940 45618 33952
rect 45741 33949 45753 33952
rect 45787 33949 45799 33983
rect 45741 33943 45799 33949
rect 49329 33983 49387 33989
rect 49329 33949 49341 33983
rect 49375 33949 49387 33983
rect 49329 33943 49387 33949
rect 48685 33915 48743 33921
rect 48685 33912 48697 33915
rect 45296 33884 48697 33912
rect 45296 33844 45324 33884
rect 48685 33881 48697 33884
rect 48731 33912 48743 33915
rect 49234 33912 49240 33924
rect 48731 33884 49240 33912
rect 48731 33881 48743 33884
rect 48685 33875 48743 33881
rect 49234 33872 49240 33884
rect 49292 33912 49298 33924
rect 49344 33912 49372 33943
rect 49292 33884 49372 33912
rect 49436 33912 49464 34020
rect 49513 34017 49525 34020
rect 49559 34048 49571 34051
rect 50065 34051 50123 34057
rect 50065 34048 50077 34051
rect 49559 34020 50077 34048
rect 49559 34017 49571 34020
rect 49513 34011 49571 34017
rect 50065 34017 50077 34020
rect 50111 34017 50123 34051
rect 50065 34011 50123 34017
rect 50154 34008 50160 34060
rect 50212 34048 50218 34060
rect 50249 34051 50307 34057
rect 50249 34048 50261 34051
rect 50212 34020 50261 34048
rect 50212 34008 50218 34020
rect 50249 34017 50261 34020
rect 50295 34048 50307 34051
rect 50706 34048 50712 34060
rect 50295 34020 50712 34048
rect 50295 34017 50307 34020
rect 50249 34011 50307 34017
rect 50706 34008 50712 34020
rect 50764 34008 50770 34060
rect 54757 34051 54815 34057
rect 54757 34048 54769 34051
rect 54220 34020 54769 34048
rect 54220 33921 54248 34020
rect 54757 34017 54769 34020
rect 54803 34048 54815 34051
rect 55309 34051 55367 34057
rect 55309 34048 55321 34051
rect 54803 34020 55321 34048
rect 54803 34017 54815 34020
rect 54757 34011 54815 34017
rect 55309 34017 55321 34020
rect 55355 34017 55367 34051
rect 55490 34048 55496 34060
rect 55451 34020 55496 34048
rect 55309 34011 55367 34017
rect 55490 34008 55496 34020
rect 55548 34048 55554 34060
rect 56042 34048 56048 34060
rect 55548 34020 56048 34048
rect 55548 34008 55554 34020
rect 56042 34008 56048 34020
rect 56100 34008 56106 34060
rect 56980 34057 57008 34088
rect 57072 34088 57928 34116
rect 56965 34051 57023 34057
rect 56965 34017 56977 34051
rect 57011 34017 57023 34051
rect 56965 34011 57023 34017
rect 54570 33980 54576 33992
rect 54531 33952 54576 33980
rect 54570 33940 54576 33952
rect 54628 33940 54634 33992
rect 56686 33980 56692 33992
rect 56599 33952 56692 33980
rect 56686 33940 56692 33952
rect 56744 33980 56750 33992
rect 57072 33980 57100 34088
rect 57149 34051 57207 34057
rect 57149 34017 57161 34051
rect 57195 34048 57207 34051
rect 57514 34048 57520 34060
rect 57195 34020 57520 34048
rect 57195 34017 57207 34020
rect 57149 34011 57207 34017
rect 57514 34008 57520 34020
rect 57572 34008 57578 34060
rect 57698 34048 57704 34060
rect 57659 34020 57704 34048
rect 57698 34008 57704 34020
rect 57756 34008 57762 34060
rect 57900 34057 57928 34088
rect 58253 34085 58265 34119
rect 58299 34116 58311 34119
rect 63126 34116 63132 34128
rect 58299 34088 63132 34116
rect 58299 34085 58311 34088
rect 58253 34079 58311 34085
rect 63126 34076 63132 34088
rect 63184 34076 63190 34128
rect 64693 34119 64751 34125
rect 64693 34085 64705 34119
rect 64739 34116 64751 34119
rect 65978 34116 65984 34128
rect 64739 34088 65984 34116
rect 64739 34085 64751 34088
rect 64693 34079 64751 34085
rect 65978 34076 65984 34088
rect 66036 34076 66042 34128
rect 74537 34119 74595 34125
rect 74537 34116 74549 34119
rect 73264 34088 74549 34116
rect 73264 34060 73292 34088
rect 74537 34085 74549 34088
rect 74583 34085 74595 34119
rect 74644 34116 74672 34156
rect 75178 34144 75184 34156
rect 75236 34184 75242 34196
rect 75730 34184 75736 34196
rect 75236 34156 75736 34184
rect 75236 34144 75242 34156
rect 75730 34144 75736 34156
rect 75788 34144 75794 34196
rect 82906 34184 82912 34196
rect 75840 34156 82912 34184
rect 75840 34116 75868 34156
rect 82906 34144 82912 34156
rect 82964 34144 82970 34196
rect 87966 34184 87972 34196
rect 87927 34156 87972 34184
rect 87966 34144 87972 34156
rect 88024 34144 88030 34196
rect 74644 34088 75868 34116
rect 74537 34079 74595 34085
rect 77110 34076 77116 34128
rect 77168 34116 77174 34128
rect 85022 34116 85028 34128
rect 77168 34088 77340 34116
rect 84983 34088 85028 34116
rect 77168 34076 77174 34088
rect 57885 34051 57943 34057
rect 57885 34017 57897 34051
rect 57931 34017 57943 34051
rect 63313 34051 63371 34057
rect 63313 34048 63325 34051
rect 57885 34011 57943 34017
rect 58268 34020 63325 34048
rect 56744 33952 57100 33980
rect 56744 33940 56750 33952
rect 54021 33915 54079 33921
rect 54021 33912 54033 33915
rect 49436 33884 54033 33912
rect 49292 33872 49298 33884
rect 43456 33816 45324 33844
rect 46842 33804 46848 33856
rect 46900 33844 46906 33856
rect 48961 33847 49019 33853
rect 48961 33844 48973 33847
rect 46900 33816 48973 33844
rect 46900 33804 46906 33816
rect 48961 33813 48973 33816
rect 49007 33844 49019 33847
rect 49145 33847 49203 33853
rect 49145 33844 49157 33847
rect 49007 33816 49157 33844
rect 49007 33813 49019 33816
rect 48961 33807 49019 33813
rect 49145 33813 49157 33816
rect 49191 33844 49203 33847
rect 49436 33844 49464 33884
rect 54021 33881 54033 33884
rect 54067 33912 54079 33915
rect 54205 33915 54263 33921
rect 54205 33912 54217 33915
rect 54067 33884 54217 33912
rect 54067 33881 54079 33884
rect 54021 33875 54079 33881
rect 54205 33881 54217 33884
rect 54251 33881 54263 33915
rect 54205 33875 54263 33881
rect 55769 33915 55827 33921
rect 55769 33881 55781 33915
rect 55815 33912 55827 33915
rect 58268 33912 58296 34020
rect 63313 34017 63325 34020
rect 63359 34017 63371 34051
rect 67453 34051 67511 34057
rect 67453 34048 67465 34051
rect 63313 34011 63371 34017
rect 64156 34020 67465 34048
rect 60918 33940 60924 33992
rect 60976 33980 60982 33992
rect 61286 33980 61292 33992
rect 60976 33952 61292 33980
rect 60976 33940 60982 33952
rect 61286 33940 61292 33952
rect 61344 33980 61350 33992
rect 62853 33983 62911 33989
rect 62853 33980 62865 33983
rect 61344 33952 62865 33980
rect 61344 33940 61350 33952
rect 62853 33949 62865 33952
rect 62899 33980 62911 33983
rect 63037 33983 63095 33989
rect 63037 33980 63049 33983
rect 62899 33952 63049 33980
rect 62899 33949 62911 33952
rect 62853 33943 62911 33949
rect 63037 33949 63049 33952
rect 63083 33949 63095 33983
rect 63037 33943 63095 33949
rect 55815 33884 58296 33912
rect 55815 33881 55827 33884
rect 55769 33875 55827 33881
rect 58434 33872 58440 33924
rect 58492 33912 58498 33924
rect 58492 33884 63080 33912
rect 58492 33872 58498 33884
rect 49191 33816 49464 33844
rect 49191 33813 49203 33816
rect 49145 33807 49203 33813
rect 57698 33804 57704 33856
rect 57756 33844 57762 33856
rect 58526 33844 58532 33856
rect 57756 33816 58532 33844
rect 57756 33804 57762 33816
rect 58526 33804 58532 33816
rect 58584 33804 58590 33856
rect 58618 33804 58624 33856
rect 58676 33844 58682 33856
rect 63052 33844 63080 33884
rect 64156 33844 64184 34020
rect 67453 34017 67465 34020
rect 67499 34017 67511 34051
rect 68925 34051 68983 34057
rect 68925 34048 68937 34051
rect 67453 34011 67511 34017
rect 67928 34020 68937 34048
rect 67177 33983 67235 33989
rect 67177 33949 67189 33983
rect 67223 33980 67235 33983
rect 67634 33980 67640 33992
rect 67223 33952 67640 33980
rect 67223 33949 67235 33952
rect 67177 33943 67235 33949
rect 67634 33940 67640 33952
rect 67692 33980 67698 33992
rect 67928 33980 67956 34020
rect 68925 34017 68937 34020
rect 68971 34017 68983 34051
rect 73246 34048 73252 34060
rect 73207 34020 73252 34048
rect 68925 34011 68983 34017
rect 73246 34008 73252 34020
rect 73304 34008 73310 34060
rect 73985 34051 74043 34057
rect 73985 34017 73997 34051
rect 74031 34048 74043 34051
rect 74442 34048 74448 34060
rect 74031 34020 74448 34048
rect 74031 34017 74043 34020
rect 73985 34011 74043 34017
rect 74442 34008 74448 34020
rect 74500 34048 74506 34060
rect 75365 34051 75423 34057
rect 75365 34048 75377 34051
rect 74500 34020 75377 34048
rect 74500 34008 74506 34020
rect 75365 34017 75377 34020
rect 75411 34017 75423 34051
rect 75365 34011 75423 34017
rect 75546 34008 75552 34060
rect 75604 34048 75610 34060
rect 77312 34057 77340 34088
rect 85022 34076 85028 34088
rect 85080 34076 85086 34128
rect 77205 34051 77263 34057
rect 77205 34048 77217 34051
rect 75604 34020 77217 34048
rect 75604 34008 75610 34020
rect 77205 34017 77217 34020
rect 77251 34017 77263 34051
rect 77205 34011 77263 34017
rect 77297 34051 77355 34057
rect 77297 34017 77309 34051
rect 77343 34017 77355 34051
rect 87138 34048 87144 34060
rect 87099 34020 87144 34048
rect 77297 34011 77355 34017
rect 87138 34008 87144 34020
rect 87196 34008 87202 34060
rect 87414 34008 87420 34060
rect 87472 34048 87478 34060
rect 87984 34048 88012 34144
rect 88245 34051 88303 34057
rect 88245 34048 88257 34051
rect 87472 34020 88257 34048
rect 87472 34008 87478 34020
rect 88245 34017 88257 34020
rect 88291 34017 88303 34051
rect 88426 34048 88432 34060
rect 88387 34020 88432 34048
rect 88245 34011 88303 34017
rect 88426 34008 88432 34020
rect 88484 34008 88490 34060
rect 88518 34008 88524 34060
rect 88576 34048 88582 34060
rect 89806 34048 89812 34060
rect 88576 34020 88621 34048
rect 89767 34020 89812 34048
rect 88576 34008 88582 34020
rect 89806 34008 89812 34020
rect 89864 34008 89870 34060
rect 68554 33980 68560 33992
rect 67692 33952 67956 33980
rect 68515 33952 68560 33980
rect 67692 33940 67698 33952
rect 68554 33940 68560 33952
rect 68612 33940 68618 33992
rect 74258 33980 74264 33992
rect 74171 33952 74264 33980
rect 74258 33940 74264 33952
rect 74316 33980 74322 33992
rect 75564 33980 75592 34008
rect 75730 33980 75736 33992
rect 74316 33952 75592 33980
rect 75691 33952 75736 33980
rect 74316 33940 74322 33952
rect 75730 33940 75736 33952
rect 75788 33940 75794 33992
rect 76101 33983 76159 33989
rect 76101 33949 76113 33983
rect 76147 33980 76159 33983
rect 78674 33980 78680 33992
rect 76147 33952 78680 33980
rect 76147 33949 76159 33952
rect 76101 33943 76159 33949
rect 78674 33940 78680 33952
rect 78732 33940 78738 33992
rect 83369 33983 83427 33989
rect 83369 33980 83381 33983
rect 83200 33952 83381 33980
rect 73525 33915 73583 33921
rect 73525 33881 73537 33915
rect 73571 33912 73583 33915
rect 73982 33912 73988 33924
rect 73571 33884 73988 33912
rect 73571 33881 73583 33884
rect 73525 33875 73583 33881
rect 73982 33872 73988 33884
rect 74040 33872 74046 33924
rect 75641 33915 75699 33921
rect 75641 33881 75653 33915
rect 75687 33912 75699 33915
rect 76834 33912 76840 33924
rect 75687 33884 76840 33912
rect 75687 33881 75699 33884
rect 75641 33875 75699 33881
rect 76834 33872 76840 33884
rect 76892 33872 76898 33924
rect 77021 33915 77079 33921
rect 77021 33881 77033 33915
rect 77067 33912 77079 33915
rect 77202 33912 77208 33924
rect 77067 33884 77208 33912
rect 77067 33881 77079 33884
rect 77021 33875 77079 33881
rect 77202 33872 77208 33884
rect 77260 33872 77266 33924
rect 83200 33856 83228 33952
rect 83369 33949 83381 33952
rect 83415 33949 83427 33983
rect 83369 33943 83427 33949
rect 83645 33983 83703 33989
rect 83645 33949 83657 33983
rect 83691 33980 83703 33983
rect 85482 33980 85488 33992
rect 83691 33952 85488 33980
rect 83691 33949 83703 33952
rect 83645 33943 83703 33949
rect 85482 33940 85488 33952
rect 85540 33940 85546 33992
rect 88334 33872 88340 33924
rect 88392 33912 88398 33924
rect 89993 33915 90051 33921
rect 89993 33912 90005 33915
rect 88392 33884 90005 33912
rect 88392 33872 88398 33884
rect 89993 33881 90005 33884
rect 90039 33881 90051 33915
rect 89993 33875 90051 33881
rect 75546 33853 75552 33856
rect 58676 33816 58721 33844
rect 63052 33816 64184 33844
rect 75530 33847 75552 33853
rect 58676 33804 58682 33816
rect 75530 33813 75542 33847
rect 75604 33844 75610 33856
rect 75822 33844 75828 33856
rect 75604 33816 75828 33844
rect 75530 33807 75552 33813
rect 75546 33804 75552 33807
rect 75604 33804 75610 33816
rect 75822 33804 75828 33816
rect 75880 33844 75886 33856
rect 76193 33847 76251 33853
rect 76193 33844 76205 33847
rect 75880 33816 76205 33844
rect 75880 33804 75886 33816
rect 76193 33813 76205 33816
rect 76239 33813 76251 33847
rect 77478 33844 77484 33856
rect 77439 33816 77484 33844
rect 76193 33807 76251 33813
rect 77478 33804 77484 33816
rect 77536 33804 77542 33856
rect 83182 33844 83188 33856
rect 83143 33816 83188 33844
rect 83182 33804 83188 33816
rect 83240 33804 83246 33856
rect 87230 33844 87236 33856
rect 87191 33816 87236 33844
rect 87230 33804 87236 33816
rect 87288 33804 87294 33856
rect 88518 33804 88524 33856
rect 88576 33844 88582 33856
rect 88705 33847 88763 33853
rect 88705 33844 88717 33847
rect 88576 33816 88717 33844
rect 88576 33804 88582 33816
rect 88705 33813 88717 33816
rect 88751 33813 88763 33847
rect 88705 33807 88763 33813
rect 1104 33754 108008 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 65686 33754
rect 65738 33702 65750 33754
rect 65802 33702 65814 33754
rect 65866 33702 65878 33754
rect 65930 33702 96406 33754
rect 96458 33702 96470 33754
rect 96522 33702 96534 33754
rect 96586 33702 96598 33754
rect 96650 33702 108008 33754
rect 1104 33680 108008 33702
rect 4433 33643 4491 33649
rect 4433 33640 4445 33643
rect 2608 33612 4445 33640
rect 2608 33513 2636 33612
rect 4433 33609 4445 33612
rect 4479 33640 4491 33643
rect 4706 33640 4712 33652
rect 4479 33612 4712 33640
rect 4479 33609 4491 33612
rect 4433 33603 4491 33609
rect 4706 33600 4712 33612
rect 4764 33600 4770 33652
rect 22738 33600 22744 33652
rect 22796 33640 22802 33652
rect 46934 33640 46940 33652
rect 22796 33612 46940 33640
rect 22796 33600 22802 33612
rect 46934 33600 46940 33612
rect 46992 33600 46998 33652
rect 49234 33640 49240 33652
rect 49195 33612 49240 33640
rect 49234 33600 49240 33612
rect 49292 33600 49298 33652
rect 50617 33643 50675 33649
rect 50617 33609 50629 33643
rect 50663 33640 50675 33643
rect 50798 33640 50804 33652
rect 50663 33612 50804 33640
rect 50663 33609 50675 33612
rect 50617 33603 50675 33609
rect 50798 33600 50804 33612
rect 50856 33600 50862 33652
rect 50982 33600 50988 33652
rect 51040 33640 51046 33652
rect 53929 33643 53987 33649
rect 51040 33612 51396 33640
rect 51040 33600 51046 33612
rect 9306 33532 9312 33584
rect 9364 33572 9370 33584
rect 9677 33575 9735 33581
rect 9677 33572 9689 33575
rect 9364 33544 9689 33572
rect 9364 33532 9370 33544
rect 9677 33541 9689 33544
rect 9723 33572 9735 33575
rect 12894 33572 12900 33584
rect 9723 33544 12900 33572
rect 9723 33541 9735 33544
rect 9677 33535 9735 33541
rect 12894 33532 12900 33544
rect 12952 33532 12958 33584
rect 14918 33532 14924 33584
rect 14976 33572 14982 33584
rect 15013 33575 15071 33581
rect 15013 33572 15025 33575
rect 14976 33544 15025 33572
rect 14976 33532 14982 33544
rect 15013 33541 15025 33544
rect 15059 33541 15071 33575
rect 17310 33572 17316 33584
rect 17271 33544 17316 33572
rect 15013 33535 15071 33541
rect 17310 33532 17316 33544
rect 17368 33532 17374 33584
rect 18141 33575 18199 33581
rect 18141 33541 18153 33575
rect 18187 33572 18199 33575
rect 18966 33572 18972 33584
rect 18187 33544 18972 33572
rect 18187 33541 18199 33544
rect 18141 33535 18199 33541
rect 18966 33532 18972 33544
rect 19024 33532 19030 33584
rect 24670 33532 24676 33584
rect 24728 33572 24734 33584
rect 24857 33575 24915 33581
rect 24857 33572 24869 33575
rect 24728 33544 24869 33572
rect 24728 33532 24734 33544
rect 24857 33541 24869 33544
rect 24903 33541 24915 33575
rect 24857 33535 24915 33541
rect 26050 33532 26056 33584
rect 26108 33572 26114 33584
rect 26329 33575 26387 33581
rect 26329 33572 26341 33575
rect 26108 33544 26341 33572
rect 26108 33532 26114 33544
rect 26329 33541 26341 33544
rect 26375 33541 26387 33575
rect 32122 33572 32128 33584
rect 32083 33544 32128 33572
rect 26329 33535 26387 33541
rect 32122 33532 32128 33544
rect 32180 33532 32186 33584
rect 33134 33572 33140 33584
rect 33095 33544 33140 33572
rect 33134 33532 33140 33544
rect 33192 33532 33198 33584
rect 36262 33532 36268 33584
rect 36320 33572 36326 33584
rect 38746 33572 38752 33584
rect 36320 33544 38752 33572
rect 36320 33532 36326 33544
rect 38746 33532 38752 33544
rect 38804 33532 38810 33584
rect 2593 33507 2651 33513
rect 2593 33473 2605 33507
rect 2639 33473 2651 33507
rect 2593 33467 2651 33473
rect 2869 33507 2927 33513
rect 2869 33473 2881 33507
rect 2915 33504 2927 33507
rect 3602 33504 3608 33516
rect 2915 33476 3608 33504
rect 2915 33473 2927 33476
rect 2869 33467 2927 33473
rect 3602 33464 3608 33476
rect 3660 33464 3666 33516
rect 3970 33464 3976 33516
rect 4028 33504 4034 33516
rect 19242 33504 19248 33516
rect 4028 33476 19248 33504
rect 4028 33464 4034 33476
rect 19242 33464 19248 33476
rect 19300 33464 19306 33516
rect 19334 33464 19340 33516
rect 19392 33504 19398 33516
rect 32858 33504 32864 33516
rect 19392 33476 32864 33504
rect 19392 33464 19398 33476
rect 32858 33464 32864 33476
rect 32916 33464 32922 33516
rect 35526 33464 35532 33516
rect 35584 33504 35590 33516
rect 37277 33507 37335 33513
rect 37277 33504 37289 33507
rect 35584 33476 37289 33504
rect 35584 33464 35590 33476
rect 37277 33473 37289 33476
rect 37323 33473 37335 33507
rect 37277 33467 37335 33473
rect 38013 33507 38071 33513
rect 38013 33473 38025 33507
rect 38059 33504 38071 33507
rect 38654 33504 38660 33516
rect 38059 33476 38660 33504
rect 38059 33473 38071 33476
rect 38013 33467 38071 33473
rect 38654 33464 38660 33476
rect 38712 33464 38718 33516
rect 49234 33464 49240 33516
rect 49292 33504 49298 33516
rect 51368 33513 51396 33612
rect 53929 33609 53941 33643
rect 53975 33640 53987 33643
rect 54570 33640 54576 33652
rect 53975 33612 54576 33640
rect 53975 33609 53987 33612
rect 53929 33603 53987 33609
rect 54570 33600 54576 33612
rect 54628 33600 54634 33652
rect 56870 33640 56876 33652
rect 56831 33612 56876 33640
rect 56870 33600 56876 33612
rect 56928 33600 56934 33652
rect 57514 33600 57520 33652
rect 57572 33640 57578 33652
rect 58618 33640 58624 33652
rect 57572 33612 58624 33640
rect 57572 33600 57578 33612
rect 58618 33600 58624 33612
rect 58676 33640 58682 33652
rect 58989 33643 59047 33649
rect 58989 33640 59001 33643
rect 58676 33612 59001 33640
rect 58676 33600 58682 33612
rect 58989 33609 59001 33612
rect 59035 33609 59047 33643
rect 68002 33640 68008 33652
rect 58989 33603 59047 33609
rect 59096 33612 68008 33640
rect 55490 33572 55496 33584
rect 54404 33544 55496 33572
rect 49421 33507 49479 33513
rect 49421 33504 49433 33507
rect 49292 33476 49433 33504
rect 49292 33464 49298 33476
rect 49421 33473 49433 33476
rect 49467 33473 49479 33507
rect 49421 33467 49479 33473
rect 51353 33507 51411 33513
rect 51353 33473 51365 33507
rect 51399 33504 51411 33507
rect 52549 33507 52607 33513
rect 51399 33476 52500 33504
rect 51399 33473 51411 33476
rect 51353 33467 51411 33473
rect 7098 33396 7104 33448
rect 7156 33436 7162 33448
rect 7377 33439 7435 33445
rect 7377 33436 7389 33439
rect 7156 33408 7389 33436
rect 7156 33396 7162 33408
rect 7377 33405 7389 33408
rect 7423 33405 7435 33439
rect 8757 33439 8815 33445
rect 8757 33436 8769 33439
rect 7377 33399 7435 33405
rect 8036 33408 8769 33436
rect 8036 33312 8064 33408
rect 8757 33405 8769 33408
rect 8803 33405 8815 33439
rect 9306 33436 9312 33448
rect 9267 33408 9312 33436
rect 8757 33399 8815 33405
rect 9306 33396 9312 33408
rect 9364 33396 9370 33448
rect 14918 33396 14924 33448
rect 14976 33436 14982 33448
rect 15197 33439 15255 33445
rect 15197 33436 15209 33439
rect 14976 33408 15209 33436
rect 14976 33396 14982 33408
rect 15197 33405 15209 33408
rect 15243 33405 15255 33439
rect 15197 33399 15255 33405
rect 15289 33439 15347 33445
rect 15289 33405 15301 33439
rect 15335 33436 15347 33439
rect 16206 33436 16212 33448
rect 15335 33408 16212 33436
rect 15335 33405 15347 33408
rect 15289 33399 15347 33405
rect 16206 33396 16212 33408
rect 16264 33436 16270 33448
rect 16577 33439 16635 33445
rect 16577 33436 16589 33439
rect 16264 33408 16589 33436
rect 16264 33396 16270 33408
rect 16577 33405 16589 33408
rect 16623 33436 16635 33439
rect 16666 33436 16672 33448
rect 16623 33408 16672 33436
rect 16623 33405 16635 33408
rect 16577 33399 16635 33405
rect 16666 33396 16672 33408
rect 16724 33396 16730 33448
rect 16761 33439 16819 33445
rect 16761 33405 16773 33439
rect 16807 33436 16819 33439
rect 17310 33436 17316 33448
rect 16807 33408 17316 33436
rect 16807 33405 16819 33408
rect 16761 33399 16819 33405
rect 17310 33396 17316 33408
rect 17368 33396 17374 33448
rect 18046 33436 18052 33448
rect 18007 33408 18052 33436
rect 18046 33396 18052 33408
rect 18104 33396 18110 33448
rect 18322 33436 18328 33448
rect 18283 33408 18328 33436
rect 18322 33396 18328 33408
rect 18380 33396 18386 33448
rect 19886 33436 19892 33448
rect 19847 33408 19892 33436
rect 19886 33396 19892 33408
rect 19944 33396 19950 33448
rect 21358 33396 21364 33448
rect 21416 33436 21422 33448
rect 24854 33436 24860 33448
rect 21416 33408 24860 33436
rect 21416 33396 21422 33408
rect 24854 33396 24860 33408
rect 24912 33396 24918 33448
rect 24949 33439 25007 33445
rect 24949 33405 24961 33439
rect 24995 33405 25007 33439
rect 24949 33399 25007 33405
rect 25225 33439 25283 33445
rect 25225 33405 25237 33439
rect 25271 33436 25283 33439
rect 26050 33436 26056 33448
rect 25271 33408 26056 33436
rect 25271 33405 25283 33408
rect 25225 33399 25283 33405
rect 8938 33328 8944 33380
rect 8996 33368 9002 33380
rect 8996 33340 24072 33368
rect 8996 33328 9002 33340
rect 4154 33300 4160 33312
rect 4115 33272 4160 33300
rect 4154 33260 4160 33272
rect 4212 33260 4218 33312
rect 7561 33303 7619 33309
rect 7561 33269 7573 33303
rect 7607 33300 7619 33303
rect 8018 33300 8024 33312
rect 7607 33272 8024 33300
rect 7607 33269 7619 33272
rect 7561 33263 7619 33269
rect 8018 33260 8024 33272
rect 8076 33260 8082 33312
rect 9033 33303 9091 33309
rect 9033 33269 9045 33303
rect 9079 33300 9091 33303
rect 9214 33300 9220 33312
rect 9079 33272 9220 33300
rect 9079 33269 9091 33272
rect 9033 33263 9091 33269
rect 9214 33260 9220 33272
rect 9272 33260 9278 33312
rect 10778 33260 10784 33312
rect 10836 33300 10842 33312
rect 16390 33300 16396 33312
rect 10836 33272 16396 33300
rect 10836 33260 10842 33272
rect 16390 33260 16396 33272
rect 16448 33260 16454 33312
rect 16482 33260 16488 33312
rect 16540 33300 16546 33312
rect 16853 33303 16911 33309
rect 16853 33300 16865 33303
rect 16540 33272 16865 33300
rect 16540 33260 16546 33272
rect 16853 33269 16865 33272
rect 16899 33269 16911 33303
rect 16853 33263 16911 33269
rect 17865 33303 17923 33309
rect 17865 33269 17877 33303
rect 17911 33300 17923 33303
rect 17954 33300 17960 33312
rect 17911 33272 17960 33300
rect 17911 33269 17923 33272
rect 17865 33263 17923 33269
rect 17954 33260 17960 33272
rect 18012 33300 18018 33312
rect 18322 33300 18328 33312
rect 18012 33272 18328 33300
rect 18012 33260 18018 33272
rect 18322 33260 18328 33272
rect 18380 33260 18386 33312
rect 18506 33300 18512 33312
rect 18467 33272 18512 33300
rect 18506 33260 18512 33272
rect 18564 33260 18570 33312
rect 19978 33300 19984 33312
rect 19939 33272 19984 33300
rect 19978 33260 19984 33272
rect 20036 33260 20042 33312
rect 24044 33300 24072 33340
rect 24118 33328 24124 33380
rect 24176 33368 24182 33380
rect 24670 33368 24676 33380
rect 24176 33340 24676 33368
rect 24176 33328 24182 33340
rect 24670 33328 24676 33340
rect 24728 33368 24734 33380
rect 24964 33368 24992 33399
rect 26050 33396 26056 33408
rect 26108 33396 26114 33448
rect 27433 33439 27491 33445
rect 27433 33405 27445 33439
rect 27479 33436 27491 33439
rect 27614 33436 27620 33448
rect 27479 33408 27620 33436
rect 27479 33405 27491 33408
rect 27433 33399 27491 33405
rect 27614 33396 27620 33408
rect 27672 33396 27678 33448
rect 30558 33436 30564 33448
rect 30519 33408 30564 33436
rect 30558 33396 30564 33408
rect 30616 33396 30622 33448
rect 30834 33396 30840 33448
rect 30892 33436 30898 33448
rect 33045 33439 33103 33445
rect 30892 33408 30937 33436
rect 30892 33396 30898 33408
rect 33045 33405 33057 33439
rect 33091 33436 33103 33439
rect 33226 33436 33232 33448
rect 33091 33408 33232 33436
rect 33091 33405 33103 33408
rect 33045 33399 33103 33405
rect 33226 33396 33232 33408
rect 33284 33396 33290 33448
rect 35434 33436 35440 33448
rect 35395 33408 35440 33436
rect 35434 33396 35440 33408
rect 35492 33436 35498 33448
rect 35621 33439 35679 33445
rect 35621 33436 35633 33439
rect 35492 33408 35633 33436
rect 35492 33396 35498 33408
rect 35621 33405 35633 33408
rect 35667 33405 35679 33439
rect 35621 33399 35679 33405
rect 37001 33439 37059 33445
rect 37001 33405 37013 33439
rect 37047 33436 37059 33439
rect 37366 33436 37372 33448
rect 37047 33408 37372 33436
rect 37047 33405 37059 33408
rect 37001 33399 37059 33405
rect 37366 33396 37372 33408
rect 37424 33436 37430 33448
rect 37921 33439 37979 33445
rect 37921 33436 37933 33439
rect 37424 33408 37933 33436
rect 37424 33396 37430 33408
rect 37921 33405 37933 33408
rect 37967 33405 37979 33439
rect 38286 33436 38292 33448
rect 38247 33408 38292 33436
rect 37921 33399 37979 33405
rect 38286 33396 38292 33408
rect 38344 33396 38350 33448
rect 38473 33439 38531 33445
rect 38473 33405 38485 33439
rect 38519 33436 38531 33439
rect 38519 33408 38700 33436
rect 38519 33405 38531 33408
rect 38473 33399 38531 33405
rect 24728 33340 24992 33368
rect 25884 33340 27660 33368
rect 24728 33328 24734 33340
rect 25884 33300 25912 33340
rect 24044 33272 25912 33300
rect 27246 33260 27252 33312
rect 27304 33300 27310 33312
rect 27522 33300 27528 33312
rect 27304 33272 27528 33300
rect 27304 33260 27310 33272
rect 27522 33260 27528 33272
rect 27580 33260 27586 33312
rect 27632 33300 27660 33340
rect 27706 33328 27712 33380
rect 27764 33368 27770 33380
rect 30650 33368 30656 33380
rect 27764 33340 30656 33368
rect 27764 33328 27770 33340
rect 30650 33328 30656 33340
rect 30708 33328 30714 33380
rect 38562 33368 38568 33380
rect 32048 33340 38568 33368
rect 32048 33300 32076 33340
rect 38562 33328 38568 33340
rect 38620 33328 38626 33380
rect 38672 33368 38700 33408
rect 41874 33396 41880 33448
rect 41932 33436 41938 33448
rect 46842 33436 46848 33448
rect 41932 33408 46848 33436
rect 41932 33396 41938 33408
rect 46842 33396 46848 33408
rect 46900 33396 46906 33448
rect 49605 33439 49663 33445
rect 49605 33436 49617 33439
rect 49068 33408 49617 33436
rect 38838 33368 38844 33380
rect 38672 33340 38844 33368
rect 38838 33328 38844 33340
rect 38896 33328 38902 33380
rect 27632 33272 32076 33300
rect 32122 33260 32128 33312
rect 32180 33300 32186 33312
rect 32306 33300 32312 33312
rect 32180 33272 32312 33300
rect 32180 33260 32186 33272
rect 32306 33260 32312 33272
rect 32364 33260 32370 33312
rect 33226 33260 33232 33312
rect 33284 33300 33290 33312
rect 33321 33303 33379 33309
rect 33321 33300 33333 33303
rect 33284 33272 33333 33300
rect 33284 33260 33290 33272
rect 33321 33269 33333 33272
rect 33367 33269 33379 33303
rect 33321 33263 33379 33269
rect 35805 33303 35863 33309
rect 35805 33269 35817 33303
rect 35851 33300 35863 33303
rect 37185 33303 37243 33309
rect 37185 33300 37197 33303
rect 35851 33272 37197 33300
rect 35851 33269 35863 33272
rect 35805 33263 35863 33269
rect 37185 33269 37197 33272
rect 37231 33300 37243 33303
rect 38286 33300 38292 33312
rect 37231 33272 38292 33300
rect 37231 33269 37243 33272
rect 37185 33263 37243 33269
rect 38286 33260 38292 33272
rect 38344 33260 38350 33312
rect 42334 33260 42340 33312
rect 42392 33300 42398 33312
rect 49068 33309 49096 33408
rect 49605 33405 49617 33408
rect 49651 33436 49663 33439
rect 50157 33439 50215 33445
rect 50157 33436 50169 33439
rect 49651 33408 50169 33436
rect 49651 33405 49663 33408
rect 49605 33399 49663 33405
rect 50157 33405 50169 33408
rect 50203 33436 50215 33439
rect 50341 33439 50399 33445
rect 50203 33408 50292 33436
rect 50203 33405 50215 33408
rect 50157 33399 50215 33405
rect 48869 33303 48927 33309
rect 48869 33300 48881 33303
rect 42392 33272 48881 33300
rect 42392 33260 42398 33272
rect 48869 33269 48881 33272
rect 48915 33300 48927 33303
rect 49053 33303 49111 33309
rect 49053 33300 49065 33303
rect 48915 33272 49065 33300
rect 48915 33269 48927 33272
rect 48869 33263 48927 33269
rect 49053 33269 49065 33272
rect 49099 33269 49111 33303
rect 50264 33300 50292 33408
rect 50341 33405 50353 33439
rect 50387 33436 50399 33439
rect 51166 33436 51172 33448
rect 50387 33408 51172 33436
rect 50387 33405 50399 33408
rect 50341 33399 50399 33405
rect 51166 33396 51172 33408
rect 51224 33396 51230 33448
rect 52472 33445 52500 33476
rect 52549 33473 52561 33507
rect 52595 33504 52607 33507
rect 53285 33507 53343 33513
rect 53285 33504 53297 33507
rect 52595 33476 53297 33504
rect 52595 33473 52607 33476
rect 52549 33467 52607 33473
rect 53285 33473 53297 33476
rect 53331 33504 53343 33507
rect 54404 33504 54432 33544
rect 55490 33532 55496 33544
rect 55548 33532 55554 33584
rect 53331 33476 54432 33504
rect 55309 33507 55367 33513
rect 53331 33473 53343 33476
rect 53285 33467 53343 33473
rect 55309 33473 55321 33507
rect 55355 33473 55367 33507
rect 56888 33504 56916 33600
rect 58434 33572 58440 33584
rect 57440 33544 58440 33572
rect 57333 33507 57391 33513
rect 57333 33504 57345 33507
rect 56888 33476 57345 33504
rect 55309 33467 55367 33473
rect 57333 33473 57345 33476
rect 57379 33473 57391 33507
rect 57333 33467 57391 33473
rect 52457 33439 52515 33445
rect 51460 33408 52040 33436
rect 51460 33380 51488 33408
rect 51442 33368 51448 33380
rect 51403 33340 51448 33368
rect 51442 33328 51448 33340
rect 51500 33328 51506 33380
rect 51810 33368 51816 33380
rect 51771 33340 51816 33368
rect 51810 33328 51816 33340
rect 51868 33328 51874 33380
rect 52012 33368 52040 33408
rect 52457 33405 52469 33439
rect 52503 33405 52515 33439
rect 52822 33436 52828 33448
rect 52735 33408 52828 33436
rect 52457 33399 52515 33405
rect 52822 33396 52828 33408
rect 52880 33396 52886 33448
rect 53006 33436 53012 33448
rect 52967 33408 53012 33436
rect 53006 33396 53012 33408
rect 53064 33396 53070 33448
rect 54205 33439 54263 33445
rect 54205 33405 54217 33439
rect 54251 33405 54263 33439
rect 54205 33399 54263 33405
rect 54297 33439 54355 33445
rect 54297 33405 54309 33439
rect 54343 33436 54355 33439
rect 54570 33436 54576 33448
rect 54343 33408 54576 33436
rect 54343 33405 54355 33408
rect 54297 33399 54355 33405
rect 52840 33368 52868 33396
rect 53469 33371 53527 33377
rect 53469 33368 53481 33371
rect 52012 33340 52868 33368
rect 52932 33340 53481 33368
rect 52932 33300 52960 33340
rect 53469 33337 53481 33340
rect 53515 33368 53527 33371
rect 53653 33371 53711 33377
rect 53653 33368 53665 33371
rect 53515 33340 53665 33368
rect 53515 33337 53527 33340
rect 53469 33331 53527 33337
rect 53653 33337 53665 33340
rect 53699 33368 53711 33371
rect 54220 33368 54248 33399
rect 54570 33396 54576 33408
rect 54628 33396 54634 33448
rect 54757 33439 54815 33445
rect 54757 33405 54769 33439
rect 54803 33405 54815 33439
rect 54757 33399 54815 33405
rect 54941 33439 54999 33445
rect 54941 33405 54953 33439
rect 54987 33405 54999 33439
rect 55324 33436 55352 33467
rect 57440 33436 57468 33544
rect 58434 33532 58440 33544
rect 58492 33532 58498 33584
rect 55324 33408 57468 33436
rect 54941 33399 54999 33405
rect 54772 33368 54800 33399
rect 53699 33340 54800 33368
rect 54956 33368 54984 33399
rect 57514 33396 57520 33448
rect 57572 33436 57578 33448
rect 57977 33439 58035 33445
rect 57977 33436 57989 33439
rect 57572 33408 57617 33436
rect 57716 33408 57989 33436
rect 57572 33396 57578 33408
rect 57054 33368 57060 33380
rect 54956 33340 55628 33368
rect 56967 33340 57060 33368
rect 53699 33337 53711 33340
rect 53653 33331 53711 33337
rect 50264 33272 52960 33300
rect 49053 33263 49111 33269
rect 53006 33260 53012 33312
rect 53064 33300 53070 33312
rect 53193 33303 53251 33309
rect 53193 33300 53205 33303
rect 53064 33272 53205 33300
rect 53064 33260 53070 33272
rect 53193 33269 53205 33272
rect 53239 33300 53251 33303
rect 54956 33300 54984 33340
rect 55600 33309 55628 33340
rect 57054 33328 57060 33340
rect 57112 33368 57118 33380
rect 57716 33368 57744 33408
rect 57977 33405 57989 33408
rect 58023 33405 58035 33439
rect 57977 33399 58035 33405
rect 58157 33439 58215 33445
rect 58157 33405 58169 33439
rect 58203 33405 58215 33439
rect 58157 33399 58215 33405
rect 58066 33368 58072 33380
rect 57112 33340 57744 33368
rect 57808 33340 58072 33368
rect 57112 33328 57118 33340
rect 53239 33272 54984 33300
rect 55585 33303 55643 33309
rect 53239 33269 53251 33272
rect 53193 33263 53251 33269
rect 55585 33269 55597 33303
rect 55631 33300 55643 33303
rect 57808 33300 57836 33340
rect 58066 33328 58072 33340
rect 58124 33328 58130 33380
rect 55631 33272 57836 33300
rect 58176 33300 58204 33399
rect 58250 33396 58256 33448
rect 58308 33436 58314 33448
rect 59096 33436 59124 33612
rect 68002 33600 68008 33612
rect 68060 33600 68066 33652
rect 68722 33643 68780 33649
rect 68722 33609 68734 33643
rect 68768 33640 68780 33643
rect 69474 33640 69480 33652
rect 68768 33612 69480 33640
rect 68768 33609 68780 33612
rect 68722 33603 68780 33609
rect 69474 33600 69480 33612
rect 69532 33600 69538 33652
rect 85482 33640 85488 33652
rect 85443 33612 85488 33640
rect 85482 33600 85488 33612
rect 85540 33600 85546 33652
rect 87049 33643 87107 33649
rect 87049 33609 87061 33643
rect 87095 33640 87107 33643
rect 87138 33640 87144 33652
rect 87095 33612 87144 33640
rect 87095 33609 87107 33612
rect 87049 33603 87107 33609
rect 87138 33600 87144 33612
rect 87196 33600 87202 33652
rect 89806 33640 89812 33652
rect 89767 33612 89812 33640
rect 89806 33600 89812 33612
rect 89864 33600 89870 33652
rect 60921 33575 60979 33581
rect 60921 33541 60933 33575
rect 60967 33572 60979 33575
rect 61654 33572 61660 33584
rect 60967 33544 61660 33572
rect 60967 33541 60979 33544
rect 60921 33535 60979 33541
rect 61654 33532 61660 33544
rect 61712 33532 61718 33584
rect 68833 33575 68891 33581
rect 68833 33541 68845 33575
rect 68879 33572 68891 33575
rect 69658 33572 69664 33584
rect 68879 33544 69664 33572
rect 68879 33541 68891 33544
rect 68833 33535 68891 33541
rect 69658 33532 69664 33544
rect 69716 33532 69722 33584
rect 61013 33507 61071 33513
rect 61013 33473 61025 33507
rect 61059 33504 61071 33507
rect 62574 33504 62580 33516
rect 61059 33476 62580 33504
rect 61059 33473 61071 33476
rect 61013 33467 61071 33473
rect 62574 33464 62580 33476
rect 62632 33464 62638 33516
rect 68925 33507 68983 33513
rect 68925 33473 68937 33507
rect 68971 33504 68983 33507
rect 69750 33504 69756 33516
rect 68971 33476 69756 33504
rect 68971 33473 68983 33476
rect 68925 33467 68983 33473
rect 69750 33464 69756 33476
rect 69808 33464 69814 33516
rect 76285 33507 76343 33513
rect 76285 33473 76297 33507
rect 76331 33504 76343 33507
rect 77478 33504 77484 33516
rect 76331 33476 77484 33504
rect 76331 33473 76343 33476
rect 76285 33467 76343 33473
rect 77478 33464 77484 33476
rect 77536 33464 77542 33516
rect 80793 33507 80851 33513
rect 80793 33473 80805 33507
rect 80839 33504 80851 33507
rect 80885 33507 80943 33513
rect 80885 33504 80897 33507
rect 80839 33476 80897 33504
rect 80839 33473 80851 33476
rect 80793 33467 80851 33473
rect 80885 33473 80897 33476
rect 80931 33504 80943 33507
rect 83182 33504 83188 33516
rect 80931 33476 83188 33504
rect 80931 33473 80943 33476
rect 80885 33467 80943 33473
rect 58308 33408 59124 33436
rect 60792 33439 60850 33445
rect 58308 33396 58314 33408
rect 60792 33405 60804 33439
rect 60838 33436 60850 33439
rect 61102 33436 61108 33448
rect 60838 33408 61108 33436
rect 60838 33405 60850 33408
rect 60792 33399 60850 33405
rect 61102 33396 61108 33408
rect 61160 33396 61166 33448
rect 61378 33436 61384 33448
rect 61339 33408 61384 33436
rect 61378 33396 61384 33408
rect 61436 33396 61442 33448
rect 69290 33436 69296 33448
rect 69251 33408 69296 33436
rect 69290 33396 69296 33408
rect 69348 33396 69354 33448
rect 75914 33396 75920 33448
rect 75972 33436 75978 33448
rect 76009 33439 76067 33445
rect 76009 33436 76021 33439
rect 75972 33408 76021 33436
rect 75972 33396 75978 33408
rect 76009 33405 76021 33408
rect 76055 33436 76067 33439
rect 77294 33436 77300 33448
rect 76055 33408 77300 33436
rect 76055 33405 76067 33408
rect 76009 33399 76067 33405
rect 77294 33396 77300 33408
rect 77352 33436 77358 33448
rect 77754 33436 77760 33448
rect 77352 33408 77760 33436
rect 77352 33396 77358 33408
rect 77754 33396 77760 33408
rect 77812 33436 77818 33448
rect 80808 33436 80836 33467
rect 83182 33464 83188 33476
rect 83240 33504 83246 33516
rect 88518 33504 88524 33516
rect 83240 33476 88104 33504
rect 88479 33476 88524 33504
rect 83240 33464 83246 33476
rect 77812 33408 80836 33436
rect 81161 33439 81219 33445
rect 77812 33396 77818 33408
rect 81161 33405 81173 33439
rect 81207 33436 81219 33439
rect 81526 33436 81532 33448
rect 81207 33408 81532 33436
rect 81207 33405 81219 33408
rect 81161 33399 81219 33405
rect 81526 33396 81532 33408
rect 81584 33396 81590 33448
rect 85393 33439 85451 33445
rect 85393 33405 85405 33439
rect 85439 33436 85451 33439
rect 85666 33436 85672 33448
rect 85439 33408 85672 33436
rect 85439 33405 85451 33408
rect 85393 33399 85451 33405
rect 85666 33396 85672 33408
rect 85724 33396 85730 33448
rect 86957 33439 87015 33445
rect 86957 33436 86969 33439
rect 86696 33408 86969 33436
rect 58621 33371 58679 33377
rect 58621 33337 58633 33371
rect 58667 33368 58679 33371
rect 60645 33371 60703 33377
rect 60645 33368 60657 33371
rect 58667 33340 60657 33368
rect 58667 33337 58679 33340
rect 58621 33331 58679 33337
rect 60645 33337 60657 33340
rect 60691 33337 60703 33371
rect 60645 33331 60703 33337
rect 63126 33328 63132 33380
rect 63184 33368 63190 33380
rect 68557 33371 68615 33377
rect 68557 33368 68569 33371
rect 63184 33340 68569 33368
rect 63184 33328 63190 33340
rect 68557 33337 68569 33340
rect 68603 33337 68615 33371
rect 75546 33368 75552 33380
rect 68557 33331 68615 33337
rect 68664 33340 75552 33368
rect 58526 33300 58532 33312
rect 58176 33272 58532 33300
rect 55631 33269 55643 33272
rect 55585 33263 55643 33269
rect 58526 33260 58532 33272
rect 58584 33300 58590 33312
rect 58897 33303 58955 33309
rect 58897 33300 58909 33303
rect 58584 33272 58909 33300
rect 58584 33260 58590 33272
rect 58897 33269 58909 33272
rect 58943 33300 58955 33303
rect 68664 33300 68692 33340
rect 75546 33328 75552 33340
rect 75604 33328 75610 33380
rect 86696 33312 86724 33408
rect 86957 33405 86969 33408
rect 87003 33405 87015 33439
rect 86957 33399 87015 33405
rect 88076 33436 88104 33476
rect 88518 33464 88524 33476
rect 88576 33464 88582 33516
rect 88245 33439 88303 33445
rect 88245 33436 88257 33439
rect 88076 33408 88257 33436
rect 86770 33328 86776 33380
rect 86828 33368 86834 33380
rect 86828 33340 86873 33368
rect 86828 33328 86834 33340
rect 77386 33300 77392 33312
rect 58943 33272 68692 33300
rect 77347 33272 77392 33300
rect 58943 33269 58955 33272
rect 58897 33263 58955 33269
rect 77386 33260 77392 33272
rect 77444 33260 77450 33312
rect 82262 33300 82268 33312
rect 82223 33272 82268 33300
rect 82262 33260 82268 33272
rect 82320 33260 82326 33312
rect 86678 33300 86684 33312
rect 86639 33272 86684 33300
rect 86678 33260 86684 33272
rect 86736 33260 86742 33312
rect 87966 33260 87972 33312
rect 88024 33300 88030 33312
rect 88076 33309 88104 33408
rect 88245 33405 88257 33408
rect 88291 33405 88303 33439
rect 88245 33399 88303 33405
rect 88061 33303 88119 33309
rect 88061 33300 88073 33303
rect 88024 33272 88073 33300
rect 88024 33260 88030 33272
rect 88061 33269 88073 33272
rect 88107 33269 88119 33303
rect 88061 33263 88119 33269
rect 1104 33210 108008 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 50326 33210
rect 50378 33158 50390 33210
rect 50442 33158 50454 33210
rect 50506 33158 50518 33210
rect 50570 33158 81046 33210
rect 81098 33158 81110 33210
rect 81162 33158 81174 33210
rect 81226 33158 81238 33210
rect 81290 33158 108008 33210
rect 1104 33136 108008 33158
rect 3786 33056 3792 33108
rect 3844 33096 3850 33108
rect 7558 33096 7564 33108
rect 3844 33068 7564 33096
rect 3844 33056 3850 33068
rect 7558 33056 7564 33068
rect 7616 33056 7622 33108
rect 8938 33096 8944 33108
rect 8899 33068 8944 33096
rect 8938 33056 8944 33068
rect 8996 33056 9002 33108
rect 10597 33099 10655 33105
rect 10597 33065 10609 33099
rect 10643 33096 10655 33099
rect 49421 33099 49479 33105
rect 49421 33096 49433 33099
rect 10643 33068 49433 33096
rect 10643 33065 10655 33068
rect 10597 33059 10655 33065
rect 49421 33065 49433 33068
rect 49467 33065 49479 33099
rect 49421 33059 49479 33065
rect 8036 33000 9720 33028
rect 8036 32972 8064 33000
rect 8018 32960 8024 32972
rect 7979 32932 8024 32960
rect 8018 32920 8024 32932
rect 8076 32920 8082 32972
rect 8573 32963 8631 32969
rect 8573 32929 8585 32963
rect 8619 32960 8631 32963
rect 8938 32960 8944 32972
rect 8619 32932 8944 32960
rect 8619 32929 8631 32932
rect 8573 32923 8631 32929
rect 8938 32920 8944 32932
rect 8996 32920 9002 32972
rect 9692 32969 9720 33000
rect 9677 32963 9735 32969
rect 9677 32929 9689 32963
rect 9723 32929 9735 32963
rect 9677 32923 9735 32929
rect 10229 32963 10287 32969
rect 10229 32929 10241 32963
rect 10275 32960 10287 32963
rect 10612 32960 10640 33059
rect 62022 33056 62028 33108
rect 62080 33096 62086 33108
rect 63681 33099 63739 33105
rect 63681 33096 63693 33099
rect 62080 33068 63693 33096
rect 62080 33056 62086 33068
rect 63681 33065 63693 33068
rect 63727 33065 63739 33099
rect 63681 33059 63739 33065
rect 11698 32988 11704 33040
rect 11756 33028 11762 33040
rect 15013 33031 15071 33037
rect 15013 33028 15025 33031
rect 11756 33000 15025 33028
rect 11756 32988 11762 33000
rect 15013 32997 15025 33000
rect 15059 33028 15071 33031
rect 17865 33031 17923 33037
rect 15059 33000 15332 33028
rect 15059 32997 15071 33000
rect 15013 32991 15071 32997
rect 15304 32969 15332 33000
rect 17865 32997 17877 33031
rect 17911 33028 17923 33031
rect 18414 33028 18420 33040
rect 17911 33000 18420 33028
rect 17911 32997 17923 33000
rect 17865 32991 17923 32997
rect 18414 32988 18420 33000
rect 18472 32988 18478 33040
rect 24854 32988 24860 33040
rect 24912 33028 24918 33040
rect 25314 33028 25320 33040
rect 24912 33000 25320 33028
rect 24912 32988 24918 33000
rect 25314 32988 25320 33000
rect 25372 33028 25378 33040
rect 27706 33028 27712 33040
rect 25372 33000 27712 33028
rect 25372 32988 25378 33000
rect 27706 32988 27712 33000
rect 27764 32988 27770 33040
rect 29270 33028 29276 33040
rect 29231 33000 29276 33028
rect 29270 32988 29276 33000
rect 29328 33028 29334 33040
rect 29365 33031 29423 33037
rect 29365 33028 29377 33031
rect 29328 33000 29377 33028
rect 29328 32988 29334 33000
rect 29365 32997 29377 33000
rect 29411 33028 29423 33031
rect 29411 33000 30512 33028
rect 29411 32997 29423 33000
rect 29365 32991 29423 32997
rect 10275 32932 10640 32960
rect 15289 32963 15347 32969
rect 10275 32929 10287 32932
rect 10229 32923 10287 32929
rect 15289 32929 15301 32963
rect 15335 32929 15347 32963
rect 17773 32963 17831 32969
rect 17773 32960 17785 32963
rect 15289 32923 15347 32929
rect 17604 32932 17785 32960
rect 8662 32892 8668 32904
rect 8623 32864 8668 32892
rect 8662 32852 8668 32864
rect 8720 32852 8726 32904
rect 10410 32892 10416 32904
rect 10371 32864 10416 32892
rect 10410 32852 10416 32864
rect 10468 32852 10474 32904
rect 15565 32895 15623 32901
rect 15565 32861 15577 32895
rect 15611 32892 15623 32895
rect 16850 32892 16856 32904
rect 15611 32864 16856 32892
rect 15611 32861 15623 32864
rect 15565 32855 15623 32861
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 16666 32756 16672 32768
rect 16627 32728 16672 32756
rect 16666 32716 16672 32728
rect 16724 32756 16730 32768
rect 17604 32765 17632 32932
rect 17773 32929 17785 32932
rect 17819 32929 17831 32963
rect 19610 32960 19616 32972
rect 19571 32932 19616 32960
rect 17773 32923 17831 32929
rect 19610 32920 19616 32932
rect 19668 32960 19674 32972
rect 20901 32963 20959 32969
rect 20901 32960 20913 32963
rect 19668 32932 20913 32960
rect 19668 32920 19674 32932
rect 20901 32929 20913 32932
rect 20947 32929 20959 32963
rect 20901 32923 20959 32929
rect 21542 32920 21548 32972
rect 21600 32960 21606 32972
rect 29932 32969 29960 33000
rect 30484 32969 30512 33000
rect 30834 32988 30840 33040
rect 30892 33028 30898 33040
rect 31021 33031 31079 33037
rect 31021 33028 31033 33031
rect 30892 33000 31033 33028
rect 30892 32988 30898 33000
rect 31021 32997 31033 33000
rect 31067 32997 31079 33031
rect 31570 33028 31576 33040
rect 31021 32991 31079 32997
rect 31312 33000 31576 33028
rect 29917 32963 29975 32969
rect 21600 32932 29868 32960
rect 21600 32920 21606 32932
rect 25222 32852 25228 32904
rect 25280 32892 25286 32904
rect 26142 32892 26148 32904
rect 25280 32864 26148 32892
rect 25280 32852 25286 32864
rect 26142 32852 26148 32864
rect 26200 32852 26206 32904
rect 29733 32895 29791 32901
rect 29733 32892 29745 32895
rect 29564 32864 29745 32892
rect 19797 32827 19855 32833
rect 19797 32793 19809 32827
rect 19843 32824 19855 32827
rect 20622 32824 20628 32836
rect 19843 32796 20628 32824
rect 19843 32793 19855 32796
rect 19797 32787 19855 32793
rect 20622 32784 20628 32796
rect 20680 32784 20686 32836
rect 21085 32827 21143 32833
rect 21085 32793 21097 32827
rect 21131 32824 21143 32827
rect 23750 32824 23756 32836
rect 21131 32796 23756 32824
rect 21131 32793 21143 32796
rect 21085 32787 21143 32793
rect 23750 32784 23756 32796
rect 23808 32784 23814 32836
rect 17589 32759 17647 32765
rect 17589 32756 17601 32759
rect 16724 32728 17601 32756
rect 16724 32716 16730 32728
rect 17589 32725 17601 32728
rect 17635 32725 17647 32759
rect 17589 32719 17647 32725
rect 24302 32716 24308 32768
rect 24360 32756 24366 32768
rect 29564 32765 29592 32864
rect 29733 32861 29745 32864
rect 29779 32861 29791 32895
rect 29840 32892 29868 32932
rect 29917 32929 29929 32963
rect 29963 32929 29975 32963
rect 30377 32963 30435 32969
rect 30377 32960 30389 32963
rect 29917 32923 29975 32929
rect 30116 32932 30389 32960
rect 30116 32892 30144 32932
rect 30377 32929 30389 32932
rect 30423 32929 30435 32963
rect 30377 32923 30435 32929
rect 30469 32963 30527 32969
rect 30469 32929 30481 32963
rect 30515 32929 30527 32963
rect 30469 32923 30527 32929
rect 30558 32920 30564 32972
rect 30616 32960 30622 32972
rect 31312 32960 31340 33000
rect 31570 32988 31576 33000
rect 31628 33028 31634 33040
rect 32122 33028 32128 33040
rect 31628 33000 32128 33028
rect 31628 32988 31634 33000
rect 32122 32988 32128 33000
rect 32180 32988 32186 33040
rect 33134 33028 33140 33040
rect 33060 33000 33140 33028
rect 30616 32932 31340 32960
rect 30616 32920 30622 32932
rect 31386 32920 31392 32972
rect 31444 32960 31450 32972
rect 33060 32969 33088 33000
rect 33134 32988 33140 33000
rect 33192 32988 33198 33040
rect 49142 33028 49148 33040
rect 49103 33000 49148 33028
rect 49142 32988 49148 33000
rect 49200 33028 49206 33040
rect 51442 33028 51448 33040
rect 49200 33000 51448 33028
rect 49200 32988 49206 33000
rect 31849 32963 31907 32969
rect 31849 32960 31861 32963
rect 31444 32932 31861 32960
rect 31444 32920 31450 32932
rect 31849 32929 31861 32932
rect 31895 32960 31907 32963
rect 32309 32963 32367 32969
rect 32309 32960 32321 32963
rect 31895 32932 32321 32960
rect 31895 32929 31907 32932
rect 31849 32923 31907 32929
rect 32309 32929 32321 32932
rect 32355 32929 32367 32963
rect 32861 32963 32919 32969
rect 32861 32960 32873 32963
rect 32309 32923 32367 32929
rect 32508 32932 32873 32960
rect 29840 32864 30144 32892
rect 29733 32855 29791 32861
rect 30116 32824 30144 32864
rect 31481 32895 31539 32901
rect 31481 32861 31493 32895
rect 31527 32892 31539 32895
rect 32125 32895 32183 32901
rect 32125 32892 32137 32895
rect 31527 32864 32137 32892
rect 31527 32861 31539 32864
rect 31481 32855 31539 32861
rect 32125 32861 32137 32864
rect 32171 32861 32183 32895
rect 32125 32855 32183 32861
rect 31202 32824 31208 32836
rect 30116 32796 31208 32824
rect 31202 32784 31208 32796
rect 31260 32784 31266 32836
rect 32508 32824 32536 32932
rect 32861 32929 32873 32932
rect 32907 32929 32919 32963
rect 32861 32923 32919 32929
rect 33045 32963 33103 32969
rect 33045 32929 33057 32963
rect 33091 32929 33103 32963
rect 33045 32923 33103 32929
rect 37918 32920 37924 32972
rect 37976 32960 37982 32972
rect 38105 32963 38163 32969
rect 38105 32960 38117 32963
rect 37976 32932 38117 32960
rect 37976 32920 37982 32932
rect 38105 32929 38117 32932
rect 38151 32929 38163 32963
rect 38105 32923 38163 32929
rect 41966 32920 41972 32972
rect 42024 32960 42030 32972
rect 42153 32963 42211 32969
rect 42153 32960 42165 32963
rect 42024 32932 42165 32960
rect 42024 32920 42030 32932
rect 42153 32929 42165 32932
rect 42199 32929 42211 32963
rect 42153 32923 42211 32929
rect 45465 32963 45523 32969
rect 45465 32929 45477 32963
rect 45511 32960 45523 32963
rect 46293 32963 46351 32969
rect 46293 32960 46305 32963
rect 45511 32932 46305 32960
rect 45511 32929 45523 32932
rect 45465 32923 45523 32929
rect 46293 32929 46305 32932
rect 46339 32929 46351 32963
rect 46293 32923 46351 32929
rect 49053 32963 49111 32969
rect 49053 32929 49065 32963
rect 49099 32960 49111 32963
rect 49694 32960 49700 32972
rect 49099 32932 49700 32960
rect 49099 32929 49111 32932
rect 49053 32923 49111 32929
rect 49694 32920 49700 32932
rect 49752 32960 49758 32972
rect 50356 32969 50384 33000
rect 51442 32988 51448 33000
rect 51500 32988 51506 33040
rect 49973 32963 50031 32969
rect 49973 32960 49985 32963
rect 49752 32932 49985 32960
rect 49752 32920 49758 32932
rect 49973 32929 49985 32932
rect 50019 32960 50031 32963
rect 50341 32963 50399 32969
rect 50019 32932 50292 32960
rect 50019 32929 50031 32932
rect 49973 32923 50031 32929
rect 43438 32852 43444 32904
rect 43496 32892 43502 32904
rect 43806 32892 43812 32904
rect 43496 32864 43812 32892
rect 43496 32852 43502 32864
rect 43806 32852 43812 32864
rect 43864 32852 43870 32904
rect 44082 32892 44088 32904
rect 44043 32864 44088 32892
rect 44082 32852 44088 32864
rect 44140 32852 44146 32904
rect 50065 32895 50123 32901
rect 50065 32861 50077 32895
rect 50111 32892 50123 32895
rect 50154 32892 50160 32904
rect 50111 32864 50160 32892
rect 50111 32861 50123 32864
rect 50065 32855 50123 32861
rect 50154 32852 50160 32864
rect 50212 32852 50218 32904
rect 50264 32892 50292 32932
rect 50341 32929 50353 32963
rect 50387 32929 50399 32963
rect 50341 32923 50399 32929
rect 50525 32963 50583 32969
rect 50525 32929 50537 32963
rect 50571 32960 50583 32963
rect 51166 32960 51172 32972
rect 50571 32932 51172 32960
rect 50571 32929 50583 32932
rect 50525 32923 50583 32929
rect 51166 32920 51172 32932
rect 51224 32920 51230 32972
rect 55858 32920 55864 32972
rect 55916 32960 55922 32972
rect 61562 32960 61568 32972
rect 55916 32932 61568 32960
rect 55916 32920 55922 32932
rect 61562 32920 61568 32932
rect 61620 32920 61626 32972
rect 61838 32960 61844 32972
rect 61799 32932 61844 32960
rect 61838 32920 61844 32932
rect 61896 32920 61902 32972
rect 62022 32960 62028 32972
rect 61983 32932 62028 32960
rect 62022 32920 62028 32932
rect 62080 32920 62086 32972
rect 62390 32960 62396 32972
rect 62224 32932 62396 32960
rect 50982 32892 50988 32904
rect 50264 32864 50988 32892
rect 50982 32852 50988 32864
rect 51040 32852 51046 32904
rect 53374 32852 53380 32904
rect 53432 32892 53438 32904
rect 56686 32892 56692 32904
rect 53432 32864 56692 32892
rect 53432 32852 53438 32864
rect 56686 32852 56692 32864
rect 56744 32852 56750 32904
rect 62224 32892 62252 32932
rect 62390 32920 62396 32932
rect 62448 32960 62454 32972
rect 62485 32963 62543 32969
rect 62485 32960 62497 32963
rect 62448 32932 62497 32960
rect 62448 32920 62454 32932
rect 62485 32929 62497 32932
rect 62531 32929 62543 32963
rect 62485 32923 62543 32929
rect 62577 32963 62635 32969
rect 62577 32929 62589 32963
rect 62623 32960 62635 32963
rect 63034 32960 63040 32972
rect 62623 32932 63040 32960
rect 62623 32929 62635 32932
rect 62577 32923 62635 32929
rect 63034 32920 63040 32932
rect 63092 32960 63098 32972
rect 63313 32963 63371 32969
rect 63313 32960 63325 32963
rect 63092 32932 63325 32960
rect 63092 32920 63098 32932
rect 63313 32929 63325 32932
rect 63359 32929 63371 32963
rect 63696 32960 63724 33059
rect 67910 33056 67916 33108
rect 67968 33096 67974 33108
rect 68738 33096 68744 33108
rect 67968 33068 68744 33096
rect 67968 33056 67974 33068
rect 68738 33056 68744 33068
rect 68796 33056 68802 33108
rect 75546 33096 75552 33108
rect 75507 33068 75552 33096
rect 75546 33056 75552 33068
rect 75604 33056 75610 33108
rect 77754 33096 77760 33108
rect 77715 33068 77760 33096
rect 77754 33056 77760 33068
rect 77812 33056 77818 33108
rect 85206 33056 85212 33108
rect 85264 33096 85270 33108
rect 85301 33099 85359 33105
rect 85301 33096 85313 33099
rect 85264 33068 85313 33096
rect 85264 33056 85270 33068
rect 85301 33065 85313 33068
rect 85347 33065 85359 33099
rect 85301 33059 85359 33065
rect 66990 33028 66996 33040
rect 66951 33000 66996 33028
rect 66990 32988 66996 33000
rect 67048 32988 67054 33040
rect 68833 33031 68891 33037
rect 68833 33028 68845 33031
rect 67376 33000 68845 33028
rect 67376 32969 67404 33000
rect 68833 32997 68845 33000
rect 68879 33028 68891 33031
rect 69290 33028 69296 33040
rect 68879 33000 69296 33028
rect 68879 32997 68891 33000
rect 68833 32991 68891 32997
rect 69290 32988 69296 33000
rect 69348 32988 69354 33040
rect 76006 32988 76012 33040
rect 76064 33028 76070 33040
rect 82262 33028 82268 33040
rect 76064 33000 77984 33028
rect 76064 32988 76070 33000
rect 67361 32963 67419 32969
rect 67361 32960 67373 32963
rect 63696 32932 67373 32960
rect 63313 32923 63371 32929
rect 67361 32929 67373 32932
rect 67407 32929 67419 32963
rect 67361 32923 67419 32929
rect 67450 32920 67456 32972
rect 67508 32960 67514 32972
rect 67910 32960 67916 32972
rect 67508 32932 67553 32960
rect 67871 32932 67916 32960
rect 67508 32920 67514 32932
rect 67910 32920 67916 32932
rect 67968 32920 67974 32972
rect 68094 32960 68100 32972
rect 68055 32932 68100 32960
rect 68094 32920 68100 32932
rect 68152 32920 68158 32972
rect 73982 32960 73988 32972
rect 73943 32932 73988 32960
rect 73982 32920 73988 32932
rect 74040 32920 74046 32972
rect 74258 32960 74264 32972
rect 74219 32932 74264 32960
rect 74258 32920 74264 32932
rect 74316 32920 74322 32972
rect 74442 32960 74448 32972
rect 74403 32932 74448 32960
rect 74442 32920 74448 32932
rect 74500 32920 74506 32972
rect 75457 32963 75515 32969
rect 75457 32960 75469 32963
rect 74828 32932 75469 32960
rect 61672 32864 62252 32892
rect 68465 32895 68523 32901
rect 33597 32827 33655 32833
rect 33597 32824 33609 32827
rect 32508 32796 33609 32824
rect 33597 32793 33609 32796
rect 33643 32824 33655 32827
rect 37182 32824 37188 32836
rect 33643 32796 37188 32824
rect 33643 32793 33655 32796
rect 33597 32787 33655 32793
rect 37182 32784 37188 32796
rect 37240 32784 37246 32836
rect 42334 32824 42340 32836
rect 42295 32796 42340 32824
rect 42334 32784 42340 32796
rect 42392 32784 42398 32836
rect 61672 32833 61700 32864
rect 68465 32861 68477 32895
rect 68511 32892 68523 32895
rect 68830 32892 68836 32904
rect 68511 32864 68836 32892
rect 68511 32861 68523 32864
rect 68465 32855 68523 32861
rect 68830 32852 68836 32864
rect 68888 32852 68894 32904
rect 73433 32895 73491 32901
rect 73433 32861 73445 32895
rect 73479 32861 73491 32895
rect 73433 32855 73491 32861
rect 61657 32827 61715 32833
rect 61657 32824 61669 32827
rect 56520 32796 61669 32824
rect 29549 32759 29607 32765
rect 29549 32756 29561 32759
rect 24360 32728 29561 32756
rect 24360 32716 24366 32728
rect 29549 32725 29561 32728
rect 29595 32756 29607 32759
rect 31481 32759 31539 32765
rect 31481 32756 31493 32759
rect 29595 32728 31493 32756
rect 29595 32725 29607 32728
rect 29549 32719 29607 32725
rect 31481 32725 31493 32728
rect 31527 32756 31539 32759
rect 31573 32759 31631 32765
rect 31573 32756 31585 32759
rect 31527 32728 31585 32756
rect 31527 32725 31539 32728
rect 31481 32719 31539 32725
rect 31573 32725 31585 32728
rect 31619 32725 31631 32759
rect 31573 32719 31631 32725
rect 31846 32716 31852 32768
rect 31904 32756 31910 32768
rect 33321 32759 33379 32765
rect 33321 32756 33333 32759
rect 31904 32728 33333 32756
rect 31904 32716 31910 32728
rect 33321 32725 33333 32728
rect 33367 32725 33379 32759
rect 37918 32756 37924 32768
rect 37879 32728 37924 32756
rect 33321 32719 33379 32725
rect 37918 32716 37924 32728
rect 37976 32716 37982 32768
rect 38289 32759 38347 32765
rect 38289 32725 38301 32759
rect 38335 32756 38347 32759
rect 41782 32756 41788 32768
rect 38335 32728 41788 32756
rect 38335 32725 38347 32728
rect 38289 32719 38347 32725
rect 41782 32716 41788 32728
rect 41840 32716 41846 32768
rect 41966 32756 41972 32768
rect 41927 32728 41972 32756
rect 41966 32716 41972 32728
rect 42024 32716 42030 32768
rect 42426 32716 42432 32768
rect 42484 32756 42490 32768
rect 46385 32759 46443 32765
rect 46385 32756 46397 32759
rect 42484 32728 46397 32756
rect 42484 32716 42490 32728
rect 46385 32725 46397 32728
rect 46431 32756 46443 32759
rect 56520 32756 56548 32796
rect 61657 32793 61669 32796
rect 61703 32793 61715 32827
rect 73448 32824 73476 32855
rect 74258 32824 74264 32836
rect 73448 32796 74264 32824
rect 61657 32787 61715 32793
rect 74258 32784 74264 32796
rect 74316 32784 74322 32836
rect 46431 32728 56548 32756
rect 63037 32759 63095 32765
rect 46431 32725 46443 32728
rect 46385 32719 46443 32725
rect 63037 32725 63049 32759
rect 63083 32756 63095 32759
rect 63218 32756 63224 32768
rect 63083 32728 63224 32756
rect 63083 32725 63095 32728
rect 63037 32719 63095 32725
rect 63218 32716 63224 32728
rect 63276 32716 63282 32768
rect 63494 32756 63500 32768
rect 63455 32728 63500 32756
rect 63494 32716 63500 32728
rect 63552 32716 63558 32768
rect 66990 32716 66996 32768
rect 67048 32756 67054 32768
rect 68094 32756 68100 32768
rect 67048 32728 68100 32756
rect 67048 32716 67054 32728
rect 68094 32716 68100 32728
rect 68152 32716 68158 32768
rect 69934 32716 69940 32768
rect 69992 32756 69998 32768
rect 74828 32756 74856 32932
rect 75457 32929 75469 32932
rect 75503 32960 75515 32963
rect 75733 32963 75791 32969
rect 75733 32960 75745 32963
rect 75503 32932 75745 32960
rect 75503 32929 75515 32932
rect 75457 32923 75515 32929
rect 75733 32929 75745 32932
rect 75779 32960 75791 32963
rect 77386 32960 77392 32972
rect 75779 32932 77392 32960
rect 75779 32929 75791 32932
rect 75733 32923 75791 32929
rect 77386 32920 77392 32932
rect 77444 32920 77450 32972
rect 77956 32969 77984 33000
rect 80440 33000 82268 33028
rect 80440 32969 80468 33000
rect 82262 32988 82268 33000
rect 82320 32988 82326 33040
rect 82538 32988 82544 33040
rect 82596 33028 82602 33040
rect 82596 33000 83228 33028
rect 82596 32988 82602 33000
rect 77941 32963 77999 32969
rect 77941 32929 77953 32963
rect 77987 32929 77999 32963
rect 77941 32923 77999 32929
rect 80425 32963 80483 32969
rect 80425 32929 80437 32963
rect 80471 32929 80483 32963
rect 80425 32923 80483 32929
rect 80514 32920 80520 32972
rect 80572 32960 80578 32972
rect 81437 32963 81495 32969
rect 81437 32960 81449 32963
rect 80572 32932 81449 32960
rect 80572 32920 80578 32932
rect 81437 32929 81449 32932
rect 81483 32929 81495 32963
rect 81437 32923 81495 32929
rect 82173 32963 82231 32969
rect 82173 32929 82185 32963
rect 82219 32960 82231 32963
rect 82354 32960 82360 32972
rect 82219 32932 82360 32960
rect 82219 32929 82231 32932
rect 82173 32923 82231 32929
rect 82354 32920 82360 32932
rect 82412 32960 82418 32972
rect 83200 32969 83228 33000
rect 82633 32963 82691 32969
rect 82633 32960 82645 32963
rect 82412 32932 82645 32960
rect 82412 32920 82418 32932
rect 82633 32929 82645 32932
rect 82679 32929 82691 32963
rect 82633 32923 82691 32929
rect 83185 32963 83243 32969
rect 83185 32929 83197 32963
rect 83231 32929 83243 32963
rect 83185 32923 83243 32929
rect 82446 32852 82452 32904
rect 82504 32892 82510 32904
rect 83461 32895 83519 32901
rect 83461 32892 83473 32895
rect 82504 32864 83473 32892
rect 82504 32852 82510 32864
rect 83461 32861 83473 32864
rect 83507 32861 83519 32895
rect 83461 32855 83519 32861
rect 85022 32852 85028 32904
rect 85080 32892 85086 32904
rect 85316 32892 85344 33059
rect 88426 33056 88432 33108
rect 88484 33096 88490 33108
rect 88521 33099 88579 33105
rect 88521 33096 88533 33099
rect 88484 33068 88533 33096
rect 88484 33056 88490 33068
rect 88521 33065 88533 33068
rect 88567 33065 88579 33099
rect 88521 33059 88579 33065
rect 85666 33028 85672 33040
rect 85627 33000 85672 33028
rect 85666 32988 85672 33000
rect 85724 32988 85730 33040
rect 87230 33028 87236 33040
rect 86328 33000 87236 33028
rect 86328 32969 86356 33000
rect 87230 32988 87236 33000
rect 87288 33028 87294 33040
rect 88245 33031 88303 33037
rect 88245 33028 88257 33031
rect 87288 33000 88257 33028
rect 87288 32988 87294 33000
rect 88245 32997 88257 33000
rect 88291 32997 88303 33031
rect 88245 32991 88303 32997
rect 86313 32963 86371 32969
rect 86313 32929 86325 32963
rect 86359 32929 86371 32963
rect 86678 32960 86684 32972
rect 86591 32932 86684 32960
rect 86313 32923 86371 32929
rect 86678 32920 86684 32932
rect 86736 32920 86742 32972
rect 86770 32920 86776 32972
rect 86828 32960 86834 32972
rect 86828 32932 86873 32960
rect 86828 32920 86834 32932
rect 88334 32920 88340 32972
rect 88392 32960 88398 32972
rect 88429 32963 88487 32969
rect 88429 32960 88441 32963
rect 88392 32932 88441 32960
rect 88392 32920 88398 32932
rect 88429 32929 88441 32932
rect 88475 32960 88487 32963
rect 88889 32963 88947 32969
rect 88889 32960 88901 32963
rect 88475 32932 88901 32960
rect 88475 32929 88487 32932
rect 88429 32923 88487 32929
rect 88889 32929 88901 32932
rect 88935 32929 88947 32963
rect 88889 32923 88947 32929
rect 86221 32895 86279 32901
rect 86221 32892 86233 32895
rect 85080 32864 86233 32892
rect 85080 32852 85086 32864
rect 86221 32861 86233 32864
rect 86267 32861 86279 32895
rect 86221 32855 86279 32861
rect 75178 32784 75184 32836
rect 75236 32824 75242 32836
rect 81621 32827 81679 32833
rect 81621 32824 81633 32827
rect 75236 32796 81633 32824
rect 75236 32784 75242 32796
rect 81621 32793 81633 32796
rect 81667 32793 81679 32827
rect 81621 32787 81679 32793
rect 69992 32728 74856 32756
rect 81636 32756 81664 32787
rect 82078 32784 82084 32836
rect 82136 32824 82142 32836
rect 82725 32827 82783 32833
rect 82725 32824 82737 32827
rect 82136 32796 82737 32824
rect 82136 32784 82142 32796
rect 82725 32793 82737 32796
rect 82771 32793 82783 32827
rect 86696 32824 86724 32920
rect 82725 32787 82783 32793
rect 85592 32796 86724 32824
rect 85592 32768 85620 32796
rect 82357 32759 82415 32765
rect 82357 32756 82369 32759
rect 81636 32728 82369 32756
rect 69992 32716 69998 32728
rect 82357 32725 82369 32728
rect 82403 32756 82415 32759
rect 82538 32756 82544 32768
rect 82403 32728 82544 32756
rect 82403 32725 82415 32728
rect 82357 32719 82415 32725
rect 82538 32716 82544 32728
rect 82596 32716 82602 32768
rect 85574 32756 85580 32768
rect 85535 32728 85580 32756
rect 85574 32716 85580 32728
rect 85632 32716 85638 32768
rect 1104 32666 108008 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 65686 32666
rect 65738 32614 65750 32666
rect 65802 32614 65814 32666
rect 65866 32614 65878 32666
rect 65930 32614 96406 32666
rect 96458 32614 96470 32666
rect 96522 32614 96534 32666
rect 96586 32614 96598 32666
rect 96650 32614 108008 32666
rect 1104 32592 108008 32614
rect 3786 32512 3792 32564
rect 3844 32552 3850 32564
rect 3844 32524 9904 32552
rect 3844 32512 3850 32524
rect 6546 32444 6552 32496
rect 6604 32484 6610 32496
rect 9876 32484 9904 32524
rect 9950 32512 9956 32564
rect 10008 32552 10014 32564
rect 10413 32555 10471 32561
rect 10413 32552 10425 32555
rect 10008 32524 10425 32552
rect 10008 32512 10014 32524
rect 10413 32521 10425 32524
rect 10459 32552 10471 32555
rect 10778 32552 10784 32564
rect 10459 32524 10784 32552
rect 10459 32521 10471 32524
rect 10413 32515 10471 32521
rect 10778 32512 10784 32524
rect 10836 32512 10842 32564
rect 35437 32555 35495 32561
rect 10888 32524 33180 32552
rect 10888 32484 10916 32524
rect 15838 32484 15844 32496
rect 6604 32456 9812 32484
rect 9876 32456 10916 32484
rect 15799 32456 15844 32484
rect 6604 32444 6610 32456
rect 3142 32416 3148 32428
rect 3103 32388 3148 32416
rect 3142 32376 3148 32388
rect 3200 32376 3206 32428
rect 8478 32416 8484 32428
rect 8439 32388 8484 32416
rect 8478 32376 8484 32388
rect 8536 32376 8542 32428
rect 8849 32419 8907 32425
rect 8849 32385 8861 32419
rect 8895 32416 8907 32419
rect 9398 32416 9404 32428
rect 8895 32388 9404 32416
rect 8895 32385 8907 32388
rect 8849 32379 8907 32385
rect 2869 32351 2927 32357
rect 2869 32317 2881 32351
rect 2915 32348 2927 32351
rect 2958 32348 2964 32360
rect 2915 32320 2964 32348
rect 2915 32317 2927 32320
rect 2869 32311 2927 32317
rect 2958 32308 2964 32320
rect 3016 32308 3022 32360
rect 8018 32348 8024 32360
rect 7979 32320 8024 32348
rect 8018 32308 8024 32320
rect 8076 32308 8082 32360
rect 8389 32351 8447 32357
rect 8389 32317 8401 32351
rect 8435 32348 8447 32351
rect 8864 32348 8892 32379
rect 9398 32376 9404 32388
rect 9456 32376 9462 32428
rect 8435 32320 8892 32348
rect 9677 32351 9735 32357
rect 8435 32317 8447 32320
rect 8389 32311 8447 32317
rect 9677 32317 9689 32351
rect 9723 32317 9735 32351
rect 9677 32311 9735 32317
rect 8036 32280 8064 32308
rect 9692 32280 9720 32311
rect 8036 32252 9720 32280
rect 9784 32280 9812 32456
rect 15838 32444 15844 32456
rect 15896 32444 15902 32496
rect 16850 32484 16856 32496
rect 16811 32456 16856 32484
rect 16850 32444 16856 32456
rect 16908 32444 16914 32496
rect 18693 32487 18751 32493
rect 18693 32453 18705 32487
rect 18739 32484 18751 32487
rect 19610 32484 19616 32496
rect 18739 32456 19616 32484
rect 18739 32453 18751 32456
rect 18693 32447 18751 32453
rect 19610 32444 19616 32456
rect 19668 32444 19674 32496
rect 21358 32484 21364 32496
rect 20180 32456 21364 32484
rect 10042 32416 10048 32428
rect 10003 32388 10048 32416
rect 10042 32376 10048 32388
rect 10100 32376 10106 32428
rect 9950 32348 9956 32360
rect 9911 32320 9956 32348
rect 9950 32308 9956 32320
rect 10008 32308 10014 32360
rect 15654 32348 15660 32360
rect 15615 32320 15660 32348
rect 15654 32308 15660 32320
rect 15712 32308 15718 32360
rect 16761 32351 16819 32357
rect 16761 32317 16773 32351
rect 16807 32348 16819 32351
rect 18506 32348 18512 32360
rect 16807 32320 18512 32348
rect 16807 32317 16819 32320
rect 16761 32311 16819 32317
rect 18506 32308 18512 32320
rect 18564 32308 18570 32360
rect 18601 32351 18659 32357
rect 18601 32317 18613 32351
rect 18647 32317 18659 32351
rect 19978 32348 19984 32360
rect 19939 32320 19984 32348
rect 18601 32311 18659 32317
rect 16666 32280 16672 32292
rect 9784 32252 16672 32280
rect 16666 32240 16672 32252
rect 16724 32240 16730 32292
rect 17954 32240 17960 32292
rect 18012 32280 18018 32292
rect 18616 32280 18644 32311
rect 19978 32308 19984 32320
rect 20036 32308 20042 32360
rect 20073 32351 20131 32357
rect 20073 32317 20085 32351
rect 20119 32317 20131 32351
rect 20180 32348 20208 32456
rect 21358 32444 21364 32456
rect 21416 32444 21422 32496
rect 21542 32484 21548 32496
rect 21503 32456 21548 32484
rect 21542 32444 21548 32456
rect 21600 32444 21606 32496
rect 25590 32444 25596 32496
rect 25648 32484 25654 32496
rect 25648 32456 26464 32484
rect 25648 32444 25654 32456
rect 20533 32351 20591 32357
rect 20533 32348 20545 32351
rect 20180 32320 20545 32348
rect 20073 32311 20131 32317
rect 20533 32317 20545 32320
rect 20579 32317 20591 32351
rect 20533 32311 20591 32317
rect 20717 32351 20775 32357
rect 20717 32317 20729 32351
rect 20763 32348 20775 32351
rect 21560 32348 21588 32444
rect 24765 32419 24823 32425
rect 24765 32385 24777 32419
rect 24811 32416 24823 32419
rect 24949 32419 25007 32425
rect 24949 32416 24961 32419
rect 24811 32388 24961 32416
rect 24811 32385 24823 32388
rect 24765 32379 24823 32385
rect 24949 32385 24961 32388
rect 24995 32416 25007 32419
rect 25222 32416 25228 32428
rect 24995 32388 25228 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 25222 32376 25228 32388
rect 25280 32376 25286 32428
rect 26050 32416 26056 32428
rect 26011 32388 26056 32416
rect 26050 32376 26056 32388
rect 26108 32376 26114 32428
rect 26436 32425 26464 32456
rect 27154 32444 27160 32496
rect 27212 32484 27218 32496
rect 27249 32487 27307 32493
rect 27249 32484 27261 32487
rect 27212 32456 27261 32484
rect 27212 32444 27218 32456
rect 27249 32453 27261 32456
rect 27295 32453 27307 32487
rect 27249 32447 27307 32453
rect 29362 32444 29368 32496
rect 29420 32484 29426 32496
rect 31386 32484 31392 32496
rect 29420 32456 31392 32484
rect 29420 32444 29426 32456
rect 31386 32444 31392 32456
rect 31444 32444 31450 32496
rect 33152 32484 33180 32524
rect 35437 32521 35449 32555
rect 35483 32552 35495 32555
rect 36170 32552 36176 32564
rect 35483 32524 36176 32552
rect 35483 32521 35495 32524
rect 35437 32515 35495 32521
rect 36170 32512 36176 32524
rect 36228 32512 36234 32564
rect 37182 32512 37188 32564
rect 37240 32552 37246 32564
rect 37645 32555 37703 32561
rect 37645 32552 37657 32555
rect 37240 32524 37657 32552
rect 37240 32512 37246 32524
rect 37645 32521 37657 32524
rect 37691 32521 37703 32555
rect 37645 32515 37703 32521
rect 42153 32555 42211 32561
rect 42153 32521 42165 32555
rect 42199 32552 42211 32555
rect 44082 32552 44088 32564
rect 42199 32524 44088 32552
rect 42199 32521 42211 32524
rect 42153 32515 42211 32521
rect 44082 32512 44088 32524
rect 44140 32512 44146 32564
rect 53558 32512 53564 32564
rect 53616 32512 53622 32564
rect 53650 32512 53656 32564
rect 53708 32552 53714 32564
rect 54573 32555 54631 32561
rect 54573 32552 54585 32555
rect 53708 32524 54585 32552
rect 53708 32512 53714 32524
rect 54573 32521 54585 32524
rect 54619 32521 54631 32555
rect 54573 32515 54631 32521
rect 62298 32512 62304 32564
rect 62356 32552 62362 32564
rect 69934 32552 69940 32564
rect 62356 32524 69940 32552
rect 62356 32512 62362 32524
rect 69934 32512 69940 32524
rect 69992 32512 69998 32564
rect 86954 32552 86960 32564
rect 70044 32524 86960 32552
rect 40773 32487 40831 32493
rect 40773 32484 40785 32487
rect 33152 32456 40785 32484
rect 40773 32453 40785 32456
rect 40819 32484 40831 32487
rect 40819 32456 41000 32484
rect 40819 32453 40831 32456
rect 40773 32447 40831 32453
rect 26421 32419 26479 32425
rect 26421 32385 26433 32419
rect 26467 32416 26479 32419
rect 26605 32419 26663 32425
rect 26605 32416 26617 32419
rect 26467 32388 26617 32416
rect 26467 32385 26479 32388
rect 26421 32379 26479 32385
rect 26605 32385 26617 32388
rect 26651 32416 26663 32419
rect 29380 32416 29408 32444
rect 40972 32428 41000 32456
rect 41598 32444 41604 32496
rect 41656 32484 41662 32496
rect 42426 32484 42432 32496
rect 41656 32456 42432 32484
rect 41656 32444 41662 32456
rect 42426 32444 42432 32456
rect 42484 32444 42490 32496
rect 42978 32484 42984 32496
rect 42939 32456 42984 32484
rect 42978 32444 42984 32456
rect 43036 32444 43042 32496
rect 53576 32484 53604 32512
rect 54757 32487 54815 32493
rect 54757 32484 54769 32487
rect 53208 32456 54769 32484
rect 31570 32416 31576 32428
rect 26651 32388 29408 32416
rect 31531 32388 31576 32416
rect 26651 32385 26663 32388
rect 26605 32379 26663 32385
rect 31570 32376 31576 32388
rect 31628 32376 31634 32428
rect 31846 32416 31852 32428
rect 31807 32388 31852 32416
rect 31846 32376 31852 32388
rect 31904 32376 31910 32428
rect 34330 32376 34336 32428
rect 34388 32416 34394 32428
rect 37277 32419 37335 32425
rect 37277 32416 37289 32419
rect 34388 32388 37289 32416
rect 34388 32376 34394 32388
rect 37277 32385 37289 32388
rect 37323 32385 37335 32419
rect 40954 32416 40960 32428
rect 40867 32388 40960 32416
rect 37277 32379 37335 32385
rect 20763 32320 21588 32348
rect 25041 32351 25099 32357
rect 20763 32317 20775 32320
rect 20717 32311 20775 32317
rect 25041 32317 25053 32351
rect 25087 32348 25099 32351
rect 25590 32348 25596 32360
rect 25087 32320 25596 32348
rect 25087 32317 25099 32320
rect 25041 32311 25099 32317
rect 18012 32252 18644 32280
rect 20088 32280 20116 32311
rect 25590 32308 25596 32320
rect 25648 32308 25654 32360
rect 25777 32351 25835 32357
rect 25777 32317 25789 32351
rect 25823 32348 25835 32351
rect 26326 32348 26332 32360
rect 25823 32320 26332 32348
rect 25823 32317 25835 32320
rect 25777 32311 25835 32317
rect 26326 32308 26332 32320
rect 26384 32308 26390 32360
rect 27062 32348 27068 32360
rect 26896 32320 27068 32348
rect 21726 32280 21732 32292
rect 20088 32252 21732 32280
rect 18012 32240 18018 32252
rect 21726 32240 21732 32252
rect 21784 32240 21790 32292
rect 2866 32172 2872 32224
rect 2924 32212 2930 32224
rect 4249 32215 4307 32221
rect 4249 32212 4261 32215
rect 2924 32184 4261 32212
rect 2924 32172 2930 32184
rect 4249 32181 4261 32184
rect 4295 32181 4307 32215
rect 4706 32212 4712 32224
rect 4667 32184 4712 32212
rect 4249 32175 4307 32181
rect 4706 32172 4712 32184
rect 4764 32172 4770 32224
rect 20990 32212 20996 32224
rect 20951 32184 20996 32212
rect 20990 32172 20996 32184
rect 21048 32172 21054 32224
rect 22278 32172 22284 32224
rect 22336 32212 22342 32224
rect 26896 32221 26924 32320
rect 27062 32308 27068 32320
rect 27120 32308 27126 32360
rect 27154 32308 27160 32360
rect 27212 32348 27218 32360
rect 33226 32348 33232 32360
rect 27212 32320 33232 32348
rect 27212 32308 27218 32320
rect 33226 32308 33232 32320
rect 33284 32308 33290 32360
rect 35253 32351 35311 32357
rect 35253 32348 35265 32351
rect 35084 32320 35265 32348
rect 35084 32224 35112 32320
rect 35253 32317 35265 32320
rect 35299 32317 35311 32351
rect 35253 32311 35311 32317
rect 36170 32308 36176 32360
rect 36228 32348 36234 32360
rect 36357 32351 36415 32357
rect 36357 32348 36369 32351
rect 36228 32320 36369 32348
rect 36228 32308 36234 32320
rect 36357 32317 36369 32320
rect 36403 32317 36415 32351
rect 37292 32348 37320 32379
rect 40954 32376 40960 32388
rect 41012 32376 41018 32428
rect 53208 32425 53236 32456
rect 54757 32453 54769 32456
rect 54803 32453 54815 32487
rect 61654 32484 61660 32496
rect 61615 32456 61660 32484
rect 54757 32447 54815 32453
rect 61654 32444 61660 32456
rect 61712 32444 61718 32496
rect 69658 32484 69664 32496
rect 69619 32456 69664 32484
rect 69658 32444 69664 32456
rect 69716 32444 69722 32496
rect 53193 32419 53251 32425
rect 53193 32385 53205 32419
rect 53239 32385 53251 32419
rect 54294 32416 54300 32428
rect 54255 32388 54300 32416
rect 53193 32379 53251 32385
rect 54294 32376 54300 32388
rect 54352 32376 54358 32428
rect 54846 32376 54852 32428
rect 54904 32416 54910 32428
rect 57054 32416 57060 32428
rect 54904 32388 57060 32416
rect 54904 32376 54910 32388
rect 57054 32376 57060 32388
rect 57112 32376 57118 32428
rect 67082 32376 67088 32428
rect 67140 32416 67146 32428
rect 67450 32416 67456 32428
rect 67140 32388 67456 32416
rect 67140 32376 67146 32388
rect 67450 32376 67456 32388
rect 67508 32416 67514 32428
rect 67508 32388 68876 32416
rect 67508 32376 67514 32388
rect 37461 32351 37519 32357
rect 37461 32348 37473 32351
rect 37292 32320 37473 32348
rect 36357 32311 36415 32317
rect 37461 32317 37473 32320
rect 37507 32348 37519 32351
rect 37918 32348 37924 32360
rect 37507 32320 37924 32348
rect 37507 32317 37519 32320
rect 37461 32311 37519 32317
rect 37918 32308 37924 32320
rect 37976 32308 37982 32360
rect 41141 32351 41199 32357
rect 41141 32348 41153 32351
rect 40604 32320 41153 32348
rect 40604 32289 40632 32320
rect 41141 32317 41153 32320
rect 41187 32317 41199 32351
rect 41598 32348 41604 32360
rect 41559 32320 41604 32348
rect 41141 32311 41199 32317
rect 41598 32308 41604 32320
rect 41656 32308 41662 32360
rect 41693 32351 41751 32357
rect 41693 32317 41705 32351
rect 41739 32348 41751 32351
rect 42334 32348 42340 32360
rect 41739 32320 42340 32348
rect 41739 32317 41751 32320
rect 41693 32311 41751 32317
rect 42334 32308 42340 32320
rect 42392 32348 42398 32360
rect 42613 32351 42671 32357
rect 42613 32348 42625 32351
rect 42392 32320 42625 32348
rect 42392 32308 42398 32320
rect 42613 32317 42625 32320
rect 42659 32317 42671 32351
rect 42613 32311 42671 32317
rect 42978 32308 42984 32360
rect 43036 32348 43042 32360
rect 43165 32351 43223 32357
rect 43165 32348 43177 32351
rect 43036 32320 43177 32348
rect 43036 32308 43042 32320
rect 43165 32317 43177 32320
rect 43211 32317 43223 32351
rect 44358 32348 44364 32360
rect 44319 32320 44364 32348
rect 43165 32311 43223 32317
rect 44358 32308 44364 32320
rect 44416 32308 44422 32360
rect 48038 32308 48044 32360
rect 48096 32348 48102 32360
rect 48133 32351 48191 32357
rect 48133 32348 48145 32351
rect 48096 32320 48145 32348
rect 48096 32308 48102 32320
rect 48133 32317 48145 32320
rect 48179 32317 48191 32351
rect 48133 32311 48191 32317
rect 53285 32351 53343 32357
rect 53285 32317 53297 32351
rect 53331 32348 53343 32351
rect 53466 32348 53472 32360
rect 53331 32320 53472 32348
rect 53331 32317 53343 32320
rect 53285 32311 53343 32317
rect 53466 32308 53472 32320
rect 53524 32308 53530 32360
rect 53742 32348 53748 32360
rect 53703 32320 53748 32348
rect 53742 32308 53748 32320
rect 53800 32308 53806 32360
rect 53837 32351 53895 32357
rect 53837 32317 53849 32351
rect 53883 32348 53895 32351
rect 55030 32348 55036 32360
rect 53883 32320 55036 32348
rect 53883 32317 53895 32320
rect 53837 32311 53895 32317
rect 55030 32308 55036 32320
rect 55088 32308 55094 32360
rect 60553 32351 60611 32357
rect 60553 32348 60565 32351
rect 60384 32320 60565 32348
rect 40589 32283 40647 32289
rect 40589 32280 40601 32283
rect 36556 32252 40601 32280
rect 36556 32224 36584 32252
rect 40589 32249 40601 32252
rect 40635 32249 40647 32283
rect 40589 32243 40647 32249
rect 41230 32240 41236 32292
rect 41288 32280 41294 32292
rect 41288 32252 42104 32280
rect 41288 32240 41294 32252
rect 26881 32215 26939 32221
rect 26881 32212 26893 32215
rect 22336 32184 26893 32212
rect 22336 32172 22342 32184
rect 26881 32181 26893 32184
rect 26927 32181 26939 32215
rect 26881 32175 26939 32181
rect 31570 32172 31576 32224
rect 31628 32212 31634 32224
rect 33321 32215 33379 32221
rect 33321 32212 33333 32215
rect 31628 32184 33333 32212
rect 31628 32172 31634 32184
rect 33321 32181 33333 32184
rect 33367 32181 33379 32215
rect 35066 32212 35072 32224
rect 35027 32184 35072 32212
rect 33321 32175 33379 32181
rect 35066 32172 35072 32184
rect 35124 32172 35130 32224
rect 36538 32212 36544 32224
rect 36499 32184 36544 32212
rect 36538 32172 36544 32184
rect 36596 32172 36602 32224
rect 36630 32172 36636 32224
rect 36688 32212 36694 32224
rect 41966 32212 41972 32224
rect 36688 32184 41972 32212
rect 36688 32172 36694 32184
rect 41966 32172 41972 32184
rect 42024 32172 42030 32224
rect 42076 32212 42104 32252
rect 42702 32240 42708 32292
rect 42760 32280 42766 32292
rect 44453 32283 44511 32289
rect 44453 32280 44465 32283
rect 42760 32252 44465 32280
rect 42760 32240 42766 32252
rect 44453 32249 44465 32252
rect 44499 32280 44511 32283
rect 55858 32280 55864 32292
rect 44499 32252 55864 32280
rect 44499 32249 44511 32252
rect 44453 32243 44511 32249
rect 55858 32240 55864 32252
rect 55916 32240 55922 32292
rect 42794 32212 42800 32224
rect 42076 32184 42800 32212
rect 42794 32172 42800 32184
rect 42852 32212 42858 32224
rect 43349 32215 43407 32221
rect 43349 32212 43361 32215
rect 42852 32184 43361 32212
rect 42852 32172 42858 32184
rect 43349 32181 43361 32184
rect 43395 32212 43407 32215
rect 44542 32212 44548 32224
rect 43395 32184 44548 32212
rect 43395 32181 43407 32184
rect 43349 32175 43407 32181
rect 44542 32172 44548 32184
rect 44600 32172 44606 32224
rect 47949 32215 48007 32221
rect 47949 32181 47961 32215
rect 47995 32212 48007 32215
rect 48498 32212 48504 32224
rect 47995 32184 48504 32212
rect 47995 32181 48007 32184
rect 47949 32175 48007 32181
rect 48498 32172 48504 32184
rect 48556 32172 48562 32224
rect 55030 32212 55036 32224
rect 54991 32184 55036 32212
rect 55030 32172 55036 32184
rect 55088 32172 55094 32224
rect 60274 32172 60280 32224
rect 60332 32212 60338 32224
rect 60384 32221 60412 32320
rect 60553 32317 60565 32320
rect 60599 32317 60611 32351
rect 60553 32311 60611 32317
rect 60737 32351 60795 32357
rect 60737 32317 60749 32351
rect 60783 32317 60795 32351
rect 60737 32311 60795 32317
rect 61289 32351 61347 32357
rect 61289 32317 61301 32351
rect 61335 32317 61347 32351
rect 61289 32311 61347 32317
rect 61473 32351 61531 32357
rect 61473 32317 61485 32351
rect 61519 32348 61531 32351
rect 61838 32348 61844 32360
rect 61519 32320 61844 32348
rect 61519 32317 61531 32320
rect 61473 32311 61531 32317
rect 60369 32215 60427 32221
rect 60369 32212 60381 32215
rect 60332 32184 60381 32212
rect 60332 32172 60338 32184
rect 60369 32181 60381 32184
rect 60415 32181 60427 32215
rect 60752 32212 60780 32311
rect 61304 32280 61332 32311
rect 61838 32308 61844 32320
rect 61896 32348 61902 32360
rect 62117 32351 62175 32357
rect 62117 32348 62129 32351
rect 61896 32320 62129 32348
rect 61896 32308 61902 32320
rect 62117 32317 62129 32320
rect 62163 32348 62175 32351
rect 63494 32348 63500 32360
rect 62163 32320 63500 32348
rect 62163 32317 62175 32320
rect 62117 32311 62175 32317
rect 63494 32308 63500 32320
rect 63552 32308 63558 32360
rect 68557 32351 68615 32357
rect 68557 32348 68569 32351
rect 68296 32320 68569 32348
rect 62022 32280 62028 32292
rect 61304 32252 62028 32280
rect 62022 32240 62028 32252
rect 62080 32280 62086 32292
rect 62209 32283 62267 32289
rect 62209 32280 62221 32283
rect 62080 32252 62221 32280
rect 62080 32240 62086 32252
rect 62209 32249 62221 32252
rect 62255 32249 62267 32283
rect 62209 32243 62267 32249
rect 62114 32212 62120 32224
rect 60752 32184 62120 32212
rect 60369 32175 60427 32181
rect 62114 32172 62120 32184
rect 62172 32212 62178 32224
rect 62390 32212 62396 32224
rect 62172 32184 62396 32212
rect 62172 32172 62178 32184
rect 62390 32172 62396 32184
rect 62448 32172 62454 32224
rect 67542 32172 67548 32224
rect 67600 32212 67606 32224
rect 68296 32221 68324 32320
rect 68557 32317 68569 32320
rect 68603 32317 68615 32351
rect 68557 32311 68615 32317
rect 68741 32351 68799 32357
rect 68741 32317 68753 32351
rect 68787 32317 68799 32351
rect 68848 32348 68876 32388
rect 69201 32351 69259 32357
rect 69201 32348 69213 32351
rect 68848 32320 69213 32348
rect 68741 32311 68799 32317
rect 69201 32317 69213 32320
rect 69247 32317 69259 32351
rect 69201 32311 69259 32317
rect 68756 32280 68784 32311
rect 69290 32308 69296 32360
rect 69348 32348 69354 32360
rect 70044 32357 70072 32524
rect 86954 32512 86960 32524
rect 87012 32512 87018 32564
rect 76006 32444 76012 32496
rect 76064 32484 76070 32496
rect 85574 32484 85580 32496
rect 76064 32456 85580 32484
rect 76064 32444 76070 32456
rect 85574 32444 85580 32456
rect 85632 32444 85638 32496
rect 80514 32416 80520 32428
rect 72988 32388 80520 32416
rect 70029 32351 70087 32357
rect 70029 32348 70041 32351
rect 69348 32320 70041 32348
rect 69348 32308 69354 32320
rect 70029 32317 70041 32320
rect 70075 32317 70087 32351
rect 72988 32348 73016 32388
rect 80514 32376 80520 32388
rect 80572 32376 80578 32428
rect 81526 32416 81532 32428
rect 81487 32388 81532 32416
rect 81526 32376 81532 32388
rect 81584 32376 81590 32428
rect 82078 32416 82084 32428
rect 82039 32388 82084 32416
rect 82078 32376 82084 32388
rect 82136 32376 82142 32428
rect 82538 32416 82544 32428
rect 82499 32388 82544 32416
rect 82538 32376 82544 32388
rect 82596 32416 82602 32428
rect 82633 32419 82691 32425
rect 82633 32416 82645 32419
rect 82596 32388 82645 32416
rect 82596 32376 82602 32388
rect 82633 32385 82645 32388
rect 82679 32385 82691 32419
rect 82633 32379 82691 32385
rect 70029 32311 70087 32317
rect 70320 32320 73016 32348
rect 74169 32351 74227 32357
rect 70320 32280 70348 32320
rect 74169 32317 74181 32351
rect 74215 32317 74227 32351
rect 74169 32311 74227 32317
rect 68756 32252 70348 32280
rect 68281 32215 68339 32221
rect 68281 32212 68293 32215
rect 67600 32184 68293 32212
rect 67600 32172 67606 32184
rect 68281 32181 68293 32184
rect 68327 32181 68339 32215
rect 74184 32212 74212 32311
rect 74258 32308 74264 32360
rect 74316 32348 74322 32360
rect 74445 32351 74503 32357
rect 74445 32348 74457 32351
rect 74316 32320 74457 32348
rect 74316 32308 74322 32320
rect 74445 32317 74457 32320
rect 74491 32317 74503 32351
rect 74445 32311 74503 32317
rect 82357 32351 82415 32357
rect 82357 32317 82369 32351
rect 82403 32348 82415 32351
rect 82446 32348 82452 32360
rect 82403 32320 82452 32348
rect 82403 32317 82415 32320
rect 82357 32311 82415 32317
rect 82446 32308 82452 32320
rect 82504 32308 82510 32360
rect 75914 32280 75920 32292
rect 75380 32252 75920 32280
rect 75380 32212 75408 32252
rect 75914 32240 75920 32252
rect 75972 32240 75978 32292
rect 82464 32280 82492 32308
rect 82722 32280 82728 32292
rect 82464 32252 82728 32280
rect 82722 32240 82728 32252
rect 82780 32240 82786 32292
rect 75546 32212 75552 32224
rect 74184 32184 75408 32212
rect 75507 32184 75552 32212
rect 68281 32175 68339 32181
rect 75546 32172 75552 32184
rect 75604 32172 75610 32224
rect 80882 32172 80888 32224
rect 80940 32212 80946 32224
rect 85390 32212 85396 32224
rect 80940 32184 85396 32212
rect 80940 32172 80946 32184
rect 85390 32172 85396 32184
rect 85448 32172 85454 32224
rect 1104 32122 108008 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 50326 32122
rect 50378 32070 50390 32122
rect 50442 32070 50454 32122
rect 50506 32070 50518 32122
rect 50570 32070 81046 32122
rect 81098 32070 81110 32122
rect 81162 32070 81174 32122
rect 81226 32070 81238 32122
rect 81290 32070 108008 32122
rect 1104 32048 108008 32070
rect 10873 32011 10931 32017
rect 10873 31977 10885 32011
rect 10919 32008 10931 32011
rect 11698 32008 11704 32020
rect 10919 31980 11704 32008
rect 10919 31977 10931 31980
rect 10873 31971 10931 31977
rect 10980 31881 11008 31980
rect 11698 31968 11704 31980
rect 11756 31968 11762 32020
rect 32950 31968 32956 32020
rect 33008 32008 33014 32020
rect 34885 32011 34943 32017
rect 34885 32008 34897 32011
rect 33008 31980 34897 32008
rect 33008 31968 33014 31980
rect 34885 31977 34897 31980
rect 34931 32008 34943 32011
rect 36630 32008 36636 32020
rect 34931 31980 36636 32008
rect 34931 31977 34943 31980
rect 34885 31971 34943 31977
rect 36630 31968 36636 31980
rect 36688 31968 36694 32020
rect 40954 32008 40960 32020
rect 40915 31980 40960 32008
rect 40954 31968 40960 31980
rect 41012 31968 41018 32020
rect 42613 32011 42671 32017
rect 42613 31977 42625 32011
rect 42659 32008 42671 32011
rect 42702 32008 42708 32020
rect 42659 31980 42708 32008
rect 42659 31977 42671 31980
rect 42613 31971 42671 31977
rect 42702 31968 42708 31980
rect 42760 31968 42766 32020
rect 42794 31968 42800 32020
rect 42852 32008 42858 32020
rect 42852 31980 42897 32008
rect 42852 31968 42858 31980
rect 44358 31968 44364 32020
rect 44416 32008 44422 32020
rect 44729 32011 44787 32017
rect 44729 32008 44741 32011
rect 44416 31980 44741 32008
rect 44416 31968 44422 31980
rect 44729 31977 44741 31980
rect 44775 31977 44787 32011
rect 44729 31971 44787 31977
rect 52362 31968 52368 32020
rect 52420 32008 52426 32020
rect 53377 32011 53435 32017
rect 53377 32008 53389 32011
rect 52420 31980 53389 32008
rect 52420 31968 52426 31980
rect 53377 31977 53389 31980
rect 53423 32008 53435 32011
rect 53742 32008 53748 32020
rect 53423 31980 53748 32008
rect 53423 31977 53435 31980
rect 53377 31971 53435 31977
rect 53742 31968 53748 31980
rect 53800 31968 53806 32020
rect 54389 32011 54447 32017
rect 54389 31977 54401 32011
rect 54435 32008 54447 32011
rect 54846 32008 54852 32020
rect 54435 31980 54852 32008
rect 54435 31977 54447 31980
rect 54389 31971 54447 31977
rect 54846 31968 54852 31980
rect 54904 31968 54910 32020
rect 55030 31968 55036 32020
rect 55088 32008 55094 32020
rect 62298 32008 62304 32020
rect 55088 31980 62304 32008
rect 55088 31968 55094 31980
rect 62298 31968 62304 31980
rect 62356 31968 62362 32020
rect 62390 31968 62396 32020
rect 62448 32008 62454 32020
rect 68741 32011 68799 32017
rect 68741 32008 68753 32011
rect 62448 31980 68753 32008
rect 62448 31968 62454 31980
rect 16114 31900 16120 31952
rect 16172 31940 16178 31952
rect 16172 31912 17632 31940
rect 16172 31900 16178 31912
rect 10965 31875 11023 31881
rect 10965 31841 10977 31875
rect 11011 31841 11023 31875
rect 10965 31835 11023 31841
rect 16485 31875 16543 31881
rect 16485 31841 16497 31875
rect 16531 31872 16543 31875
rect 17034 31872 17040 31884
rect 16531 31844 17040 31872
rect 16531 31841 16543 31844
rect 16485 31835 16543 31841
rect 17034 31832 17040 31844
rect 17092 31832 17098 31884
rect 17221 31875 17279 31881
rect 17221 31841 17233 31875
rect 17267 31841 17279 31875
rect 17402 31872 17408 31884
rect 17363 31844 17408 31872
rect 17221 31835 17279 31841
rect 11238 31804 11244 31816
rect 11199 31776 11244 31804
rect 11238 31764 11244 31776
rect 11296 31764 11302 31816
rect 15378 31764 15384 31816
rect 15436 31804 15442 31816
rect 16209 31807 16267 31813
rect 16209 31804 16221 31807
rect 15436 31776 16221 31804
rect 15436 31764 15442 31776
rect 16209 31773 16221 31776
rect 16255 31804 16267 31807
rect 16574 31804 16580 31816
rect 16255 31776 16289 31804
rect 16535 31776 16580 31804
rect 16255 31773 16267 31776
rect 16209 31767 16267 31773
rect 12434 31696 12440 31748
rect 12492 31736 12498 31748
rect 16224 31736 16252 31767
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 17236 31804 17264 31835
rect 17402 31832 17408 31844
rect 17460 31832 17466 31884
rect 16776 31776 17264 31804
rect 17604 31804 17632 31912
rect 41506 31900 41512 31952
rect 41564 31940 41570 31952
rect 42337 31943 42395 31949
rect 41564 31912 42012 31940
rect 41564 31900 41570 31912
rect 17865 31875 17923 31881
rect 17865 31841 17877 31875
rect 17911 31872 17923 31875
rect 19521 31875 19579 31881
rect 17911 31844 18276 31872
rect 17911 31841 17923 31844
rect 17865 31835 17923 31841
rect 17954 31804 17960 31816
rect 17604 31776 17960 31804
rect 16776 31736 16804 31776
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18248 31748 18276 31844
rect 19521 31841 19533 31875
rect 19567 31872 19579 31875
rect 19978 31872 19984 31884
rect 19567 31844 19984 31872
rect 19567 31841 19579 31844
rect 19521 31835 19579 31841
rect 19978 31832 19984 31844
rect 20036 31832 20042 31884
rect 34701 31875 34759 31881
rect 34701 31872 34713 31875
rect 34532 31844 34713 31872
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31804 19487 31807
rect 25406 31804 25412 31816
rect 19475 31776 25412 31804
rect 19475 31773 19487 31776
rect 19429 31767 19487 31773
rect 25406 31764 25412 31776
rect 25464 31764 25470 31816
rect 27062 31764 27068 31816
rect 27120 31804 27126 31816
rect 34532 31813 34560 31844
rect 34701 31841 34713 31844
rect 34747 31872 34759 31875
rect 35066 31872 35072 31884
rect 34747 31844 35072 31872
rect 34747 31841 34759 31844
rect 34701 31835 34759 31841
rect 35066 31832 35072 31844
rect 35124 31832 35130 31884
rect 41230 31832 41236 31884
rect 41288 31872 41294 31884
rect 41874 31881 41880 31884
rect 41873 31872 41880 31881
rect 41288 31844 41333 31872
rect 41835 31844 41880 31872
rect 41288 31832 41294 31844
rect 41873 31835 41880 31844
rect 41874 31832 41880 31835
rect 41932 31832 41938 31884
rect 41984 31881 42012 31912
rect 42337 31909 42349 31943
rect 42383 31909 42395 31943
rect 42337 31903 42395 31909
rect 41969 31875 42027 31881
rect 41969 31841 41981 31875
rect 42015 31872 42027 31875
rect 42352 31872 42380 31903
rect 44542 31900 44548 31952
rect 44600 31940 44606 31952
rect 56226 31940 56232 31952
rect 44600 31912 56232 31940
rect 44600 31900 44606 31912
rect 56226 31900 56232 31912
rect 56284 31900 56290 31952
rect 67542 31940 67548 31952
rect 66916 31912 67548 31940
rect 43625 31875 43683 31881
rect 43625 31872 43637 31875
rect 42015 31844 42288 31872
rect 42352 31844 43637 31872
rect 42015 31841 42027 31844
rect 41969 31835 42027 31841
rect 34517 31807 34575 31813
rect 34517 31804 34529 31807
rect 27120 31776 34529 31804
rect 27120 31764 27126 31776
rect 34517 31773 34529 31776
rect 34563 31773 34575 31807
rect 34517 31767 34575 31773
rect 40954 31764 40960 31816
rect 41012 31804 41018 31816
rect 41049 31807 41107 31813
rect 41049 31804 41061 31807
rect 41012 31776 41061 31804
rect 41012 31764 41018 31776
rect 41049 31773 41061 31776
rect 41095 31773 41107 31807
rect 41049 31767 41107 31773
rect 18230 31736 18236 31748
rect 12492 31708 16160 31736
rect 16224 31708 16804 31736
rect 18143 31708 18236 31736
rect 12492 31696 12498 31708
rect 12529 31671 12587 31677
rect 12529 31637 12541 31671
rect 12575 31668 12587 31671
rect 12986 31668 12992 31680
rect 12575 31640 12992 31668
rect 12575 31637 12587 31640
rect 12529 31631 12587 31637
rect 12986 31628 12992 31640
rect 13044 31628 13050 31680
rect 16132 31668 16160 31708
rect 18230 31696 18236 31708
rect 18288 31736 18294 31748
rect 18288 31708 19840 31736
rect 18288 31696 18294 31708
rect 17402 31668 17408 31680
rect 16132 31640 17408 31668
rect 17402 31628 17408 31640
rect 17460 31628 17466 31680
rect 19426 31628 19432 31680
rect 19484 31668 19490 31680
rect 19705 31671 19763 31677
rect 19705 31668 19717 31671
rect 19484 31640 19717 31668
rect 19484 31628 19490 31640
rect 19705 31637 19717 31640
rect 19751 31637 19763 31671
rect 19812 31668 19840 31708
rect 21358 31696 21364 31748
rect 21416 31736 21422 31748
rect 34790 31736 34796 31748
rect 21416 31708 34796 31736
rect 21416 31696 21422 31708
rect 34790 31696 34796 31708
rect 34848 31696 34854 31748
rect 40773 31739 40831 31745
rect 40773 31705 40785 31739
rect 40819 31736 40831 31739
rect 41874 31736 41880 31748
rect 40819 31708 41880 31736
rect 40819 31705 40831 31708
rect 40773 31699 40831 31705
rect 41874 31696 41880 31708
rect 41932 31696 41938 31748
rect 42260 31736 42288 31844
rect 43625 31841 43637 31844
rect 43671 31841 43683 31875
rect 43625 31835 43683 31841
rect 53190 31832 53196 31884
rect 53248 31872 53254 31884
rect 53285 31875 53343 31881
rect 53285 31872 53297 31875
rect 53248 31844 53297 31872
rect 53248 31832 53254 31844
rect 53285 31841 53297 31844
rect 53331 31872 53343 31875
rect 53374 31872 53380 31884
rect 53331 31844 53380 31872
rect 53331 31841 53343 31844
rect 53285 31835 53343 31841
rect 53374 31832 53380 31844
rect 53432 31832 53438 31884
rect 54389 31875 54447 31881
rect 54389 31872 54401 31875
rect 53484 31844 54401 31872
rect 42702 31804 42708 31816
rect 42444 31776 42708 31804
rect 42444 31736 42472 31776
rect 42702 31764 42708 31776
rect 42760 31764 42766 31816
rect 43346 31804 43352 31816
rect 43307 31776 43352 31804
rect 43346 31764 43352 31776
rect 43404 31764 43410 31816
rect 48314 31764 48320 31816
rect 48372 31804 48378 31816
rect 53484 31804 53512 31844
rect 54389 31841 54401 31844
rect 54435 31872 54447 31875
rect 54573 31875 54631 31881
rect 54573 31872 54585 31875
rect 54435 31844 54585 31872
rect 54435 31841 54447 31844
rect 54389 31835 54447 31841
rect 54573 31841 54585 31844
rect 54619 31841 54631 31875
rect 54573 31835 54631 31841
rect 54772 31844 55076 31872
rect 48372 31776 53512 31804
rect 48372 31764 48378 31776
rect 53650 31764 53656 31816
rect 53708 31804 53714 31816
rect 54772 31804 54800 31844
rect 53708 31776 54800 31804
rect 53708 31764 53714 31776
rect 54938 31736 54944 31748
rect 42260 31708 42472 31736
rect 46216 31708 54944 31736
rect 46216 31668 46244 31708
rect 54938 31696 54944 31708
rect 54996 31696 55002 31748
rect 55048 31736 55076 31844
rect 66916 31816 66944 31912
rect 67542 31900 67548 31912
rect 67600 31940 67606 31952
rect 67600 31912 67956 31940
rect 67600 31900 67606 31912
rect 67174 31832 67180 31884
rect 67232 31872 67238 31884
rect 67928 31881 67956 31912
rect 68020 31881 68048 31980
rect 68741 31977 68753 31980
rect 68787 31977 68799 32011
rect 74442 32008 74448 32020
rect 74403 31980 74448 32008
rect 68741 31971 68799 31977
rect 68756 31940 68784 31971
rect 74442 31968 74448 31980
rect 74500 31968 74506 32020
rect 76006 32008 76012 32020
rect 75967 31980 76012 32008
rect 76006 31968 76012 31980
rect 76064 31968 76070 32020
rect 76285 32011 76343 32017
rect 76285 31977 76297 32011
rect 76331 32008 76343 32011
rect 80882 32008 80888 32020
rect 76331 31980 80888 32008
rect 76331 31977 76343 31980
rect 76285 31971 76343 31977
rect 75178 31940 75184 31952
rect 68756 31912 75184 31940
rect 75178 31900 75184 31912
rect 75236 31900 75242 31952
rect 67453 31875 67511 31881
rect 67453 31872 67465 31875
rect 67232 31844 67465 31872
rect 67232 31832 67238 31844
rect 67453 31841 67465 31844
rect 67499 31841 67511 31875
rect 67453 31835 67511 31841
rect 67913 31875 67971 31881
rect 67913 31841 67925 31875
rect 67959 31841 67971 31875
rect 67913 31835 67971 31841
rect 68005 31875 68063 31881
rect 68005 31841 68017 31875
rect 68051 31841 68063 31875
rect 68005 31835 68063 31841
rect 69014 31832 69020 31884
rect 69072 31872 69078 31884
rect 74353 31875 74411 31881
rect 74353 31872 74365 31875
rect 69072 31844 74365 31872
rect 69072 31832 69078 31844
rect 74353 31841 74365 31844
rect 74399 31872 74411 31875
rect 74629 31875 74687 31881
rect 74629 31872 74641 31875
rect 74399 31844 74641 31872
rect 74399 31841 74411 31844
rect 74353 31835 74411 31841
rect 74629 31841 74641 31844
rect 74675 31872 74687 31875
rect 75546 31872 75552 31884
rect 74675 31844 75552 31872
rect 74675 31841 74687 31844
rect 74629 31835 74687 31841
rect 75546 31832 75552 31844
rect 75604 31832 75610 31884
rect 75730 31832 75736 31884
rect 75788 31872 75794 31884
rect 75825 31875 75883 31881
rect 75825 31872 75837 31875
rect 75788 31844 75837 31872
rect 75788 31832 75794 31844
rect 75825 31841 75837 31844
rect 75871 31872 75883 31875
rect 76300 31872 76328 31971
rect 80882 31968 80888 31980
rect 80940 31968 80946 32020
rect 81161 32011 81219 32017
rect 81161 31977 81173 32011
rect 81207 32008 81219 32011
rect 81434 32008 81440 32020
rect 81207 31980 81440 32008
rect 81207 31977 81219 31980
rect 81161 31971 81219 31977
rect 81434 31968 81440 31980
rect 81492 31968 81498 32020
rect 88429 32011 88487 32017
rect 88429 31977 88441 32011
rect 88475 31977 88487 32011
rect 88429 31971 88487 31977
rect 82262 31940 82268 31952
rect 80808 31912 82268 31940
rect 75871 31844 76328 31872
rect 75871 31841 75883 31844
rect 75825 31835 75883 31841
rect 78674 31832 78680 31884
rect 78732 31872 78738 31884
rect 79778 31872 79784 31884
rect 78732 31844 79784 31872
rect 78732 31832 78738 31844
rect 79778 31832 79784 31844
rect 79836 31872 79842 31884
rect 80517 31875 80575 31881
rect 80517 31872 80529 31875
rect 79836 31844 80529 31872
rect 79836 31832 79842 31844
rect 80517 31841 80529 31844
rect 80563 31841 80575 31875
rect 80517 31835 80575 31841
rect 80664 31875 80722 31881
rect 80664 31841 80676 31875
rect 80710 31872 80722 31875
rect 80808 31872 80836 31912
rect 82262 31900 82268 31912
rect 82320 31900 82326 31952
rect 87417 31943 87475 31949
rect 87417 31940 87429 31943
rect 86972 31912 87429 31940
rect 86972 31884 87000 31912
rect 87417 31909 87429 31912
rect 87463 31940 87475 31943
rect 88444 31940 88472 31971
rect 87463 31912 88472 31940
rect 87463 31909 87475 31912
rect 87417 31903 87475 31909
rect 81345 31875 81403 31881
rect 81345 31872 81357 31875
rect 80710 31844 80836 31872
rect 80900 31844 81357 31872
rect 80710 31841 80722 31844
rect 80664 31835 80722 31841
rect 80900 31816 80928 31844
rect 81345 31841 81357 31844
rect 81391 31841 81403 31875
rect 85390 31872 85396 31884
rect 85351 31844 85396 31872
rect 81345 31835 81403 31841
rect 85390 31832 85396 31844
rect 85448 31832 85454 31884
rect 86773 31875 86831 31881
rect 86773 31872 86785 31875
rect 85500 31844 86785 31872
rect 66898 31804 66904 31816
rect 66859 31776 66904 31804
rect 66898 31764 66904 31776
rect 66956 31764 66962 31816
rect 67266 31804 67272 31816
rect 67227 31776 67272 31804
rect 67266 31764 67272 31776
rect 67324 31764 67330 31816
rect 80882 31804 80888 31816
rect 80795 31776 80888 31804
rect 80882 31764 80888 31776
rect 80940 31764 80946 31816
rect 82814 31764 82820 31816
rect 82872 31804 82878 31816
rect 85500 31813 85528 31844
rect 86773 31841 86785 31844
rect 86819 31841 86831 31875
rect 86954 31872 86960 31884
rect 86915 31844 86960 31872
rect 86773 31835 86831 31841
rect 86954 31832 86960 31844
rect 87012 31832 87018 31884
rect 87325 31875 87383 31881
rect 87325 31841 87337 31875
rect 87371 31872 87383 31875
rect 87690 31872 87696 31884
rect 87371 31844 87696 31872
rect 87371 31841 87383 31844
rect 87325 31835 87383 31841
rect 87690 31832 87696 31844
rect 87748 31832 87754 31884
rect 88242 31872 88248 31884
rect 88203 31844 88248 31872
rect 88242 31832 88248 31844
rect 88300 31832 88306 31884
rect 85485 31807 85543 31813
rect 85485 31804 85497 31807
rect 82872 31776 85497 31804
rect 82872 31764 82878 31776
rect 85485 31773 85497 31776
rect 85531 31773 85543 31807
rect 85485 31767 85543 31773
rect 55048 31708 80928 31736
rect 19812 31640 46244 31668
rect 19705 31631 19763 31637
rect 50154 31628 50160 31680
rect 50212 31668 50218 31680
rect 53101 31671 53159 31677
rect 53101 31668 53113 31671
rect 50212 31640 53113 31668
rect 50212 31628 50218 31640
rect 53101 31637 53113 31640
rect 53147 31668 53159 31671
rect 53190 31668 53196 31680
rect 53147 31640 53196 31668
rect 53147 31637 53159 31640
rect 53101 31631 53159 31637
rect 53190 31628 53196 31640
rect 53248 31628 53254 31680
rect 54110 31628 54116 31680
rect 54168 31668 54174 31680
rect 54665 31671 54723 31677
rect 54665 31668 54677 31671
rect 54168 31640 54677 31668
rect 54168 31628 54174 31640
rect 54665 31637 54677 31640
rect 54711 31637 54723 31671
rect 54665 31631 54723 31637
rect 55398 31628 55404 31680
rect 55456 31668 55462 31680
rect 67085 31671 67143 31677
rect 67085 31668 67097 31671
rect 55456 31640 67097 31668
rect 55456 31628 55462 31640
rect 67085 31637 67097 31640
rect 67131 31668 67143 31671
rect 67266 31668 67272 31680
rect 67131 31640 67272 31668
rect 67131 31637 67143 31640
rect 67085 31631 67143 31637
rect 67266 31628 67272 31640
rect 67324 31668 67330 31680
rect 67542 31668 67548 31680
rect 67324 31640 67548 31668
rect 67324 31628 67330 31640
rect 67542 31628 67548 31640
rect 67600 31628 67606 31680
rect 68462 31668 68468 31680
rect 68423 31640 68468 31668
rect 68462 31628 68468 31640
rect 68520 31628 68526 31680
rect 69014 31668 69020 31680
rect 68975 31640 69020 31668
rect 69014 31628 69020 31640
rect 69072 31628 69078 31680
rect 80514 31628 80520 31680
rect 80572 31668 80578 31680
rect 80793 31671 80851 31677
rect 80793 31668 80805 31671
rect 80572 31640 80805 31668
rect 80572 31628 80578 31640
rect 80793 31637 80805 31640
rect 80839 31637 80851 31671
rect 80900 31668 80928 31708
rect 85114 31668 85120 31680
rect 80900 31640 85120 31668
rect 80793 31631 80851 31637
rect 85114 31628 85120 31640
rect 85172 31628 85178 31680
rect 1104 31578 108008 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 65686 31578
rect 65738 31526 65750 31578
rect 65802 31526 65814 31578
rect 65866 31526 65878 31578
rect 65930 31526 96406 31578
rect 96458 31526 96470 31578
rect 96522 31526 96534 31578
rect 96586 31526 96598 31578
rect 96650 31526 108008 31578
rect 1104 31504 108008 31526
rect 12069 31467 12127 31473
rect 12069 31433 12081 31467
rect 12115 31464 12127 31467
rect 12161 31467 12219 31473
rect 12161 31464 12173 31467
rect 12115 31436 12173 31464
rect 12115 31433 12127 31436
rect 12069 31427 12127 31433
rect 12161 31433 12173 31436
rect 12207 31464 12219 31467
rect 17494 31464 17500 31476
rect 12207 31436 17500 31464
rect 12207 31433 12219 31436
rect 12161 31427 12219 31433
rect 17494 31424 17500 31436
rect 17552 31424 17558 31476
rect 17954 31424 17960 31476
rect 18012 31464 18018 31476
rect 57149 31467 57207 31473
rect 18012 31436 55536 31464
rect 18012 31424 18018 31436
rect 4062 31356 4068 31408
rect 4120 31396 4126 31408
rect 23658 31396 23664 31408
rect 4120 31368 23664 31396
rect 4120 31356 4126 31368
rect 23658 31356 23664 31368
rect 23716 31356 23722 31408
rect 23753 31399 23811 31405
rect 23753 31365 23765 31399
rect 23799 31396 23811 31399
rect 25498 31396 25504 31408
rect 23799 31368 25504 31396
rect 23799 31365 23811 31368
rect 23753 31359 23811 31365
rect 3145 31331 3203 31337
rect 3145 31297 3157 31331
rect 3191 31328 3203 31331
rect 7006 31328 7012 31340
rect 3191 31300 7012 31328
rect 3191 31297 3203 31300
rect 3145 31291 3203 31297
rect 7006 31288 7012 31300
rect 7064 31288 7070 31340
rect 16114 31328 16120 31340
rect 16075 31300 16120 31328
rect 16114 31288 16120 31300
rect 16172 31288 16178 31340
rect 16390 31288 16396 31340
rect 16448 31328 16454 31340
rect 22738 31328 22744 31340
rect 16448 31300 22744 31328
rect 16448 31288 16454 31300
rect 22738 31288 22744 31300
rect 22796 31288 22802 31340
rect 24780 31337 24808 31368
rect 25498 31356 25504 31368
rect 25556 31356 25562 31408
rect 35250 31396 35256 31408
rect 35211 31368 35256 31396
rect 35250 31356 35256 31368
rect 35308 31356 35314 31408
rect 35529 31399 35587 31405
rect 35529 31365 35541 31399
rect 35575 31365 35587 31399
rect 41966 31396 41972 31408
rect 41927 31368 41972 31396
rect 35529 31359 35587 31365
rect 24765 31331 24823 31337
rect 24765 31297 24777 31331
rect 24811 31297 24823 31331
rect 24765 31291 24823 31297
rect 25406 31288 25412 31340
rect 25464 31328 25470 31340
rect 35158 31328 35164 31340
rect 25464 31300 35164 31328
rect 25464 31288 25470 31300
rect 35158 31288 35164 31300
rect 35216 31288 35222 31340
rect 2869 31263 2927 31269
rect 2869 31229 2881 31263
rect 2915 31260 2927 31263
rect 2958 31260 2964 31272
rect 2915 31232 2964 31260
rect 2915 31229 2927 31232
rect 2869 31223 2927 31229
rect 2958 31220 2964 31232
rect 3016 31260 3022 31272
rect 4706 31260 4712 31272
rect 3016 31232 4712 31260
rect 3016 31220 3022 31232
rect 4706 31220 4712 31232
rect 4764 31220 4770 31272
rect 11885 31263 11943 31269
rect 11885 31229 11897 31263
rect 11931 31260 11943 31263
rect 12161 31263 12219 31269
rect 12161 31260 12173 31263
rect 11931 31232 12173 31260
rect 11931 31229 11943 31232
rect 11885 31223 11943 31229
rect 12161 31229 12173 31232
rect 12207 31229 12219 31263
rect 12161 31223 12219 31229
rect 15654 31220 15660 31272
rect 15712 31260 15718 31272
rect 15749 31263 15807 31269
rect 15749 31260 15761 31263
rect 15712 31232 15761 31260
rect 15712 31220 15718 31232
rect 15749 31229 15761 31232
rect 15795 31229 15807 31263
rect 15749 31223 15807 31229
rect 17678 31220 17684 31272
rect 17736 31220 17742 31272
rect 18322 31220 18328 31272
rect 18380 31260 18386 31272
rect 23753 31263 23811 31269
rect 23753 31260 23765 31263
rect 18380 31232 23765 31260
rect 18380 31220 18386 31232
rect 23753 31229 23765 31232
rect 23799 31260 23811 31263
rect 23845 31263 23903 31269
rect 23845 31260 23857 31263
rect 23799 31232 23857 31260
rect 23799 31229 23811 31232
rect 23753 31223 23811 31229
rect 23845 31229 23857 31232
rect 23891 31229 23903 31263
rect 24670 31260 24676 31272
rect 24631 31232 24676 31260
rect 23845 31223 23903 31229
rect 24670 31220 24676 31232
rect 24728 31220 24734 31272
rect 24946 31220 24952 31272
rect 25004 31260 25010 31272
rect 25042 31263 25100 31269
rect 25042 31260 25054 31263
rect 25004 31232 25054 31260
rect 25004 31220 25010 31232
rect 25042 31229 25054 31232
rect 25088 31229 25100 31263
rect 25042 31223 25100 31229
rect 25133 31263 25191 31269
rect 25133 31229 25145 31263
rect 25179 31229 25191 31263
rect 25133 31223 25191 31229
rect 29273 31263 29331 31269
rect 29273 31229 29285 31263
rect 29319 31260 29331 31263
rect 29454 31260 29460 31272
rect 29319 31232 29460 31260
rect 29319 31229 29331 31232
rect 29273 31223 29331 31229
rect 15562 31192 15568 31204
rect 15523 31164 15568 31192
rect 15562 31152 15568 31164
rect 15620 31192 15626 31204
rect 16482 31192 16488 31204
rect 15620 31164 16488 31192
rect 15620 31152 15626 31164
rect 16482 31152 16488 31164
rect 16540 31152 16546 31204
rect 17034 31152 17040 31204
rect 17092 31192 17098 31204
rect 17696 31192 17724 31220
rect 22738 31192 22744 31204
rect 17092 31164 22744 31192
rect 17092 31152 17098 31164
rect 22738 31152 22744 31164
rect 22796 31152 22802 31204
rect 24026 31192 24032 31204
rect 23987 31164 24032 31192
rect 24026 31152 24032 31164
rect 24084 31152 24090 31204
rect 3510 31084 3516 31136
rect 3568 31124 3574 31136
rect 4249 31127 4307 31133
rect 4249 31124 4261 31127
rect 3568 31096 4261 31124
rect 3568 31084 3574 31096
rect 4249 31093 4261 31096
rect 4295 31093 4307 31127
rect 4706 31124 4712 31136
rect 4667 31096 4712 31124
rect 4249 31087 4307 31093
rect 4706 31084 4712 31096
rect 4764 31084 4770 31136
rect 9582 31084 9588 31136
rect 9640 31124 9646 31136
rect 11701 31127 11759 31133
rect 11701 31124 11713 31127
rect 9640 31096 11713 31124
rect 9640 31084 9646 31096
rect 11701 31093 11713 31096
rect 11747 31093 11759 31127
rect 11701 31087 11759 31093
rect 12894 31084 12900 31136
rect 12952 31124 12958 31136
rect 18322 31124 18328 31136
rect 12952 31096 18328 31124
rect 12952 31084 12958 31096
rect 18322 31084 18328 31096
rect 18380 31084 18386 31136
rect 24946 31084 24952 31136
rect 25004 31124 25010 31136
rect 25148 31124 25176 31223
rect 29454 31220 29460 31232
rect 29512 31220 29518 31272
rect 35268 31260 35296 31356
rect 35544 31328 35572 31359
rect 41966 31356 41972 31368
rect 42024 31356 42030 31408
rect 55398 31396 55404 31408
rect 42168 31368 55404 31396
rect 35618 31328 35624 31340
rect 35531 31300 35624 31328
rect 35618 31288 35624 31300
rect 35676 31328 35682 31340
rect 41230 31328 41236 31340
rect 35676 31300 41236 31328
rect 35676 31288 35682 31300
rect 41230 31288 41236 31300
rect 41288 31328 41294 31340
rect 41782 31328 41788 31340
rect 41288 31300 41788 31328
rect 41288 31288 41294 31300
rect 41782 31288 41788 31300
rect 41840 31288 41846 31340
rect 35345 31263 35403 31269
rect 35345 31260 35357 31263
rect 35268 31232 35357 31260
rect 35345 31229 35357 31232
rect 35391 31229 35403 31263
rect 35345 31223 35403 31229
rect 35894 31220 35900 31272
rect 35952 31260 35958 31272
rect 36449 31263 36507 31269
rect 36449 31260 36461 31263
rect 35952 31232 36461 31260
rect 35952 31220 35958 31232
rect 36449 31229 36461 31232
rect 36495 31229 36507 31263
rect 36722 31260 36728 31272
rect 36683 31232 36728 31260
rect 36449 31223 36507 31229
rect 36722 31220 36728 31232
rect 36780 31220 36786 31272
rect 40770 31260 40776 31272
rect 37384 31232 40776 31260
rect 25406 31152 25412 31204
rect 25464 31192 25470 31204
rect 25464 31164 32444 31192
rect 25464 31152 25470 31164
rect 25004 31096 25176 31124
rect 25004 31084 25010 31096
rect 28994 31084 29000 31136
rect 29052 31124 29058 31136
rect 29365 31127 29423 31133
rect 29365 31124 29377 31127
rect 29052 31096 29377 31124
rect 29052 31084 29058 31096
rect 29365 31093 29377 31096
rect 29411 31093 29423 31127
rect 29365 31087 29423 31093
rect 29454 31084 29460 31136
rect 29512 31124 29518 31136
rect 29641 31127 29699 31133
rect 29641 31124 29653 31127
rect 29512 31096 29653 31124
rect 29512 31084 29518 31096
rect 29641 31093 29653 31096
rect 29687 31124 29699 31127
rect 30650 31124 30656 31136
rect 29687 31096 30656 31124
rect 29687 31093 29699 31096
rect 29641 31087 29699 31093
rect 30650 31084 30656 31096
rect 30708 31084 30714 31136
rect 32416 31124 32444 31164
rect 37384 31124 37412 31232
rect 40770 31220 40776 31232
rect 40828 31220 40834 31272
rect 41984 31260 42012 31356
rect 42061 31263 42119 31269
rect 42061 31260 42073 31263
rect 41984 31232 42073 31260
rect 42061 31229 42073 31232
rect 42107 31229 42119 31263
rect 42061 31223 42119 31229
rect 38102 31192 38108 31204
rect 38063 31164 38108 31192
rect 38102 31152 38108 31164
rect 38160 31152 38166 31204
rect 42168 31192 42196 31368
rect 55398 31356 55404 31368
rect 55456 31356 55462 31408
rect 55508 31396 55536 31436
rect 57149 31433 57161 31467
rect 57195 31464 57207 31467
rect 61930 31464 61936 31476
rect 57195 31436 61936 31464
rect 57195 31433 57207 31436
rect 57149 31427 57207 31433
rect 61930 31424 61936 31436
rect 61988 31424 61994 31476
rect 62114 31464 62120 31476
rect 62075 31436 62120 31464
rect 62114 31424 62120 31436
rect 62172 31424 62178 31476
rect 63218 31464 63224 31476
rect 63179 31436 63224 31464
rect 63218 31424 63224 31436
rect 63276 31424 63282 31476
rect 63586 31464 63592 31476
rect 63547 31436 63592 31464
rect 63586 31424 63592 31436
rect 63644 31424 63650 31476
rect 68462 31424 68468 31476
rect 68520 31464 68526 31476
rect 68695 31467 68753 31473
rect 68695 31464 68707 31467
rect 68520 31436 68707 31464
rect 68520 31424 68526 31436
rect 68695 31433 68707 31436
rect 68741 31433 68753 31467
rect 68830 31464 68836 31476
rect 68791 31436 68836 31464
rect 68695 31427 68753 31433
rect 68830 31424 68836 31436
rect 68888 31424 68894 31476
rect 75730 31464 75736 31476
rect 75691 31436 75736 31464
rect 75730 31424 75736 31436
rect 75788 31424 75794 31476
rect 75917 31467 75975 31473
rect 75917 31433 75929 31467
rect 75963 31464 75975 31467
rect 76006 31464 76012 31476
rect 75963 31436 76012 31464
rect 75963 31433 75975 31436
rect 75917 31427 75975 31433
rect 66898 31396 66904 31408
rect 55508 31368 66904 31396
rect 66898 31356 66904 31368
rect 66956 31356 66962 31408
rect 68370 31356 68376 31408
rect 68428 31396 68434 31408
rect 69017 31399 69075 31405
rect 69017 31396 69029 31399
rect 68428 31368 69029 31396
rect 68428 31356 68434 31368
rect 69017 31365 69029 31368
rect 69063 31365 69075 31399
rect 69017 31359 69075 31365
rect 73614 31356 73620 31408
rect 73672 31396 73678 31408
rect 75748 31396 75776 31424
rect 73672 31368 74212 31396
rect 73672 31356 73678 31368
rect 43254 31288 43260 31340
rect 43312 31328 43318 31340
rect 46569 31331 46627 31337
rect 46569 31328 46581 31331
rect 43312 31300 46581 31328
rect 43312 31288 43318 31300
rect 46569 31297 46581 31300
rect 46615 31328 46627 31331
rect 46753 31331 46811 31337
rect 46753 31328 46765 31331
rect 46615 31300 46765 31328
rect 46615 31297 46627 31300
rect 46569 31291 46627 31297
rect 46753 31297 46765 31300
rect 46799 31328 46811 31331
rect 46799 31300 47348 31328
rect 46799 31297 46811 31300
rect 46753 31291 46811 31297
rect 47320 31269 47348 31300
rect 54938 31288 54944 31340
rect 54996 31328 55002 31340
rect 74184 31337 74212 31368
rect 74368 31368 75776 31396
rect 57149 31331 57207 31337
rect 57149 31328 57161 31331
rect 54996 31300 57161 31328
rect 54996 31288 55002 31300
rect 57149 31297 57161 31300
rect 57195 31297 57207 31331
rect 57149 31291 57207 31297
rect 61933 31331 61991 31337
rect 61933 31297 61945 31331
rect 61979 31328 61991 31331
rect 63092 31331 63150 31337
rect 63092 31328 63104 31331
rect 61979 31300 63104 31328
rect 61979 31297 61991 31300
rect 61933 31291 61991 31297
rect 63092 31297 63104 31300
rect 63138 31297 63150 31331
rect 63092 31291 63150 31297
rect 63313 31331 63371 31337
rect 63313 31297 63325 31331
rect 63359 31297 63371 31331
rect 63313 31291 63371 31297
rect 68925 31331 68983 31337
rect 68925 31297 68937 31331
rect 68971 31328 68983 31331
rect 74169 31331 74227 31337
rect 68971 31300 74028 31328
rect 68971 31297 68983 31300
rect 68925 31291 68983 31297
rect 43165 31263 43223 31269
rect 43165 31229 43177 31263
rect 43211 31260 43223 31263
rect 47121 31263 47179 31269
rect 47121 31260 47133 31263
rect 43211 31232 43576 31260
rect 43211 31229 43223 31232
rect 43165 31223 43223 31229
rect 41984 31164 42196 31192
rect 32416 31096 37412 31124
rect 37918 31084 37924 31136
rect 37976 31124 37982 31136
rect 41984 31124 42012 31164
rect 37976 31096 42012 31124
rect 37976 31084 37982 31096
rect 42058 31084 42064 31136
rect 42116 31124 42122 31136
rect 42245 31127 42303 31133
rect 42245 31124 42257 31127
rect 42116 31096 42257 31124
rect 42116 31084 42122 31096
rect 42245 31093 42257 31096
rect 42291 31093 42303 31127
rect 42245 31087 42303 31093
rect 42426 31084 42432 31136
rect 42484 31124 42490 31136
rect 43548 31133 43576 31232
rect 46952 31232 47133 31260
rect 46952 31136 46980 31232
rect 47121 31229 47133 31232
rect 47167 31229 47179 31263
rect 47121 31223 47179 31229
rect 47305 31263 47363 31269
rect 47305 31229 47317 31263
rect 47351 31260 47363 31263
rect 47857 31263 47915 31269
rect 47857 31260 47869 31263
rect 47351 31232 47869 31260
rect 47351 31229 47363 31232
rect 47305 31223 47363 31229
rect 47857 31229 47869 31232
rect 47903 31229 47915 31263
rect 47857 31223 47915 31229
rect 48041 31263 48099 31269
rect 48041 31229 48053 31263
rect 48087 31260 48099 31263
rect 52362 31260 52368 31272
rect 48087 31232 52368 31260
rect 48087 31229 48099 31232
rect 48041 31223 48099 31229
rect 52362 31220 52368 31232
rect 52420 31220 52426 31272
rect 53650 31260 53656 31272
rect 53563 31232 53656 31260
rect 53650 31220 53656 31232
rect 53708 31220 53714 31272
rect 53745 31263 53803 31269
rect 53745 31229 53757 31263
rect 53791 31260 53803 31263
rect 53834 31260 53840 31272
rect 53791 31232 53840 31260
rect 53791 31229 53803 31232
rect 53745 31223 53803 31229
rect 53834 31220 53840 31232
rect 53892 31220 53898 31272
rect 54110 31260 54116 31272
rect 54071 31232 54116 31260
rect 54110 31220 54116 31232
rect 54168 31220 54174 31272
rect 54205 31263 54263 31269
rect 54205 31229 54217 31263
rect 54251 31260 54263 31263
rect 55030 31260 55036 31272
rect 54251 31232 55036 31260
rect 54251 31229 54263 31232
rect 54205 31223 54263 31229
rect 55030 31220 55036 31232
rect 55088 31260 55094 31272
rect 55125 31263 55183 31269
rect 55125 31260 55137 31263
rect 55088 31232 55137 31260
rect 55088 31220 55094 31232
rect 55125 31229 55137 31232
rect 55171 31229 55183 31263
rect 55125 31223 55183 31229
rect 58989 31263 59047 31269
rect 58989 31229 59001 31263
rect 59035 31260 59047 31263
rect 59262 31260 59268 31272
rect 59035 31232 59268 31260
rect 59035 31229 59047 31232
rect 58989 31223 59047 31229
rect 59262 31220 59268 31232
rect 59320 31220 59326 31272
rect 60458 31220 60464 31272
rect 60516 31260 60522 31272
rect 60645 31263 60703 31269
rect 60645 31260 60657 31263
rect 60516 31232 60657 31260
rect 60516 31220 60522 31232
rect 60645 31229 60657 31232
rect 60691 31229 60703 31263
rect 60826 31260 60832 31272
rect 60787 31232 60832 31260
rect 60645 31223 60703 31229
rect 60826 31220 60832 31232
rect 60884 31220 60890 31272
rect 61289 31263 61347 31269
rect 61289 31229 61301 31263
rect 61335 31229 61347 31263
rect 61289 31223 61347 31229
rect 61381 31263 61439 31269
rect 61381 31229 61393 31263
rect 61427 31260 61439 31263
rect 62114 31260 62120 31272
rect 61427 31232 62120 31260
rect 61427 31229 61439 31232
rect 61381 31223 61439 31229
rect 48409 31195 48467 31201
rect 48409 31161 48421 31195
rect 48455 31192 48467 31195
rect 49234 31192 49240 31204
rect 48455 31164 49240 31192
rect 48455 31161 48467 31164
rect 48409 31155 48467 31161
rect 49234 31152 49240 31164
rect 49292 31152 49298 31204
rect 53668 31192 53696 31220
rect 54941 31195 54999 31201
rect 54941 31192 54953 31195
rect 53668 31164 54953 31192
rect 54941 31161 54953 31164
rect 54987 31161 54999 31195
rect 54941 31155 54999 31161
rect 57330 31152 57336 31204
rect 57388 31192 57394 31204
rect 60274 31192 60280 31204
rect 57388 31164 60280 31192
rect 57388 31152 57394 31164
rect 60274 31152 60280 31164
rect 60332 31192 60338 31204
rect 61304 31192 61332 31223
rect 62114 31220 62120 31232
rect 62172 31220 62178 31272
rect 63328 31260 63356 31291
rect 63328 31232 68692 31260
rect 60332 31164 61332 31192
rect 60332 31152 60338 31164
rect 61930 31152 61936 31204
rect 61988 31192 61994 31204
rect 62206 31192 62212 31204
rect 61988 31164 62212 31192
rect 61988 31152 61994 31164
rect 62206 31152 62212 31164
rect 62264 31152 62270 31204
rect 62390 31152 62396 31204
rect 62448 31192 62454 31204
rect 62945 31195 63003 31201
rect 62945 31192 62957 31195
rect 62448 31164 62957 31192
rect 62448 31152 62454 31164
rect 62945 31161 62957 31164
rect 62991 31161 63003 31195
rect 62945 31155 63003 31161
rect 67450 31152 67456 31204
rect 67508 31192 67514 31204
rect 68557 31195 68615 31201
rect 68557 31192 68569 31195
rect 67508 31164 68569 31192
rect 67508 31152 67514 31164
rect 68557 31161 68569 31164
rect 68603 31161 68615 31195
rect 68664 31192 68692 31232
rect 72510 31192 72516 31204
rect 68664 31164 72516 31192
rect 68557 31155 68615 31161
rect 72510 31152 72516 31164
rect 72568 31152 72574 31204
rect 43257 31127 43315 31133
rect 43257 31124 43269 31127
rect 42484 31096 43269 31124
rect 42484 31084 42490 31096
rect 43257 31093 43269 31096
rect 43303 31093 43315 31127
rect 43257 31087 43315 31093
rect 43533 31127 43591 31133
rect 43533 31093 43545 31127
rect 43579 31124 43591 31127
rect 45002 31124 45008 31136
rect 43579 31096 45008 31124
rect 43579 31093 43591 31096
rect 43533 31087 43591 31093
rect 45002 31084 45008 31096
rect 45060 31084 45066 31136
rect 46934 31124 46940 31136
rect 46895 31096 46940 31124
rect 46934 31084 46940 31096
rect 46992 31084 46998 31136
rect 53282 31084 53288 31136
rect 53340 31124 53346 31136
rect 54665 31127 54723 31133
rect 54665 31124 54677 31127
rect 53340 31096 54677 31124
rect 53340 31084 53346 31096
rect 54665 31093 54677 31096
rect 54711 31093 54723 31127
rect 54665 31087 54723 31093
rect 58434 31084 58440 31136
rect 58492 31124 58498 31136
rect 59081 31127 59139 31133
rect 59081 31124 59093 31127
rect 58492 31096 59093 31124
rect 58492 31084 58498 31096
rect 59081 31093 59093 31096
rect 59127 31093 59139 31127
rect 60458 31124 60464 31136
rect 60419 31096 60464 31124
rect 59081 31087 59139 31093
rect 60458 31084 60464 31096
rect 60516 31084 60522 31136
rect 60826 31084 60832 31136
rect 60884 31124 60890 31136
rect 62022 31124 62028 31136
rect 60884 31096 62028 31124
rect 60884 31084 60890 31096
rect 62022 31084 62028 31096
rect 62080 31124 62086 31136
rect 62301 31127 62359 31133
rect 62301 31124 62313 31127
rect 62080 31096 62313 31124
rect 62080 31084 62086 31096
rect 62301 31093 62313 31096
rect 62347 31124 62359 31127
rect 67174 31124 67180 31136
rect 62347 31096 67180 31124
rect 62347 31093 62359 31096
rect 62301 31087 62359 31093
rect 67174 31084 67180 31096
rect 67232 31124 67238 31136
rect 69014 31124 69020 31136
rect 67232 31096 69020 31124
rect 67232 31084 67238 31096
rect 69014 31084 69020 31096
rect 69072 31084 69078 31136
rect 73614 31084 73620 31136
rect 73672 31124 73678 31136
rect 73709 31127 73767 31133
rect 73709 31124 73721 31127
rect 73672 31096 73721 31124
rect 73672 31084 73678 31096
rect 73709 31093 73721 31096
rect 73755 31124 73767 31127
rect 73893 31127 73951 31133
rect 73893 31124 73905 31127
rect 73755 31096 73905 31124
rect 73755 31093 73767 31096
rect 73709 31087 73767 31093
rect 73893 31093 73905 31096
rect 73939 31093 73951 31127
rect 74000 31124 74028 31300
rect 74169 31297 74181 31331
rect 74215 31297 74227 31331
rect 74169 31291 74227 31297
rect 74184 31192 74212 31291
rect 74368 31269 74396 31368
rect 74353 31263 74411 31269
rect 74353 31229 74365 31263
rect 74399 31229 74411 31263
rect 74353 31223 74411 31229
rect 74813 31263 74871 31269
rect 74813 31229 74825 31263
rect 74859 31229 74871 31263
rect 74813 31223 74871 31229
rect 74905 31263 74963 31269
rect 74905 31229 74917 31263
rect 74951 31260 74963 31263
rect 75932 31260 75960 31427
rect 76006 31424 76012 31436
rect 76064 31424 76070 31476
rect 79594 31424 79600 31476
rect 79652 31464 79658 31476
rect 79652 31436 84056 31464
rect 79652 31424 79658 31436
rect 82722 31356 82728 31408
rect 82780 31396 82786 31408
rect 84028 31396 84056 31436
rect 84194 31424 84200 31476
rect 84252 31464 84258 31476
rect 85114 31464 85120 31476
rect 84252 31436 84297 31464
rect 85075 31436 85120 31464
rect 84252 31424 84258 31436
rect 85114 31424 85120 31436
rect 85172 31464 85178 31476
rect 85172 31436 85804 31464
rect 85172 31424 85178 31436
rect 85022 31396 85028 31408
rect 82780 31368 83964 31396
rect 84028 31368 85028 31396
rect 82780 31356 82786 31368
rect 82188 31300 83872 31328
rect 79778 31260 79784 31272
rect 74951 31232 75960 31260
rect 79739 31232 79784 31260
rect 74951 31229 74963 31232
rect 74905 31223 74963 31229
rect 74828 31192 74856 31223
rect 79778 31220 79784 31232
rect 79836 31220 79842 31272
rect 79870 31220 79876 31272
rect 79928 31260 79934 31272
rect 79965 31263 80023 31269
rect 79965 31260 79977 31263
rect 79928 31232 79977 31260
rect 79928 31220 79934 31232
rect 79965 31229 79977 31232
rect 80011 31260 80023 31263
rect 80425 31263 80483 31269
rect 80425 31260 80437 31263
rect 80011 31232 80437 31260
rect 80011 31229 80023 31232
rect 79965 31223 80023 31229
rect 80425 31229 80437 31232
rect 80471 31229 80483 31263
rect 80425 31223 80483 31229
rect 82188 31201 82216 31300
rect 82354 31260 82360 31272
rect 82315 31232 82360 31260
rect 82354 31220 82360 31232
rect 82412 31220 82418 31272
rect 82722 31260 82728 31272
rect 82683 31232 82728 31260
rect 82722 31220 82728 31232
rect 82780 31220 82786 31272
rect 83645 31263 83703 31269
rect 83645 31229 83657 31263
rect 83691 31260 83703 31263
rect 83737 31263 83795 31269
rect 83737 31260 83749 31263
rect 83691 31232 83749 31260
rect 83691 31229 83703 31232
rect 83645 31223 83703 31229
rect 83737 31229 83749 31232
rect 83783 31229 83795 31263
rect 83737 31223 83795 31229
rect 74184 31164 74856 31192
rect 80333 31195 80391 31201
rect 80333 31161 80345 31195
rect 80379 31192 80391 31195
rect 82173 31195 82231 31201
rect 82173 31192 82185 31195
rect 80379 31164 82185 31192
rect 80379 31161 80391 31164
rect 80333 31155 80391 31161
rect 82173 31161 82185 31164
rect 82219 31161 82231 31195
rect 82173 31155 82231 31161
rect 75365 31127 75423 31133
rect 75365 31124 75377 31127
rect 74000 31096 75377 31124
rect 73893 31087 73951 31093
rect 75365 31093 75377 31096
rect 75411 31093 75423 31127
rect 83752 31124 83780 31223
rect 83844 31192 83872 31300
rect 83936 31269 83964 31368
rect 85022 31356 85028 31368
rect 85080 31356 85086 31408
rect 85485 31399 85543 31405
rect 85485 31365 85497 31399
rect 85531 31365 85543 31399
rect 85485 31359 85543 31365
rect 85500 31328 85528 31359
rect 84028 31300 85528 31328
rect 84028 31269 84056 31300
rect 83921 31263 83979 31269
rect 83921 31229 83933 31263
rect 83967 31229 83979 31263
rect 83921 31223 83979 31229
rect 84013 31263 84071 31269
rect 84013 31229 84025 31263
rect 84059 31229 84071 31263
rect 84013 31223 84071 31229
rect 85669 31263 85727 31269
rect 85669 31229 85681 31263
rect 85715 31229 85727 31263
rect 85776 31260 85804 31436
rect 85945 31263 86003 31269
rect 85945 31260 85957 31263
rect 85776 31232 85957 31260
rect 85669 31223 85727 31229
rect 85945 31229 85957 31232
rect 85991 31229 86003 31263
rect 87414 31260 87420 31272
rect 87375 31232 87420 31260
rect 85945 31223 86003 31229
rect 85390 31192 85396 31204
rect 83844 31164 85396 31192
rect 85390 31152 85396 31164
rect 85448 31152 85454 31204
rect 85684 31192 85712 31223
rect 87414 31220 87420 31232
rect 87472 31220 87478 31272
rect 87690 31260 87696 31272
rect 87651 31232 87696 31260
rect 87690 31220 87696 31232
rect 87748 31220 87754 31272
rect 86678 31192 86684 31204
rect 85684 31164 86684 31192
rect 86678 31152 86684 31164
rect 86736 31192 86742 31204
rect 87601 31195 87659 31201
rect 87601 31192 87613 31195
rect 86736 31164 87613 31192
rect 86736 31152 86742 31164
rect 87601 31161 87613 31164
rect 87647 31161 87659 31195
rect 87601 31155 87659 31161
rect 88153 31195 88211 31201
rect 88153 31161 88165 31195
rect 88199 31192 88211 31195
rect 88610 31192 88616 31204
rect 88199 31164 88616 31192
rect 88199 31161 88211 31164
rect 88153 31155 88211 31161
rect 88610 31152 88616 31164
rect 88668 31152 88674 31204
rect 87233 31127 87291 31133
rect 87233 31124 87245 31127
rect 83752 31096 87245 31124
rect 75365 31087 75423 31093
rect 87233 31093 87245 31096
rect 87279 31124 87291 31127
rect 87414 31124 87420 31136
rect 87279 31096 87420 31124
rect 87279 31093 87291 31096
rect 87233 31087 87291 31093
rect 87414 31084 87420 31096
rect 87472 31084 87478 31136
rect 1104 31034 108008 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 50326 31034
rect 50378 30982 50390 31034
rect 50442 30982 50454 31034
rect 50506 30982 50518 31034
rect 50570 30982 81046 31034
rect 81098 30982 81110 31034
rect 81162 30982 81174 31034
rect 81226 30982 81238 31034
rect 81290 30982 108008 31034
rect 1104 30960 108008 30982
rect 12894 30920 12900 30932
rect 11716 30892 12900 30920
rect 11149 30855 11207 30861
rect 11149 30821 11161 30855
rect 11195 30852 11207 30855
rect 11238 30852 11244 30864
rect 11195 30824 11244 30852
rect 11195 30821 11207 30824
rect 11149 30815 11207 30821
rect 11238 30812 11244 30824
rect 11296 30812 11302 30864
rect 5169 30787 5227 30793
rect 5169 30753 5181 30787
rect 5215 30784 5227 30787
rect 7742 30784 7748 30796
rect 5215 30756 7748 30784
rect 5215 30753 5227 30756
rect 5169 30747 5227 30753
rect 7742 30744 7748 30756
rect 7800 30744 7806 30796
rect 11716 30793 11744 30892
rect 12894 30880 12900 30892
rect 12952 30880 12958 30932
rect 12986 30880 12992 30932
rect 13044 30920 13050 30932
rect 17954 30920 17960 30932
rect 13044 30892 17960 30920
rect 13044 30880 13050 30892
rect 17954 30880 17960 30892
rect 18012 30880 18018 30932
rect 18230 30920 18236 30932
rect 18191 30892 18236 30920
rect 18230 30880 18236 30892
rect 18288 30880 18294 30932
rect 25225 30923 25283 30929
rect 25225 30889 25237 30923
rect 25271 30920 25283 30923
rect 25314 30920 25320 30932
rect 25271 30892 25320 30920
rect 25271 30889 25283 30892
rect 25225 30883 25283 30889
rect 25314 30880 25320 30892
rect 25372 30880 25378 30932
rect 30929 30923 30987 30929
rect 30929 30889 30941 30923
rect 30975 30920 30987 30923
rect 31018 30920 31024 30932
rect 30975 30892 31024 30920
rect 30975 30889 30987 30892
rect 30929 30883 30987 30889
rect 31018 30880 31024 30892
rect 31076 30920 31082 30932
rect 31570 30920 31576 30932
rect 31076 30892 31576 30920
rect 31076 30880 31082 30892
rect 31570 30880 31576 30892
rect 31628 30880 31634 30932
rect 35158 30880 35164 30932
rect 35216 30920 35222 30932
rect 36909 30923 36967 30929
rect 35216 30892 36860 30920
rect 35216 30880 35222 30892
rect 12342 30852 12348 30864
rect 12084 30824 12348 30852
rect 11057 30787 11115 30793
rect 11057 30753 11069 30787
rect 11103 30784 11115 30787
rect 11701 30787 11759 30793
rect 11701 30784 11713 30787
rect 11103 30756 11713 30784
rect 11103 30753 11115 30756
rect 11057 30747 11115 30753
rect 11701 30753 11713 30756
rect 11747 30753 11759 30787
rect 11701 30747 11759 30753
rect 11790 30744 11796 30796
rect 11848 30784 11854 30796
rect 12084 30793 12112 30824
rect 12342 30812 12348 30824
rect 12400 30852 12406 30864
rect 12434 30852 12440 30864
rect 12400 30824 12440 30852
rect 12400 30812 12406 30824
rect 12434 30812 12440 30824
rect 12492 30812 12498 30864
rect 12526 30812 12532 30864
rect 12584 30852 12590 30864
rect 13004 30852 13032 30880
rect 12584 30824 13032 30852
rect 12584 30812 12590 30824
rect 34790 30812 34796 30864
rect 34848 30852 34854 30864
rect 35253 30855 35311 30861
rect 35253 30852 35265 30855
rect 34848 30824 35265 30852
rect 34848 30812 34854 30824
rect 35253 30821 35265 30824
rect 35299 30852 35311 30855
rect 36722 30852 36728 30864
rect 35299 30824 36584 30852
rect 36683 30824 36728 30852
rect 35299 30821 35311 30824
rect 35253 30815 35311 30821
rect 12069 30787 12127 30793
rect 11848 30756 11893 30784
rect 11848 30744 11854 30756
rect 12069 30753 12081 30787
rect 12115 30753 12127 30787
rect 12618 30784 12624 30796
rect 12531 30756 12624 30784
rect 12069 30747 12127 30753
rect 4706 30676 4712 30728
rect 4764 30716 4770 30728
rect 4893 30719 4951 30725
rect 4893 30716 4905 30719
rect 4764 30688 4905 30716
rect 4764 30676 4770 30688
rect 4893 30685 4905 30688
rect 4939 30716 4951 30719
rect 4939 30688 6684 30716
rect 4939 30685 4951 30688
rect 4893 30679 4951 30685
rect 6656 30592 6684 30688
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 12084 30716 12112 30747
rect 12618 30744 12624 30756
rect 12676 30784 12682 30796
rect 16114 30784 16120 30796
rect 12676 30756 16120 30784
rect 12676 30744 12682 30756
rect 16114 30744 16120 30756
rect 16172 30744 16178 30796
rect 16574 30744 16580 30796
rect 16632 30784 16638 30796
rect 16945 30787 17003 30793
rect 16945 30784 16957 30787
rect 16632 30756 16957 30784
rect 16632 30744 16638 30756
rect 16945 30753 16957 30756
rect 16991 30753 17003 30787
rect 16945 30747 17003 30753
rect 19429 30787 19487 30793
rect 19429 30753 19441 30787
rect 19475 30784 19487 30787
rect 19978 30784 19984 30796
rect 19475 30756 19984 30784
rect 19475 30753 19487 30756
rect 19429 30747 19487 30753
rect 19978 30744 19984 30756
rect 20036 30744 20042 30796
rect 24026 30784 24032 30796
rect 23987 30756 24032 30784
rect 24026 30744 24032 30756
rect 24084 30744 24090 30796
rect 25041 30787 25099 30793
rect 25041 30753 25053 30787
rect 25087 30784 25099 30787
rect 25314 30784 25320 30796
rect 25087 30756 25320 30784
rect 25087 30753 25099 30756
rect 25041 30747 25099 30753
rect 25314 30744 25320 30756
rect 25372 30744 25378 30796
rect 35452 30793 35480 30824
rect 35437 30787 35495 30793
rect 35437 30753 35449 30787
rect 35483 30753 35495 30787
rect 35618 30784 35624 30796
rect 35579 30756 35624 30784
rect 35437 30747 35495 30753
rect 35618 30744 35624 30756
rect 35676 30784 35682 30796
rect 36173 30787 36231 30793
rect 36173 30784 36185 30787
rect 35676 30756 36185 30784
rect 35676 30744 35682 30756
rect 36173 30753 36185 30756
rect 36219 30753 36231 30787
rect 36354 30784 36360 30796
rect 36315 30756 36360 30784
rect 36173 30747 36231 30753
rect 36354 30744 36360 30756
rect 36412 30744 36418 30796
rect 11204 30688 12112 30716
rect 12437 30719 12495 30725
rect 11204 30676 11210 30688
rect 12437 30685 12449 30719
rect 12483 30685 12495 30719
rect 16482 30716 16488 30728
rect 16395 30688 16488 30716
rect 12437 30679 12495 30685
rect 12452 30648 12480 30679
rect 16482 30676 16488 30688
rect 16540 30716 16546 30728
rect 16669 30719 16727 30725
rect 16669 30716 16681 30719
rect 16540 30688 16681 30716
rect 16540 30676 16546 30688
rect 16669 30685 16681 30688
rect 16715 30685 16727 30719
rect 29086 30716 29092 30728
rect 29047 30688 29092 30716
rect 16669 30679 16727 30685
rect 29086 30676 29092 30688
rect 29144 30676 29150 30728
rect 29270 30676 29276 30728
rect 29328 30716 29334 30728
rect 29365 30719 29423 30725
rect 29365 30716 29377 30719
rect 29328 30688 29377 30716
rect 29328 30676 29334 30688
rect 29365 30685 29377 30688
rect 29411 30685 29423 30719
rect 36556 30716 36584 30824
rect 36722 30812 36728 30824
rect 36780 30812 36786 30864
rect 36832 30852 36860 30892
rect 36909 30889 36921 30923
rect 36955 30920 36967 30923
rect 57330 30920 57336 30932
rect 36955 30892 57336 30920
rect 36955 30889 36967 30892
rect 36909 30883 36967 30889
rect 57330 30880 57336 30892
rect 57388 30880 57394 30932
rect 57440 30892 59124 30920
rect 41598 30852 41604 30864
rect 36832 30824 41604 30852
rect 41598 30812 41604 30824
rect 41656 30812 41662 30864
rect 41782 30812 41788 30864
rect 41840 30852 41846 30864
rect 41840 30824 46428 30852
rect 41840 30812 41846 30824
rect 37093 30787 37151 30793
rect 37093 30753 37105 30787
rect 37139 30784 37151 30787
rect 37182 30784 37188 30796
rect 37139 30756 37188 30784
rect 37139 30753 37151 30756
rect 37093 30747 37151 30753
rect 37182 30744 37188 30756
rect 37240 30784 37246 30796
rect 37277 30787 37335 30793
rect 37277 30784 37289 30787
rect 37240 30756 37289 30784
rect 37240 30744 37246 30756
rect 37277 30753 37289 30756
rect 37323 30784 37335 30787
rect 37921 30787 37979 30793
rect 37921 30784 37933 30787
rect 37323 30756 37933 30784
rect 37323 30753 37335 30756
rect 37277 30747 37335 30753
rect 37550 30716 37556 30728
rect 36556 30688 37556 30716
rect 29365 30679 29423 30685
rect 37550 30676 37556 30688
rect 37608 30716 37614 30728
rect 37737 30719 37795 30725
rect 37737 30716 37749 30719
rect 37608 30688 37749 30716
rect 37608 30676 37614 30688
rect 37737 30685 37749 30688
rect 37783 30685 37795 30719
rect 37737 30679 37795 30685
rect 12526 30648 12532 30660
rect 12452 30620 12532 30648
rect 12526 30608 12532 30620
rect 12584 30608 12590 30660
rect 12805 30651 12863 30657
rect 12805 30617 12817 30651
rect 12851 30648 12863 30651
rect 15378 30648 15384 30660
rect 12851 30620 15384 30648
rect 12851 30617 12863 30620
rect 12805 30611 12863 30617
rect 4062 30540 4068 30592
rect 4120 30580 4126 30592
rect 6273 30583 6331 30589
rect 6273 30580 6285 30583
rect 4120 30552 6285 30580
rect 4120 30540 4126 30552
rect 6273 30549 6285 30552
rect 6319 30549 6331 30583
rect 6638 30580 6644 30592
rect 6599 30552 6644 30580
rect 6273 30543 6331 30549
rect 6638 30540 6644 30552
rect 6696 30540 6702 30592
rect 11698 30540 11704 30592
rect 11756 30580 11762 30592
rect 12820 30580 12848 30611
rect 15378 30608 15384 30620
rect 15436 30608 15442 30660
rect 30650 30648 30656 30660
rect 30563 30620 30656 30648
rect 30650 30608 30656 30620
rect 30708 30648 30714 30660
rect 36909 30651 36967 30657
rect 36909 30648 36921 30651
rect 30708 30620 36921 30648
rect 30708 30608 30714 30620
rect 36909 30617 36921 30620
rect 36955 30617 36967 30651
rect 36909 30611 36967 30617
rect 11756 30552 12848 30580
rect 11756 30540 11762 30552
rect 17402 30540 17408 30592
rect 17460 30580 17466 30592
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 17460 30552 19625 30580
rect 17460 30540 17466 30552
rect 19613 30549 19625 30552
rect 19659 30580 19671 30583
rect 19886 30580 19892 30592
rect 19659 30552 19892 30580
rect 19659 30549 19671 30552
rect 19613 30543 19671 30549
rect 19886 30540 19892 30552
rect 19944 30540 19950 30592
rect 24118 30580 24124 30592
rect 24079 30552 24124 30580
rect 24118 30540 24124 30552
rect 24176 30540 24182 30592
rect 36354 30540 36360 30592
rect 36412 30580 36418 30592
rect 37458 30580 37464 30592
rect 36412 30552 37464 30580
rect 36412 30540 36418 30552
rect 37458 30540 37464 30552
rect 37516 30540 37522 30592
rect 37844 30580 37872 30756
rect 37921 30753 37933 30756
rect 37967 30753 37979 30787
rect 38381 30787 38439 30793
rect 38381 30784 38393 30787
rect 37921 30747 37979 30753
rect 38120 30756 38393 30784
rect 38010 30676 38016 30728
rect 38068 30716 38074 30728
rect 38120 30716 38148 30756
rect 38381 30753 38393 30756
rect 38427 30753 38439 30787
rect 38381 30747 38439 30753
rect 38473 30787 38531 30793
rect 38473 30753 38485 30787
rect 38519 30784 38531 30787
rect 38654 30784 38660 30796
rect 38519 30756 38660 30784
rect 38519 30753 38531 30756
rect 38473 30747 38531 30753
rect 38654 30744 38660 30756
rect 38712 30744 38718 30796
rect 40954 30744 40960 30796
rect 41012 30784 41018 30796
rect 41141 30787 41199 30793
rect 41012 30756 41057 30784
rect 41012 30744 41018 30756
rect 41141 30753 41153 30787
rect 41187 30784 41199 30787
rect 41690 30784 41696 30796
rect 41187 30756 41696 30784
rect 41187 30753 41199 30756
rect 41141 30747 41199 30753
rect 40770 30716 40776 30728
rect 38068 30688 38148 30716
rect 40731 30688 40776 30716
rect 38068 30676 38074 30688
rect 40770 30676 40776 30688
rect 40828 30676 40834 30728
rect 38286 30608 38292 30660
rect 38344 30648 38350 30660
rect 38841 30651 38899 30657
rect 38841 30648 38853 30651
rect 38344 30620 38853 30648
rect 38344 30608 38350 30620
rect 38841 30617 38853 30620
rect 38887 30617 38899 30651
rect 40494 30648 40500 30660
rect 40407 30620 40500 30648
rect 38841 30611 38899 30617
rect 40494 30608 40500 30620
rect 40552 30648 40558 30660
rect 40681 30651 40739 30657
rect 40681 30648 40693 30651
rect 40552 30620 40693 30648
rect 40552 30608 40558 30620
rect 40681 30617 40693 30620
rect 40727 30648 40739 30651
rect 41156 30648 41184 30747
rect 41690 30744 41696 30756
rect 41748 30744 41754 30796
rect 41874 30784 41880 30796
rect 41835 30756 41880 30784
rect 41874 30744 41880 30756
rect 41932 30784 41938 30796
rect 42426 30784 42432 30796
rect 41932 30756 42432 30784
rect 41932 30744 41938 30756
rect 42426 30744 42432 30756
rect 42484 30744 42490 30796
rect 43162 30744 43168 30796
rect 43220 30784 43226 30796
rect 43349 30787 43407 30793
rect 43349 30784 43361 30787
rect 43220 30756 43361 30784
rect 43220 30744 43226 30756
rect 43349 30753 43361 30756
rect 43395 30784 43407 30787
rect 43530 30784 43536 30796
rect 43395 30756 43536 30784
rect 43395 30753 43407 30756
rect 43349 30747 43407 30753
rect 43530 30744 43536 30756
rect 43588 30744 43594 30796
rect 46400 30793 46428 30824
rect 46385 30787 46443 30793
rect 46385 30753 46397 30787
rect 46431 30784 46443 30787
rect 46937 30787 46995 30793
rect 46937 30784 46949 30787
rect 46431 30756 46949 30784
rect 46431 30753 46443 30756
rect 46385 30747 46443 30753
rect 46937 30753 46949 30756
rect 46983 30753 46995 30787
rect 46937 30747 46995 30753
rect 47121 30787 47179 30793
rect 47121 30753 47133 30787
rect 47167 30784 47179 30787
rect 49234 30784 49240 30796
rect 47167 30756 49096 30784
rect 49195 30756 49240 30784
rect 47167 30753 47179 30756
rect 47121 30747 47179 30753
rect 42245 30719 42303 30725
rect 42245 30685 42257 30719
rect 42291 30716 42303 30719
rect 43622 30716 43628 30728
rect 42291 30688 43628 30716
rect 42291 30685 42303 30688
rect 42245 30679 42303 30685
rect 43622 30676 43628 30688
rect 43680 30676 43686 30728
rect 46201 30719 46259 30725
rect 46201 30685 46213 30719
rect 46247 30685 46259 30719
rect 46201 30679 46259 30685
rect 40727 30620 41184 30648
rect 40727 30617 40739 30620
rect 40681 30611 40739 30617
rect 41598 30608 41604 30660
rect 41656 30648 41662 30660
rect 46017 30651 46075 30657
rect 46017 30648 46029 30651
rect 41656 30620 46029 30648
rect 41656 30608 41662 30620
rect 46017 30617 46029 30620
rect 46063 30648 46075 30651
rect 46216 30648 46244 30679
rect 48498 30676 48504 30728
rect 48556 30716 48562 30728
rect 48961 30719 49019 30725
rect 48961 30716 48973 30719
rect 48556 30688 48973 30716
rect 48556 30676 48562 30688
rect 46934 30648 46940 30660
rect 46063 30620 46940 30648
rect 46063 30617 46075 30620
rect 46017 30611 46075 30617
rect 46934 30608 46940 30620
rect 46992 30608 46998 30660
rect 47486 30648 47492 30660
rect 47044 30620 47492 30648
rect 38654 30580 38660 30592
rect 37844 30552 38660 30580
rect 38654 30540 38660 30552
rect 38712 30580 38718 30592
rect 43254 30580 43260 30592
rect 38712 30552 43260 30580
rect 38712 30540 38718 30552
rect 43254 30540 43260 30552
rect 43312 30540 43318 30592
rect 43438 30580 43444 30592
rect 43399 30552 43444 30580
rect 43438 30540 43444 30552
rect 43496 30540 43502 30592
rect 43530 30540 43536 30592
rect 43588 30580 43594 30592
rect 43717 30583 43775 30589
rect 43717 30580 43729 30583
rect 43588 30552 43729 30580
rect 43588 30540 43594 30552
rect 43717 30549 43729 30552
rect 43763 30580 43775 30583
rect 47044 30580 47072 30620
rect 47486 30608 47492 30620
rect 47544 30608 47550 30660
rect 48792 30592 48820 30688
rect 48961 30685 48973 30688
rect 49007 30685 49019 30719
rect 49068 30716 49096 30756
rect 49234 30744 49240 30756
rect 49292 30744 49298 30796
rect 54018 30744 54024 30796
rect 54076 30784 54082 30796
rect 54573 30787 54631 30793
rect 54573 30784 54585 30787
rect 54076 30756 54585 30784
rect 54076 30744 54082 30756
rect 54573 30753 54585 30756
rect 54619 30753 54631 30787
rect 56226 30784 56232 30796
rect 56139 30756 56232 30784
rect 54573 30747 54631 30753
rect 56226 30744 56232 30756
rect 56284 30784 56290 30796
rect 57440 30793 57468 30892
rect 57624 30824 59032 30852
rect 57624 30793 57652 30824
rect 56413 30787 56471 30793
rect 56413 30784 56425 30787
rect 56284 30756 56425 30784
rect 56284 30744 56290 30756
rect 56413 30753 56425 30756
rect 56459 30784 56471 30787
rect 56873 30787 56931 30793
rect 56873 30784 56885 30787
rect 56459 30756 56885 30784
rect 56459 30753 56471 30756
rect 56413 30747 56471 30753
rect 56873 30753 56885 30756
rect 56919 30784 56931 30787
rect 57425 30787 57483 30793
rect 57425 30784 57437 30787
rect 56919 30756 57437 30784
rect 56919 30753 56931 30756
rect 56873 30747 56931 30753
rect 57425 30753 57437 30756
rect 57471 30753 57483 30787
rect 57425 30747 57483 30753
rect 57609 30787 57667 30793
rect 57609 30753 57621 30787
rect 57655 30753 57667 30787
rect 57609 30747 57667 30753
rect 58710 30744 58716 30796
rect 58768 30784 58774 30796
rect 58897 30787 58955 30793
rect 58897 30784 58909 30787
rect 58768 30756 58909 30784
rect 58768 30744 58774 30756
rect 58897 30753 58909 30756
rect 58943 30753 58955 30787
rect 58897 30747 58955 30753
rect 54110 30716 54116 30728
rect 49068 30688 54116 30716
rect 48961 30679 49019 30685
rect 54110 30676 54116 30688
rect 54168 30676 54174 30728
rect 56594 30716 56600 30728
rect 56507 30688 56600 30716
rect 56594 30676 56600 30688
rect 56652 30716 56658 30728
rect 56689 30719 56747 30725
rect 56689 30716 56701 30719
rect 56652 30688 56701 30716
rect 56652 30676 56658 30688
rect 56689 30685 56701 30688
rect 56735 30685 56747 30719
rect 56689 30679 56747 30685
rect 57790 30648 57796 30660
rect 57751 30620 57796 30648
rect 57790 30608 57796 30620
rect 57848 30608 57854 30660
rect 59004 30657 59032 30824
rect 59096 30716 59124 30892
rect 59170 30880 59176 30932
rect 59228 30920 59234 30932
rect 59228 30892 61056 30920
rect 59228 30880 59234 30892
rect 60918 30716 60924 30728
rect 59096 30688 60924 30716
rect 60918 30676 60924 30688
rect 60976 30676 60982 30728
rect 61028 30725 61056 30892
rect 62206 30880 62212 30932
rect 62264 30920 62270 30932
rect 66073 30923 66131 30929
rect 66073 30920 66085 30923
rect 62264 30892 66085 30920
rect 62264 30880 62270 30892
rect 66073 30889 66085 30892
rect 66119 30889 66131 30923
rect 67450 30920 67456 30932
rect 67411 30892 67456 30920
rect 66073 30883 66131 30889
rect 62390 30852 62396 30864
rect 61304 30824 62252 30852
rect 62351 30824 62396 30852
rect 61304 30793 61332 30824
rect 61289 30787 61347 30793
rect 61289 30753 61301 30787
rect 61335 30753 61347 30787
rect 61289 30747 61347 30753
rect 61654 30744 61660 30796
rect 61712 30784 61718 30796
rect 61930 30793 61936 30796
rect 61755 30787 61813 30793
rect 61755 30784 61767 30787
rect 61712 30756 61767 30784
rect 61712 30744 61718 30756
rect 61755 30753 61767 30756
rect 61801 30753 61813 30787
rect 61929 30784 61936 30793
rect 61891 30756 61936 30784
rect 61755 30747 61813 30753
rect 61929 30747 61936 30756
rect 61930 30744 61936 30747
rect 61988 30744 61994 30796
rect 62224 30784 62252 30824
rect 62390 30812 62396 30824
rect 62448 30812 62454 30864
rect 66088 30852 66116 30883
rect 67450 30880 67456 30892
rect 67508 30880 67514 30932
rect 67542 30880 67548 30932
rect 67600 30920 67606 30932
rect 68281 30923 68339 30929
rect 68281 30920 68293 30923
rect 67600 30892 68293 30920
rect 67600 30880 67606 30892
rect 68281 30889 68293 30892
rect 68327 30920 68339 30923
rect 68327 30892 68600 30920
rect 68327 30889 68339 30892
rect 68281 30883 68339 30889
rect 68097 30855 68155 30861
rect 68097 30852 68109 30855
rect 66088 30824 68109 30852
rect 66916 30793 66944 30824
rect 68097 30821 68109 30824
rect 68143 30852 68155 30855
rect 68143 30824 68508 30852
rect 68143 30821 68155 30824
rect 68097 30815 68155 30821
rect 62761 30787 62819 30793
rect 62761 30784 62773 30787
rect 62224 30756 62773 30784
rect 62761 30753 62773 30756
rect 62807 30784 62819 30787
rect 66441 30787 66499 30793
rect 66441 30784 66453 30787
rect 62807 30756 66453 30784
rect 62807 30753 62819 30756
rect 62761 30747 62819 30753
rect 66441 30753 66453 30756
rect 66487 30784 66499 30787
rect 66901 30787 66959 30793
rect 66487 30756 66668 30784
rect 66487 30753 66499 30756
rect 66441 30747 66499 30753
rect 61013 30719 61071 30725
rect 61013 30685 61025 30719
rect 61059 30716 61071 30719
rect 61105 30719 61163 30725
rect 61105 30716 61117 30719
rect 61059 30688 61117 30716
rect 61059 30685 61071 30688
rect 61013 30679 61071 30685
rect 61105 30685 61117 30688
rect 61151 30685 61163 30719
rect 61105 30679 61163 30685
rect 66257 30719 66315 30725
rect 66257 30685 66269 30719
rect 66303 30685 66315 30719
rect 66257 30679 66315 30685
rect 58989 30651 59047 30657
rect 58989 30617 59001 30651
rect 59035 30648 59047 30651
rect 66272 30648 66300 30679
rect 59035 30620 66300 30648
rect 66640 30648 66668 30756
rect 66901 30753 66913 30787
rect 66947 30753 66959 30787
rect 66901 30747 66959 30753
rect 66990 30744 66996 30796
rect 67048 30784 67054 30796
rect 67726 30784 67732 30796
rect 67048 30756 67732 30784
rect 67048 30744 67054 30756
rect 67726 30744 67732 30756
rect 67784 30744 67790 30796
rect 68480 30793 68508 30824
rect 68465 30787 68523 30793
rect 68465 30753 68477 30787
rect 68511 30753 68523 30787
rect 68465 30747 68523 30753
rect 68002 30716 68008 30728
rect 67376 30688 68008 30716
rect 67376 30648 67404 30688
rect 68002 30676 68008 30688
rect 68060 30676 68066 30728
rect 68572 30716 68600 30892
rect 69474 30880 69480 30932
rect 69532 30920 69538 30932
rect 69661 30923 69719 30929
rect 69661 30920 69673 30923
rect 69532 30892 69673 30920
rect 69532 30880 69538 30892
rect 69661 30889 69673 30892
rect 69707 30889 69719 30923
rect 69661 30883 69719 30889
rect 69750 30880 69756 30932
rect 69808 30920 69814 30932
rect 84654 30920 84660 30932
rect 69808 30892 84660 30920
rect 69808 30880 69814 30892
rect 84654 30880 84660 30892
rect 84712 30880 84718 30932
rect 85114 30880 85120 30932
rect 85172 30920 85178 30932
rect 86221 30923 86279 30929
rect 86221 30920 86233 30923
rect 85172 30892 86233 30920
rect 85172 30880 85178 30892
rect 86221 30889 86233 30892
rect 86267 30889 86279 30923
rect 87966 30920 87972 30932
rect 87927 30892 87972 30920
rect 86221 30883 86279 30889
rect 70026 30852 70032 30864
rect 68664 30824 70032 30852
rect 68664 30793 68692 30824
rect 70026 30812 70032 30824
rect 70084 30812 70090 30864
rect 72510 30812 72516 30864
rect 72568 30852 72574 30864
rect 74813 30855 74871 30861
rect 74813 30852 74825 30855
rect 72568 30824 74825 30852
rect 72568 30812 72574 30824
rect 74813 30821 74825 30824
rect 74859 30821 74871 30855
rect 74813 30815 74871 30821
rect 75089 30855 75147 30861
rect 75089 30821 75101 30855
rect 75135 30852 75147 30855
rect 75181 30855 75239 30861
rect 75181 30852 75193 30855
rect 75135 30824 75193 30852
rect 75135 30821 75147 30824
rect 75089 30815 75147 30821
rect 75181 30821 75193 30824
rect 75227 30852 75239 30855
rect 76006 30852 76012 30864
rect 75227 30824 76012 30852
rect 75227 30821 75239 30824
rect 75181 30815 75239 30821
rect 68649 30787 68707 30793
rect 68649 30753 68661 30787
rect 68695 30753 68707 30787
rect 69109 30787 69167 30793
rect 69109 30784 69121 30787
rect 68649 30747 68707 30753
rect 68756 30756 69121 30784
rect 68756 30716 68784 30756
rect 69109 30753 69121 30756
rect 69155 30753 69167 30787
rect 69109 30747 69167 30753
rect 69198 30744 69204 30796
rect 69256 30784 69262 30796
rect 70121 30787 70179 30793
rect 70121 30784 70133 30787
rect 69256 30756 70133 30784
rect 69256 30744 69262 30756
rect 70121 30753 70133 30756
rect 70167 30753 70179 30787
rect 73706 30784 73712 30796
rect 73667 30756 73712 30784
rect 70121 30747 70179 30753
rect 73706 30744 73712 30756
rect 73764 30744 73770 30796
rect 74169 30787 74227 30793
rect 74169 30784 74181 30787
rect 73816 30756 74181 30784
rect 68572 30688 68784 30716
rect 73154 30676 73160 30728
rect 73212 30716 73218 30728
rect 73525 30719 73583 30725
rect 73525 30716 73537 30719
rect 73212 30688 73537 30716
rect 73212 30676 73218 30688
rect 73525 30685 73537 30688
rect 73571 30716 73583 30719
rect 73816 30716 73844 30756
rect 74169 30753 74181 30756
rect 74215 30753 74227 30787
rect 74169 30747 74227 30753
rect 74258 30744 74264 30796
rect 74316 30784 74322 30796
rect 75104 30784 75132 30815
rect 76006 30812 76012 30824
rect 76064 30812 76070 30864
rect 82814 30852 82820 30864
rect 79520 30824 82820 30852
rect 79520 30793 79548 30824
rect 82814 30812 82820 30824
rect 82872 30812 82878 30864
rect 83182 30812 83188 30864
rect 83240 30852 83246 30864
rect 83737 30855 83795 30861
rect 83737 30852 83749 30855
rect 83240 30824 83749 30852
rect 83240 30812 83246 30824
rect 83737 30821 83749 30824
rect 83783 30852 83795 30855
rect 83918 30852 83924 30864
rect 83783 30824 83924 30852
rect 83783 30821 83795 30824
rect 83737 30815 83795 30821
rect 83918 30812 83924 30824
rect 83976 30812 83982 30864
rect 86236 30852 86264 30883
rect 87966 30880 87972 30892
rect 88024 30880 88030 30932
rect 88242 30880 88248 30932
rect 88300 30920 88306 30932
rect 89717 30923 89775 30929
rect 89717 30920 89729 30923
rect 88300 30892 89729 30920
rect 88300 30880 88306 30892
rect 89717 30889 89729 30892
rect 89763 30889 89775 30923
rect 89717 30883 89775 30889
rect 86405 30855 86463 30861
rect 86405 30852 86417 30855
rect 86236 30824 86417 30852
rect 86405 30821 86417 30824
rect 86451 30821 86463 30855
rect 86405 30815 86463 30821
rect 74316 30756 75132 30784
rect 79505 30787 79563 30793
rect 74316 30744 74322 30756
rect 79505 30753 79517 30787
rect 79551 30753 79563 30787
rect 79505 30747 79563 30753
rect 79594 30744 79600 30796
rect 79652 30784 79658 30796
rect 79870 30784 79876 30796
rect 79652 30756 79697 30784
rect 79783 30756 79876 30784
rect 79652 30744 79658 30756
rect 79870 30744 79876 30756
rect 79928 30784 79934 30796
rect 80882 30784 80888 30796
rect 79928 30756 80100 30784
rect 80795 30756 80888 30784
rect 79928 30744 79934 30756
rect 73571 30688 73844 30716
rect 78769 30719 78827 30725
rect 73571 30685 73583 30688
rect 73525 30679 73583 30685
rect 78769 30685 78781 30719
rect 78815 30716 78827 30719
rect 79612 30716 79640 30744
rect 78815 30688 79640 30716
rect 78815 30685 78827 30688
rect 78769 30679 78827 30685
rect 79778 30676 79784 30728
rect 79836 30716 79842 30728
rect 79965 30719 80023 30725
rect 79965 30716 79977 30719
rect 79836 30688 79977 30716
rect 79836 30676 79842 30688
rect 79965 30685 79977 30688
rect 80011 30685 80023 30719
rect 79965 30679 80023 30685
rect 66640 30620 67404 30648
rect 59035 30617 59047 30620
rect 58989 30611 59047 30617
rect 69658 30608 69664 30660
rect 69716 30648 69722 30660
rect 80072 30648 80100 30756
rect 80882 30744 80888 30756
rect 80940 30744 80946 30796
rect 84194 30744 84200 30796
rect 84252 30784 84258 30796
rect 86586 30784 86592 30796
rect 84252 30756 84297 30784
rect 86547 30756 86592 30784
rect 84252 30744 84258 30756
rect 86586 30744 86592 30756
rect 86644 30744 86650 30796
rect 87984 30784 88012 30880
rect 88337 30787 88395 30793
rect 88337 30784 88349 30787
rect 87984 30756 88349 30784
rect 88337 30753 88349 30756
rect 88383 30753 88395 30787
rect 88610 30784 88616 30796
rect 88571 30756 88616 30784
rect 88337 30747 88395 30753
rect 88610 30744 88616 30756
rect 88668 30744 88674 30796
rect 80698 30716 80704 30728
rect 80659 30688 80704 30716
rect 80698 30676 80704 30688
rect 80756 30716 80762 30728
rect 80900 30716 80928 30744
rect 83918 30716 83924 30728
rect 80756 30688 80928 30716
rect 83879 30688 83924 30716
rect 80756 30676 80762 30688
rect 83918 30676 83924 30688
rect 83976 30676 83982 30728
rect 80149 30651 80207 30657
rect 80149 30648 80161 30651
rect 69716 30620 80161 30648
rect 69716 30608 69722 30620
rect 80149 30617 80161 30620
rect 80195 30648 80207 30651
rect 81069 30651 81127 30657
rect 81069 30648 81081 30651
rect 80195 30620 81081 30648
rect 80195 30617 80207 30620
rect 80149 30611 80207 30617
rect 81069 30617 81081 30620
rect 81115 30617 81127 30651
rect 81069 30611 81127 30617
rect 82354 30608 82360 30660
rect 82412 30648 82418 30660
rect 82412 30620 83872 30648
rect 82412 30608 82418 30620
rect 43763 30552 47072 30580
rect 43763 30549 43775 30552
rect 43717 30543 43775 30549
rect 47210 30540 47216 30592
rect 47268 30580 47274 30592
rect 47397 30583 47455 30589
rect 47397 30580 47409 30583
rect 47268 30552 47409 30580
rect 47268 30540 47274 30552
rect 47397 30549 47409 30552
rect 47443 30549 47455 30583
rect 48774 30580 48780 30592
rect 48735 30552 48780 30580
rect 47397 30543 47455 30549
rect 48774 30540 48780 30552
rect 48832 30540 48838 30592
rect 50154 30540 50160 30592
rect 50212 30580 50218 30592
rect 50341 30583 50399 30589
rect 50341 30580 50353 30583
rect 50212 30552 50353 30580
rect 50212 30540 50218 30552
rect 50341 30549 50353 30552
rect 50387 30549 50399 30583
rect 54662 30580 54668 30592
rect 54623 30552 54668 30580
rect 50341 30543 50399 30549
rect 54662 30540 54668 30552
rect 54720 30580 54726 30592
rect 59078 30580 59084 30592
rect 54720 30552 59084 30580
rect 54720 30540 54726 30552
rect 59078 30540 59084 30552
rect 59136 30540 59142 30592
rect 59170 30540 59176 30592
rect 59228 30580 59234 30592
rect 59228 30552 59273 30580
rect 59228 30540 59234 30552
rect 60366 30540 60372 30592
rect 60424 30580 60430 30592
rect 60737 30583 60795 30589
rect 60737 30580 60749 30583
rect 60424 30552 60749 30580
rect 60424 30540 60430 30552
rect 60737 30549 60749 30552
rect 60783 30580 60795 30583
rect 61654 30580 61660 30592
rect 60783 30552 61660 30580
rect 60783 30549 60795 30552
rect 60737 30543 60795 30549
rect 61654 30540 61660 30552
rect 61712 30540 61718 30592
rect 61930 30540 61936 30592
rect 61988 30580 61994 30592
rect 62669 30583 62727 30589
rect 62669 30580 62681 30583
rect 61988 30552 62681 30580
rect 61988 30540 61994 30552
rect 62669 30549 62681 30552
rect 62715 30580 62727 30583
rect 66990 30580 66996 30592
rect 62715 30552 66996 30580
rect 62715 30549 62727 30552
rect 62669 30543 62727 30549
rect 66990 30540 66996 30552
rect 67048 30540 67054 30592
rect 67726 30580 67732 30592
rect 67687 30552 67732 30580
rect 67726 30540 67732 30552
rect 67784 30540 67790 30592
rect 68002 30580 68008 30592
rect 67915 30552 68008 30580
rect 68002 30540 68008 30552
rect 68060 30580 68066 30592
rect 69750 30580 69756 30592
rect 68060 30552 69756 30580
rect 68060 30540 68066 30552
rect 69750 30540 69756 30552
rect 69808 30540 69814 30592
rect 70026 30580 70032 30592
rect 69987 30552 70032 30580
rect 70026 30540 70032 30552
rect 70084 30540 70090 30592
rect 73154 30580 73160 30592
rect 73115 30552 73160 30580
rect 73154 30540 73160 30552
rect 73212 30580 73218 30592
rect 73341 30583 73399 30589
rect 73341 30580 73353 30583
rect 73212 30552 73353 30580
rect 73212 30540 73218 30552
rect 73341 30549 73353 30552
rect 73387 30549 73399 30583
rect 73341 30543 73399 30549
rect 78953 30583 79011 30589
rect 78953 30549 78965 30583
rect 78999 30580 79011 30583
rect 79226 30580 79232 30592
rect 78999 30552 79232 30580
rect 78999 30549 79011 30552
rect 78953 30543 79011 30549
rect 79226 30540 79232 30552
rect 79284 30540 79290 30592
rect 83844 30580 83872 30620
rect 85224 30620 86724 30648
rect 85224 30580 85252 30620
rect 83844 30552 85252 30580
rect 85298 30540 85304 30592
rect 85356 30580 85362 30592
rect 86696 30589 86724 30620
rect 86681 30583 86739 30589
rect 85356 30552 85401 30580
rect 85356 30540 85362 30552
rect 86681 30549 86693 30583
rect 86727 30549 86739 30583
rect 86681 30543 86739 30549
rect 1104 30490 108008 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 65686 30490
rect 65738 30438 65750 30490
rect 65802 30438 65814 30490
rect 65866 30438 65878 30490
rect 65930 30438 96406 30490
rect 96458 30438 96470 30490
rect 96522 30438 96534 30490
rect 96586 30438 96598 30490
rect 96650 30438 108008 30490
rect 1104 30416 108008 30438
rect 3602 30336 3608 30388
rect 3660 30376 3666 30388
rect 4890 30376 4896 30388
rect 3660 30348 4896 30376
rect 3660 30336 3666 30348
rect 4890 30336 4896 30348
rect 4948 30336 4954 30388
rect 10686 30336 10692 30388
rect 10744 30376 10750 30388
rect 16482 30376 16488 30388
rect 10744 30348 16488 30376
rect 10744 30336 10750 30348
rect 16482 30336 16488 30348
rect 16540 30336 16546 30388
rect 31018 30376 31024 30388
rect 30979 30348 31024 30376
rect 31018 30336 31024 30348
rect 31076 30336 31082 30388
rect 37458 30336 37464 30388
rect 37516 30376 37522 30388
rect 38197 30379 38255 30385
rect 38197 30376 38209 30379
rect 37516 30348 38209 30376
rect 37516 30336 37522 30348
rect 38197 30345 38209 30348
rect 38243 30376 38255 30379
rect 38243 30348 53972 30376
rect 38243 30345 38255 30348
rect 38197 30339 38255 30345
rect 3878 30268 3884 30320
rect 3936 30308 3942 30320
rect 20070 30308 20076 30320
rect 3936 30280 20076 30308
rect 3936 30268 3942 30280
rect 20070 30268 20076 30280
rect 20128 30268 20134 30320
rect 26786 30308 26792 30320
rect 21744 30280 26792 30308
rect 2593 30243 2651 30249
rect 2593 30209 2605 30243
rect 2639 30240 2651 30243
rect 2958 30240 2964 30252
rect 2639 30212 2964 30240
rect 2639 30209 2651 30212
rect 2593 30203 2651 30209
rect 2958 30200 2964 30212
rect 3016 30200 3022 30252
rect 4617 30243 4675 30249
rect 4617 30209 4629 30243
rect 4663 30240 4675 30243
rect 4706 30240 4712 30252
rect 4663 30212 4712 30240
rect 4663 30209 4675 30212
rect 4617 30203 4675 30209
rect 4706 30200 4712 30212
rect 4764 30200 4770 30252
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30240 10011 30243
rect 18506 30240 18512 30252
rect 9999 30212 18512 30240
rect 9999 30209 10011 30212
rect 9953 30203 10011 30209
rect 2869 30175 2927 30181
rect 2869 30141 2881 30175
rect 2915 30172 2927 30175
rect 7929 30175 7987 30181
rect 2915 30144 4476 30172
rect 2915 30141 2927 30144
rect 2869 30135 2927 30141
rect 4448 30048 4476 30144
rect 7929 30141 7941 30175
rect 7975 30172 7987 30175
rect 9582 30172 9588 30184
rect 7975 30144 9588 30172
rect 7975 30141 7987 30144
rect 7929 30135 7987 30141
rect 9582 30132 9588 30144
rect 9640 30132 9646 30184
rect 10612 30181 10640 30212
rect 18506 30200 18512 30212
rect 18564 30240 18570 30252
rect 21744 30240 21772 30280
rect 26786 30268 26792 30280
rect 26844 30268 26850 30320
rect 28169 30311 28227 30317
rect 28169 30277 28181 30311
rect 28215 30308 28227 30311
rect 29270 30308 29276 30320
rect 28215 30280 29276 30308
rect 28215 30277 28227 30280
rect 28169 30271 28227 30277
rect 29270 30268 29276 30280
rect 29328 30268 29334 30320
rect 22462 30240 22468 30252
rect 18564 30212 21772 30240
rect 21836 30212 22468 30240
rect 18564 30200 18570 30212
rect 10597 30175 10655 30181
rect 10597 30141 10609 30175
rect 10643 30141 10655 30175
rect 10597 30135 10655 30141
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30141 10839 30175
rect 10781 30135 10839 30141
rect 10965 30175 11023 30181
rect 10965 30141 10977 30175
rect 11011 30172 11023 30175
rect 11146 30172 11152 30184
rect 11011 30144 11152 30172
rect 11011 30141 11023 30144
rect 10965 30135 11023 30141
rect 9950 30064 9956 30116
rect 10008 30104 10014 30116
rect 10045 30107 10103 30113
rect 10045 30104 10057 30107
rect 10008 30076 10057 30104
rect 10008 30064 10014 30076
rect 10045 30073 10057 30076
rect 10091 30073 10103 30107
rect 10045 30067 10103 30073
rect 3142 29996 3148 30048
rect 3200 30036 3206 30048
rect 3973 30039 4031 30045
rect 3973 30036 3985 30039
rect 3200 30008 3985 30036
rect 3200 29996 3206 30008
rect 3973 30005 3985 30008
rect 4019 30005 4031 30039
rect 4430 30036 4436 30048
rect 4391 30008 4436 30036
rect 3973 29999 4031 30005
rect 4430 29996 4436 30008
rect 4488 29996 4494 30048
rect 7742 30036 7748 30048
rect 7655 30008 7748 30036
rect 7742 29996 7748 30008
rect 7800 30036 7806 30048
rect 9674 30036 9680 30048
rect 7800 30008 9680 30036
rect 7800 29996 7806 30008
rect 9674 29996 9680 30008
rect 9732 30036 9738 30048
rect 10686 30036 10692 30048
rect 9732 30008 10692 30036
rect 9732 29996 9738 30008
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 10796 30036 10824 30135
rect 11146 30132 11152 30144
rect 11204 30132 11210 30184
rect 11333 30175 11391 30181
rect 11333 30141 11345 30175
rect 11379 30141 11391 30175
rect 11333 30135 11391 30141
rect 11517 30175 11575 30181
rect 11517 30141 11529 30175
rect 11563 30172 11575 30175
rect 12618 30172 12624 30184
rect 11563 30144 12624 30172
rect 11563 30141 11575 30144
rect 11517 30135 11575 30141
rect 11348 30104 11376 30135
rect 12618 30132 12624 30144
rect 12676 30132 12682 30184
rect 15473 30175 15531 30181
rect 15473 30141 15485 30175
rect 15519 30172 15531 30175
rect 15562 30172 15568 30184
rect 15519 30144 15568 30172
rect 15519 30141 15531 30144
rect 15473 30135 15531 30141
rect 15488 30104 15516 30135
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 19797 30175 19855 30181
rect 19797 30141 19809 30175
rect 19843 30172 19855 30175
rect 19978 30172 19984 30184
rect 19843 30144 19984 30172
rect 19843 30141 19855 30144
rect 19797 30135 19855 30141
rect 19978 30132 19984 30144
rect 20036 30132 20042 30184
rect 21836 30181 21864 30212
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 24670 30200 24676 30252
rect 24728 30240 24734 30252
rect 25041 30243 25099 30249
rect 25041 30240 25053 30243
rect 24728 30212 25053 30240
rect 24728 30200 24734 30212
rect 25041 30209 25053 30212
rect 25087 30209 25099 30243
rect 28994 30240 29000 30252
rect 25041 30203 25099 30209
rect 28460 30212 29000 30240
rect 21821 30175 21879 30181
rect 21821 30141 21833 30175
rect 21867 30141 21879 30175
rect 22005 30175 22063 30181
rect 22005 30172 22017 30175
rect 21821 30135 21879 30141
rect 21928 30144 22017 30172
rect 21928 30104 21956 30144
rect 22005 30141 22017 30144
rect 22051 30141 22063 30175
rect 24762 30172 24768 30184
rect 22005 30135 22063 30141
rect 22112 30144 24624 30172
rect 24723 30144 24768 30172
rect 11348 30076 11928 30104
rect 15488 30076 21956 30104
rect 11900 30048 11928 30076
rect 11609 30039 11667 30045
rect 11609 30036 11621 30039
rect 10796 30008 11621 30036
rect 11609 30005 11621 30008
rect 11655 30036 11667 30039
rect 11698 30036 11704 30048
rect 11655 30008 11704 30036
rect 11655 30005 11667 30008
rect 11609 29999 11667 30005
rect 11698 29996 11704 30008
rect 11756 29996 11762 30048
rect 11882 30036 11888 30048
rect 11843 30008 11888 30036
rect 11882 29996 11888 30008
rect 11940 29996 11946 30048
rect 15562 30036 15568 30048
rect 15523 30008 15568 30036
rect 15562 29996 15568 30008
rect 15620 29996 15626 30048
rect 19978 30036 19984 30048
rect 19891 30008 19984 30036
rect 19978 29996 19984 30008
rect 20036 30036 20042 30048
rect 20806 30036 20812 30048
rect 20036 30008 20812 30036
rect 20036 29996 20042 30008
rect 20806 29996 20812 30008
rect 20864 29996 20870 30048
rect 20898 29996 20904 30048
rect 20956 30036 20962 30048
rect 22112 30036 22140 30144
rect 22278 30104 22284 30116
rect 22239 30076 22284 30104
rect 22278 30064 22284 30076
rect 22336 30064 22342 30116
rect 24596 30104 24624 30144
rect 24762 30132 24768 30144
rect 24820 30132 24826 30184
rect 24946 30172 24952 30184
rect 24859 30144 24952 30172
rect 24946 30132 24952 30144
rect 25004 30132 25010 30184
rect 25409 30175 25467 30181
rect 25409 30141 25421 30175
rect 25455 30172 25467 30175
rect 26326 30172 26332 30184
rect 25455 30144 26332 30172
rect 25455 30141 25467 30144
rect 25409 30135 25467 30141
rect 26326 30132 26332 30144
rect 26384 30132 26390 30184
rect 26973 30175 27031 30181
rect 26973 30141 26985 30175
rect 27019 30141 27031 30175
rect 27154 30172 27160 30184
rect 27115 30144 27160 30172
rect 26973 30135 27031 30141
rect 24964 30104 24992 30132
rect 24596 30076 24992 30104
rect 22462 30036 22468 30048
rect 20956 30008 22140 30036
rect 22375 30008 22468 30036
rect 20956 29996 20962 30008
rect 22462 29996 22468 30008
rect 22520 30036 22526 30048
rect 23290 30036 23296 30048
rect 22520 30008 23296 30036
rect 22520 29996 22526 30008
rect 23290 29996 23296 30008
rect 23348 29996 23354 30048
rect 23658 29996 23664 30048
rect 23716 30036 23722 30048
rect 26789 30039 26847 30045
rect 26789 30036 26801 30039
rect 23716 30008 26801 30036
rect 23716 29996 23722 30008
rect 26789 30005 26801 30008
rect 26835 30036 26847 30039
rect 26988 30036 27016 30135
rect 27154 30132 27160 30144
rect 27212 30132 27218 30184
rect 27246 30132 27252 30184
rect 27304 30172 27310 30184
rect 27798 30181 27804 30184
rect 27617 30175 27675 30181
rect 27617 30172 27629 30175
rect 27304 30144 27629 30172
rect 27304 30132 27310 30144
rect 27617 30141 27629 30144
rect 27663 30141 27675 30175
rect 27797 30172 27804 30181
rect 27759 30144 27804 30172
rect 27617 30135 27675 30141
rect 27797 30135 27804 30144
rect 27798 30132 27804 30135
rect 27856 30132 27862 30184
rect 26835 30008 27016 30036
rect 26835 30005 26847 30008
rect 26789 29999 26847 30005
rect 27246 29996 27252 30048
rect 27304 30036 27310 30048
rect 28460 30045 28488 30212
rect 28994 30200 29000 30212
rect 29052 30200 29058 30252
rect 29086 30200 29092 30252
rect 29144 30240 29150 30252
rect 31036 30240 31064 30336
rect 37550 30308 37556 30320
rect 37511 30280 37556 30308
rect 37550 30268 37556 30280
rect 37608 30268 37614 30320
rect 43162 30308 43168 30320
rect 43123 30280 43168 30308
rect 43162 30268 43168 30280
rect 43220 30268 43226 30320
rect 48774 30308 48780 30320
rect 48687 30280 48780 30308
rect 48774 30268 48780 30280
rect 48832 30308 48838 30320
rect 52549 30311 52607 30317
rect 52549 30308 52561 30311
rect 48832 30280 52561 30308
rect 48832 30268 48838 30280
rect 52549 30277 52561 30280
rect 52595 30308 52607 30311
rect 53944 30308 53972 30348
rect 54018 30336 54024 30388
rect 54076 30376 54082 30388
rect 54113 30379 54171 30385
rect 54113 30376 54125 30379
rect 54076 30348 54125 30376
rect 54076 30336 54082 30348
rect 54113 30345 54125 30348
rect 54159 30345 54171 30379
rect 60185 30379 60243 30385
rect 60185 30376 60197 30379
rect 54113 30339 54171 30345
rect 54220 30348 60197 30376
rect 54220 30308 54248 30348
rect 60185 30345 60197 30348
rect 60231 30376 60243 30379
rect 60458 30376 60464 30388
rect 60231 30348 60464 30376
rect 60231 30345 60243 30348
rect 60185 30339 60243 30345
rect 60458 30336 60464 30348
rect 60516 30336 60522 30388
rect 60918 30336 60924 30388
rect 60976 30376 60982 30388
rect 60976 30348 65748 30376
rect 60976 30336 60982 30348
rect 52595 30280 52776 30308
rect 53944 30280 54248 30308
rect 58636 30280 60780 30308
rect 52595 30277 52607 30280
rect 52549 30271 52607 30277
rect 52638 30240 52644 30252
rect 29144 30212 31064 30240
rect 32416 30212 52644 30240
rect 29144 30200 29150 30212
rect 29288 30181 29316 30212
rect 29273 30175 29331 30181
rect 29273 30141 29285 30175
rect 29319 30141 29331 30175
rect 29273 30135 29331 30141
rect 29362 30132 29368 30184
rect 29420 30172 29426 30184
rect 29549 30175 29607 30181
rect 29549 30172 29561 30175
rect 29420 30144 29561 30172
rect 29420 30132 29426 30144
rect 29549 30141 29561 30144
rect 29595 30141 29607 30175
rect 29549 30135 29607 30141
rect 29638 30132 29644 30184
rect 29696 30172 29702 30184
rect 32416 30172 32444 30212
rect 52638 30200 52644 30212
rect 52696 30200 52702 30252
rect 52748 30249 52776 30280
rect 52733 30243 52791 30249
rect 52733 30209 52745 30243
rect 52779 30209 52791 30243
rect 58636 30240 58664 30280
rect 52733 30203 52791 30209
rect 52840 30212 58664 30240
rect 29696 30144 32444 30172
rect 35621 30175 35679 30181
rect 29696 30132 29702 30144
rect 35621 30141 35633 30175
rect 35667 30172 35679 30175
rect 35710 30172 35716 30184
rect 35667 30144 35716 30172
rect 35667 30141 35679 30144
rect 35621 30135 35679 30141
rect 35710 30132 35716 30144
rect 35768 30132 35774 30184
rect 35897 30175 35955 30181
rect 35897 30141 35909 30175
rect 35943 30172 35955 30175
rect 37274 30172 37280 30184
rect 35943 30144 37280 30172
rect 35943 30141 35955 30144
rect 35897 30135 35955 30141
rect 37274 30132 37280 30144
rect 37332 30132 37338 30184
rect 37458 30172 37464 30184
rect 37371 30144 37464 30172
rect 37458 30132 37464 30144
rect 37516 30172 37522 30184
rect 37918 30172 37924 30184
rect 37516 30144 37924 30172
rect 37516 30132 37522 30144
rect 37918 30132 37924 30144
rect 37976 30132 37982 30184
rect 38010 30132 38016 30184
rect 38068 30172 38074 30184
rect 38105 30175 38163 30181
rect 38105 30172 38117 30175
rect 38068 30144 38117 30172
rect 38068 30132 38074 30144
rect 38105 30141 38117 30144
rect 38151 30141 38163 30175
rect 41598 30172 41604 30184
rect 41559 30144 41604 30172
rect 38105 30135 38163 30141
rect 41598 30132 41604 30144
rect 41656 30132 41662 30184
rect 41877 30175 41935 30181
rect 41877 30141 41889 30175
rect 41923 30172 41935 30175
rect 42242 30172 42248 30184
rect 41923 30144 42248 30172
rect 41923 30141 41935 30144
rect 41877 30135 41935 30141
rect 42242 30132 42248 30144
rect 42300 30132 42306 30184
rect 43346 30172 43352 30184
rect 43307 30144 43352 30172
rect 43346 30132 43352 30144
rect 43404 30132 43410 30184
rect 43622 30172 43628 30184
rect 43583 30144 43628 30172
rect 43622 30132 43628 30144
rect 43680 30132 43686 30184
rect 44726 30132 44732 30184
rect 44784 30172 44790 30184
rect 45462 30172 45468 30184
rect 44784 30144 45468 30172
rect 44784 30132 44790 30144
rect 45462 30132 45468 30144
rect 45520 30132 45526 30184
rect 46934 30172 46940 30184
rect 46895 30144 46940 30172
rect 46934 30132 46940 30144
rect 46992 30132 46998 30184
rect 47210 30172 47216 30184
rect 47171 30144 47216 30172
rect 47210 30132 47216 30144
rect 47268 30132 47274 30184
rect 47302 30132 47308 30184
rect 47360 30172 47366 30184
rect 48774 30172 48780 30184
rect 47360 30144 48780 30172
rect 47360 30132 47366 30144
rect 48774 30132 48780 30144
rect 48832 30132 48838 30184
rect 45002 30104 45008 30116
rect 36556 30076 38056 30104
rect 28445 30039 28503 30045
rect 28445 30036 28457 30039
rect 27304 30008 28457 30036
rect 27304 29996 27310 30008
rect 28445 30005 28457 30008
rect 28491 30005 28503 30039
rect 28718 30036 28724 30048
rect 28631 30008 28724 30036
rect 28445 29999 28503 30005
rect 28718 29996 28724 30008
rect 28776 30036 28782 30048
rect 28905 30039 28963 30045
rect 28905 30036 28917 30039
rect 28776 30008 28917 30036
rect 28776 29996 28782 30008
rect 28905 30005 28917 30008
rect 28951 30036 28963 30039
rect 29822 30036 29828 30048
rect 28951 30008 29828 30036
rect 28951 30005 28963 30008
rect 28905 29999 28963 30005
rect 29822 29996 29828 30008
rect 29880 29996 29886 30048
rect 30834 30036 30840 30048
rect 30747 30008 30840 30036
rect 30834 29996 30840 30008
rect 30892 30036 30898 30048
rect 36556 30036 36584 30076
rect 36998 30036 37004 30048
rect 30892 30008 36584 30036
rect 36959 30008 37004 30036
rect 30892 29996 30898 30008
rect 36998 29996 37004 30008
rect 37056 29996 37062 30048
rect 37918 30036 37924 30048
rect 37879 30008 37924 30036
rect 37918 29996 37924 30008
rect 37976 29996 37982 30048
rect 38028 30036 38056 30076
rect 42904 30076 43116 30104
rect 42904 30036 42932 30076
rect 38028 30008 42932 30036
rect 43088 30036 43116 30076
rect 44652 30076 44864 30104
rect 44915 30076 45008 30104
rect 44652 30036 44680 30076
rect 43088 30008 44680 30036
rect 44836 30036 44864 30076
rect 45002 30064 45008 30076
rect 45060 30104 45066 30116
rect 46842 30104 46848 30116
rect 45060 30076 46848 30104
rect 45060 30064 45066 30076
rect 46842 30064 46848 30076
rect 46900 30064 46906 30116
rect 52840 30104 52868 30212
rect 58710 30200 58716 30252
rect 58768 30240 58774 30252
rect 58805 30243 58863 30249
rect 58805 30240 58817 30243
rect 58768 30212 58817 30240
rect 58768 30200 58774 30212
rect 58805 30209 58817 30212
rect 58851 30240 58863 30243
rect 59170 30240 59176 30252
rect 58851 30212 59176 30240
rect 58851 30209 58863 30212
rect 58805 30203 58863 30209
rect 59170 30200 59176 30212
rect 59228 30200 59234 30252
rect 53006 30132 53012 30184
rect 53064 30172 53070 30184
rect 53064 30144 53109 30172
rect 53064 30132 53070 30144
rect 53282 30132 53288 30184
rect 53340 30172 53346 30184
rect 56778 30172 56784 30184
rect 53340 30144 56784 30172
rect 53340 30132 53346 30144
rect 56778 30132 56784 30144
rect 56836 30132 56842 30184
rect 57425 30175 57483 30181
rect 57425 30141 57437 30175
rect 57471 30141 57483 30175
rect 57425 30135 57483 30141
rect 57701 30175 57759 30181
rect 57701 30141 57713 30175
rect 57747 30172 57759 30175
rect 57790 30172 57796 30184
rect 57747 30144 57796 30172
rect 57747 30141 57759 30144
rect 57701 30135 57759 30141
rect 47872 30076 52868 30104
rect 47872 30036 47900 30076
rect 48314 30036 48320 30048
rect 44836 30008 47900 30036
rect 48275 30008 48320 30036
rect 48314 29996 48320 30008
rect 48372 29996 48378 30048
rect 51994 29996 52000 30048
rect 52052 30036 52058 30048
rect 56594 30036 56600 30048
rect 52052 30008 56600 30036
rect 52052 29996 52058 30008
rect 56594 29996 56600 30008
rect 56652 29996 56658 30048
rect 57440 30036 57468 30135
rect 57790 30132 57796 30144
rect 57848 30132 57854 30184
rect 59446 30132 59452 30184
rect 59504 30172 59510 30184
rect 59725 30175 59783 30181
rect 59725 30172 59737 30175
rect 59504 30144 59737 30172
rect 59504 30132 59510 30144
rect 59725 30141 59737 30144
rect 59771 30141 59783 30175
rect 60366 30172 60372 30184
rect 60279 30144 60372 30172
rect 59725 30135 59783 30141
rect 60366 30132 60372 30144
rect 60424 30132 60430 30184
rect 60553 30175 60611 30181
rect 60553 30141 60565 30175
rect 60599 30172 60611 30175
rect 60599 30144 60688 30172
rect 60599 30141 60611 30144
rect 60553 30135 60611 30141
rect 60182 30104 60188 30116
rect 59188 30076 60188 30104
rect 59188 30045 59216 30076
rect 60182 30064 60188 30076
rect 60240 30064 60246 30116
rect 59173 30039 59231 30045
rect 59173 30036 59185 30039
rect 57440 30008 59185 30036
rect 59173 30005 59185 30008
rect 59219 30005 59231 30039
rect 59173 29999 59231 30005
rect 59354 29996 59360 30048
rect 59412 30036 59418 30048
rect 59541 30039 59599 30045
rect 59541 30036 59553 30039
rect 59412 30008 59553 30036
rect 59412 29996 59418 30008
rect 59541 30005 59553 30008
rect 59587 30005 59599 30039
rect 59998 30036 60004 30048
rect 59959 30008 60004 30036
rect 59541 29999 59599 30005
rect 59998 29996 60004 30008
rect 60056 30036 60062 30048
rect 60384 30036 60412 30132
rect 60660 30048 60688 30144
rect 60056 30008 60412 30036
rect 60056 29996 60062 30008
rect 60642 29996 60648 30048
rect 60700 29996 60706 30048
rect 60752 30036 60780 30280
rect 61102 30268 61108 30320
rect 61160 30308 61166 30320
rect 61473 30311 61531 30317
rect 61473 30308 61485 30311
rect 61160 30280 61485 30308
rect 61160 30268 61166 30280
rect 61473 30277 61485 30280
rect 61519 30277 61531 30311
rect 61930 30308 61936 30320
rect 61891 30280 61936 30308
rect 61473 30271 61531 30277
rect 61930 30268 61936 30280
rect 61988 30268 61994 30320
rect 65720 30317 65748 30348
rect 67726 30336 67732 30388
rect 67784 30376 67790 30388
rect 69658 30376 69664 30388
rect 67784 30348 69664 30376
rect 67784 30336 67790 30348
rect 69658 30336 69664 30348
rect 69716 30336 69722 30388
rect 70026 30336 70032 30388
rect 70084 30376 70090 30388
rect 80698 30376 80704 30388
rect 70084 30348 80704 30376
rect 70084 30336 70090 30348
rect 80698 30336 80704 30348
rect 80756 30336 80762 30388
rect 84654 30376 84660 30388
rect 84567 30348 84660 30376
rect 84654 30336 84660 30348
rect 84712 30376 84718 30388
rect 85298 30376 85304 30388
rect 84712 30348 85304 30376
rect 84712 30336 84718 30348
rect 85298 30336 85304 30348
rect 85356 30336 85362 30388
rect 65705 30311 65763 30317
rect 65705 30277 65717 30311
rect 65751 30308 65763 30311
rect 65889 30311 65947 30317
rect 65889 30308 65901 30311
rect 65751 30280 65901 30308
rect 65751 30277 65763 30280
rect 65705 30271 65763 30277
rect 65889 30277 65901 30280
rect 65935 30277 65947 30311
rect 71409 30311 71467 30317
rect 71409 30308 71421 30311
rect 65889 30271 65947 30277
rect 66272 30280 71421 30308
rect 61013 30175 61071 30181
rect 61013 30141 61025 30175
rect 61059 30141 61071 30175
rect 61013 30135 61071 30141
rect 61193 30175 61251 30181
rect 61193 30141 61205 30175
rect 61239 30172 61251 30175
rect 62022 30172 62028 30184
rect 61239 30144 62028 30172
rect 61239 30141 61251 30144
rect 61193 30135 61251 30141
rect 60826 30064 60832 30116
rect 60884 30104 60890 30116
rect 61028 30104 61056 30135
rect 62022 30132 62028 30144
rect 62080 30132 62086 30184
rect 65904 30172 65932 30271
rect 66070 30200 66076 30252
rect 66128 30240 66134 30252
rect 66272 30249 66300 30280
rect 71409 30277 71421 30280
rect 71455 30308 71467 30311
rect 71590 30308 71596 30320
rect 71455 30280 71596 30308
rect 71455 30277 71467 30280
rect 71409 30271 71467 30277
rect 71590 30268 71596 30280
rect 71648 30268 71654 30320
rect 84381 30311 84439 30317
rect 84381 30277 84393 30311
rect 84427 30308 84439 30311
rect 85114 30308 85120 30320
rect 84427 30280 85120 30308
rect 84427 30277 84439 30280
rect 84381 30271 84439 30277
rect 85114 30268 85120 30280
rect 85172 30268 85178 30320
rect 66257 30243 66315 30249
rect 66257 30240 66269 30243
rect 66128 30212 66269 30240
rect 66128 30200 66134 30212
rect 66257 30209 66269 30212
rect 66303 30209 66315 30243
rect 68649 30243 68707 30249
rect 68649 30240 68661 30243
rect 66257 30203 66315 30209
rect 66456 30212 66668 30240
rect 66456 30181 66484 30212
rect 66441 30175 66499 30181
rect 66441 30172 66453 30175
rect 65904 30144 66453 30172
rect 66441 30141 66453 30144
rect 66487 30141 66499 30175
rect 66640 30172 66668 30212
rect 67560 30212 68661 30240
rect 66993 30175 67051 30181
rect 66993 30172 67005 30175
rect 66640 30144 67005 30172
rect 66441 30135 66499 30141
rect 66993 30141 67005 30144
rect 67039 30141 67051 30175
rect 66993 30135 67051 30141
rect 67082 30132 67088 30184
rect 67140 30172 67146 30184
rect 67177 30175 67235 30181
rect 67177 30172 67189 30175
rect 67140 30144 67189 30172
rect 67140 30132 67146 30144
rect 67177 30141 67189 30144
rect 67223 30172 67235 30175
rect 67560 30172 67588 30212
rect 68649 30209 68661 30212
rect 68695 30209 68707 30243
rect 73154 30240 73160 30252
rect 68649 30203 68707 30209
rect 68940 30212 73160 30240
rect 67223 30144 67588 30172
rect 68557 30175 68615 30181
rect 67223 30141 67235 30144
rect 67177 30135 67235 30141
rect 68557 30141 68569 30175
rect 68603 30172 68615 30175
rect 68830 30172 68836 30184
rect 68603 30144 68836 30172
rect 68603 30141 68615 30144
rect 68557 30135 68615 30141
rect 68830 30132 68836 30144
rect 68888 30132 68894 30184
rect 68940 30104 68968 30212
rect 73154 30200 73160 30212
rect 73212 30200 73218 30252
rect 86586 30240 86592 30252
rect 86328 30212 86592 30240
rect 74350 30172 74356 30184
rect 74311 30144 74356 30172
rect 74350 30132 74356 30144
rect 74408 30132 74414 30184
rect 79781 30175 79839 30181
rect 79781 30141 79793 30175
rect 79827 30141 79839 30175
rect 80054 30172 80060 30184
rect 80015 30144 80060 30172
rect 79781 30135 79839 30141
rect 60884 30076 61056 30104
rect 61120 30076 68968 30104
rect 60884 30064 60890 30076
rect 61120 30036 61148 30076
rect 75914 30064 75920 30116
rect 75972 30104 75978 30116
rect 79505 30107 79563 30113
rect 79505 30104 79517 30107
rect 75972 30076 79517 30104
rect 75972 30064 75978 30076
rect 79505 30073 79517 30076
rect 79551 30104 79563 30107
rect 79796 30104 79824 30135
rect 80054 30132 80060 30144
rect 80112 30132 80118 30184
rect 84289 30175 84347 30181
rect 84289 30141 84301 30175
rect 84335 30172 84347 30175
rect 84654 30172 84660 30184
rect 84335 30144 84660 30172
rect 84335 30141 84347 30144
rect 84289 30135 84347 30141
rect 84654 30132 84660 30144
rect 84712 30132 84718 30184
rect 85390 30132 85396 30184
rect 85448 30172 85454 30184
rect 86328 30181 86356 30212
rect 86586 30200 86592 30212
rect 86644 30240 86650 30252
rect 87693 30243 87751 30249
rect 87693 30240 87705 30243
rect 86644 30212 87705 30240
rect 86644 30200 86650 30212
rect 87693 30209 87705 30212
rect 87739 30209 87751 30243
rect 87693 30203 87751 30209
rect 86129 30175 86187 30181
rect 86129 30172 86141 30175
rect 85448 30144 86141 30172
rect 85448 30132 85454 30144
rect 86129 30141 86141 30144
rect 86175 30141 86187 30175
rect 86129 30135 86187 30141
rect 86313 30175 86371 30181
rect 86313 30141 86325 30175
rect 86359 30141 86371 30175
rect 86678 30172 86684 30184
rect 86639 30144 86684 30172
rect 86313 30135 86371 30141
rect 86678 30132 86684 30144
rect 86736 30132 86742 30184
rect 87601 30175 87659 30181
rect 87601 30141 87613 30175
rect 87647 30172 87659 30175
rect 88242 30172 88248 30184
rect 87647 30144 88248 30172
rect 87647 30141 87659 30144
rect 87601 30135 87659 30141
rect 88242 30132 88248 30144
rect 88300 30132 88306 30184
rect 86954 30104 86960 30116
rect 79551 30076 79824 30104
rect 86915 30076 86960 30104
rect 79551 30073 79563 30076
rect 79505 30067 79563 30073
rect 86954 30064 86960 30076
rect 87012 30064 87018 30116
rect 66070 30036 66076 30048
rect 60752 30008 61148 30036
rect 66031 30008 66076 30036
rect 66070 29996 66076 30008
rect 66128 29996 66134 30048
rect 67453 30039 67511 30045
rect 67453 30005 67465 30039
rect 67499 30036 67511 30039
rect 67910 30036 67916 30048
rect 67499 30008 67916 30036
rect 67499 30005 67511 30008
rect 67453 29999 67511 30005
rect 67910 29996 67916 30008
rect 67968 29996 67974 30048
rect 68830 30036 68836 30048
rect 68791 30008 68836 30036
rect 68830 29996 68836 30008
rect 68888 29996 68894 30048
rect 73154 29996 73160 30048
rect 73212 30036 73218 30048
rect 74445 30039 74503 30045
rect 74445 30036 74457 30039
rect 73212 30008 74457 30036
rect 73212 29996 73218 30008
rect 74445 30005 74457 30008
rect 74491 30005 74503 30039
rect 74445 29999 74503 30005
rect 80514 29996 80520 30048
rect 80572 30036 80578 30048
rect 81161 30039 81219 30045
rect 81161 30036 81173 30039
rect 80572 30008 81173 30036
rect 80572 29996 80578 30008
rect 81161 30005 81173 30008
rect 81207 30005 81219 30039
rect 87046 30036 87052 30048
rect 87007 30008 87052 30036
rect 81161 29999 81219 30005
rect 87046 29996 87052 30008
rect 87104 29996 87110 30048
rect 1104 29946 108008 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 50326 29946
rect 50378 29894 50390 29946
rect 50442 29894 50454 29946
rect 50506 29894 50518 29946
rect 50570 29894 81046 29946
rect 81098 29894 81110 29946
rect 81162 29894 81174 29946
rect 81226 29894 81238 29946
rect 81290 29894 108008 29946
rect 1104 29872 108008 29894
rect 4430 29792 4436 29844
rect 4488 29832 4494 29844
rect 13446 29832 13452 29844
rect 4488 29804 13452 29832
rect 4488 29792 4494 29804
rect 13446 29792 13452 29804
rect 13504 29792 13510 29844
rect 15378 29792 15384 29844
rect 15436 29832 15442 29844
rect 15473 29835 15531 29841
rect 15473 29832 15485 29835
rect 15436 29804 15485 29832
rect 15436 29792 15442 29804
rect 15473 29801 15485 29804
rect 15519 29801 15531 29835
rect 17954 29832 17960 29844
rect 17915 29804 17960 29832
rect 15473 29795 15531 29801
rect 17954 29792 17960 29804
rect 18012 29792 18018 29844
rect 18230 29792 18236 29844
rect 18288 29832 18294 29844
rect 19242 29832 19248 29844
rect 18288 29804 19248 29832
rect 18288 29792 18294 29804
rect 19242 29792 19248 29804
rect 19300 29832 19306 29844
rect 19337 29835 19395 29841
rect 19337 29832 19349 29835
rect 19300 29804 19349 29832
rect 19300 29792 19306 29804
rect 19337 29801 19349 29804
rect 19383 29801 19395 29835
rect 19337 29795 19395 29801
rect 27154 29792 27160 29844
rect 27212 29832 27218 29844
rect 27798 29832 27804 29844
rect 27212 29804 27804 29832
rect 27212 29792 27218 29804
rect 6549 29767 6607 29773
rect 6549 29733 6561 29767
rect 6595 29764 6607 29767
rect 6638 29764 6644 29776
rect 6595 29736 6644 29764
rect 6595 29733 6607 29736
rect 6549 29727 6607 29733
rect 6638 29724 6644 29736
rect 6696 29764 6702 29776
rect 7742 29764 7748 29776
rect 6696 29736 7748 29764
rect 6696 29724 6702 29736
rect 7742 29724 7748 29736
rect 7800 29724 7806 29776
rect 4706 29696 4712 29708
rect 4667 29668 4712 29696
rect 4706 29656 4712 29668
rect 4764 29656 4770 29708
rect 4985 29699 5043 29705
rect 4985 29665 4997 29699
rect 5031 29696 5043 29699
rect 8478 29696 8484 29708
rect 5031 29668 8484 29696
rect 5031 29665 5043 29668
rect 4985 29659 5043 29665
rect 8478 29656 8484 29668
rect 8536 29656 8542 29708
rect 9674 29656 9680 29708
rect 9732 29696 9738 29708
rect 9950 29696 9956 29708
rect 9732 29668 9777 29696
rect 9911 29668 9956 29696
rect 9732 29656 9738 29668
rect 9950 29656 9956 29668
rect 10008 29656 10014 29708
rect 11333 29699 11391 29705
rect 11333 29665 11345 29699
rect 11379 29696 11391 29699
rect 11882 29696 11888 29708
rect 11379 29668 11888 29696
rect 11379 29665 11391 29668
rect 11333 29659 11391 29665
rect 11882 29656 11888 29668
rect 11940 29656 11946 29708
rect 15289 29699 15347 29705
rect 15289 29665 15301 29699
rect 15335 29696 15347 29699
rect 15562 29696 15568 29708
rect 15335 29668 15568 29696
rect 15335 29665 15347 29668
rect 15289 29659 15347 29665
rect 15562 29656 15568 29668
rect 15620 29696 15626 29708
rect 16114 29696 16120 29708
rect 15620 29668 16120 29696
rect 15620 29656 15626 29668
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 17972 29696 18000 29792
rect 18322 29724 18328 29776
rect 18380 29764 18386 29776
rect 23658 29764 23664 29776
rect 18380 29736 23664 29764
rect 18380 29724 18386 29736
rect 23658 29724 23664 29736
rect 23716 29724 23722 29776
rect 26786 29764 26792 29776
rect 26747 29736 26792 29764
rect 26786 29724 26792 29736
rect 26844 29764 26850 29776
rect 26844 29736 27016 29764
rect 26844 29724 26850 29736
rect 18049 29699 18107 29705
rect 18049 29696 18061 29699
rect 17972 29668 18061 29696
rect 18049 29665 18061 29668
rect 18095 29665 18107 29699
rect 18049 29659 18107 29665
rect 18141 29699 18199 29705
rect 18141 29665 18153 29699
rect 18187 29696 18199 29699
rect 19521 29699 19579 29705
rect 19521 29696 19533 29699
rect 18187 29668 19533 29696
rect 18187 29665 18199 29668
rect 18141 29659 18199 29665
rect 19521 29665 19533 29668
rect 19567 29696 19579 29699
rect 19978 29696 19984 29708
rect 19567 29668 19984 29696
rect 19567 29665 19579 29668
rect 19521 29659 19579 29665
rect 19978 29656 19984 29668
rect 20036 29656 20042 29708
rect 23845 29699 23903 29705
rect 23845 29665 23857 29699
rect 23891 29696 23903 29699
rect 24118 29696 24124 29708
rect 23891 29668 24124 29696
rect 23891 29665 23903 29668
rect 23845 29659 23903 29665
rect 24118 29656 24124 29668
rect 24176 29656 24182 29708
rect 26988 29705 27016 29736
rect 26973 29699 27031 29705
rect 26973 29665 26985 29699
rect 27019 29665 27031 29699
rect 26973 29659 27031 29665
rect 27157 29699 27215 29705
rect 27157 29665 27169 29699
rect 27203 29696 27215 29699
rect 27264 29696 27292 29804
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 28169 29835 28227 29841
rect 28169 29801 28181 29835
rect 28215 29832 28227 29835
rect 29362 29832 29368 29844
rect 28215 29804 29368 29832
rect 28215 29801 28227 29804
rect 28169 29795 28227 29801
rect 29362 29792 29368 29804
rect 29420 29792 29426 29844
rect 29822 29792 29828 29844
rect 29880 29832 29886 29844
rect 36538 29832 36544 29844
rect 29880 29804 36544 29832
rect 29880 29792 29886 29804
rect 36538 29792 36544 29804
rect 36596 29792 36602 29844
rect 36725 29835 36783 29841
rect 36725 29801 36737 29835
rect 36771 29832 36783 29835
rect 37458 29832 37464 29844
rect 36771 29804 37464 29832
rect 36771 29801 36783 29804
rect 36725 29795 36783 29801
rect 37458 29792 37464 29804
rect 37516 29792 37522 29844
rect 40954 29832 40960 29844
rect 40915 29804 40960 29832
rect 40954 29792 40960 29804
rect 41012 29792 41018 29844
rect 41782 29792 41788 29844
rect 41840 29832 41846 29844
rect 42058 29832 42064 29844
rect 41840 29804 42064 29832
rect 41840 29792 41846 29804
rect 42058 29792 42064 29804
rect 42116 29792 42122 29844
rect 42242 29832 42248 29844
rect 42203 29804 42248 29832
rect 42242 29792 42248 29804
rect 42300 29792 42306 29844
rect 42613 29835 42671 29841
rect 42613 29801 42625 29835
rect 42659 29832 42671 29835
rect 42794 29832 42800 29844
rect 42659 29804 42800 29832
rect 42659 29801 42671 29804
rect 42613 29795 42671 29801
rect 42794 29792 42800 29804
rect 42852 29832 42858 29844
rect 43438 29832 43444 29844
rect 42852 29804 43444 29832
rect 42852 29792 42858 29804
rect 43438 29792 43444 29804
rect 43496 29792 43502 29844
rect 47486 29792 47492 29844
rect 47544 29832 47550 29844
rect 52638 29832 52644 29844
rect 47544 29804 52644 29832
rect 47544 29792 47550 29804
rect 52638 29792 52644 29804
rect 52696 29792 52702 29844
rect 53006 29792 53012 29844
rect 53064 29832 53070 29844
rect 53101 29835 53159 29841
rect 53101 29832 53113 29835
rect 53064 29804 53113 29832
rect 53064 29792 53070 29804
rect 53101 29801 53113 29804
rect 53147 29801 53159 29835
rect 60550 29832 60556 29844
rect 53101 29795 53159 29801
rect 54680 29804 60556 29832
rect 28445 29767 28503 29773
rect 28445 29764 28457 29767
rect 27632 29736 28457 29764
rect 27632 29705 27660 29736
rect 28445 29733 28457 29736
rect 28491 29764 28503 29767
rect 29273 29767 29331 29773
rect 29273 29764 29285 29767
rect 28491 29736 29285 29764
rect 28491 29733 28503 29736
rect 28445 29727 28503 29733
rect 29273 29733 29285 29736
rect 29319 29733 29331 29767
rect 29273 29727 29331 29733
rect 29549 29767 29607 29773
rect 29549 29733 29561 29767
rect 29595 29764 29607 29767
rect 30834 29764 30840 29776
rect 29595 29736 30840 29764
rect 29595 29733 29607 29736
rect 29549 29727 29607 29733
rect 27617 29699 27675 29705
rect 27617 29696 27629 29699
rect 27203 29668 27292 29696
rect 27356 29668 27629 29696
rect 27203 29665 27215 29668
rect 27157 29659 27215 29665
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 19300 29600 19441 29628
rect 19300 29588 19306 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 23569 29631 23627 29637
rect 23569 29628 23581 29631
rect 23523 29600 23581 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 23569 29597 23581 29600
rect 23615 29628 23627 29631
rect 24026 29628 24032 29640
rect 23615 29600 24032 29628
rect 23615 29597 23627 29600
rect 23569 29591 23627 29597
rect 24026 29588 24032 29600
rect 24084 29628 24090 29640
rect 26142 29628 26148 29640
rect 24084 29600 26148 29628
rect 24084 29588 24090 29600
rect 26142 29588 26148 29600
rect 26200 29588 26206 29640
rect 26878 29588 26884 29640
rect 26936 29628 26942 29640
rect 27356 29628 27384 29668
rect 27617 29665 27629 29668
rect 27663 29665 27675 29699
rect 27617 29659 27675 29665
rect 27709 29699 27767 29705
rect 27709 29665 27721 29699
rect 27755 29696 27767 29699
rect 27798 29696 27804 29708
rect 27755 29668 27804 29696
rect 27755 29665 27767 29668
rect 27709 29659 27767 29665
rect 27798 29656 27804 29668
rect 27856 29696 27862 29708
rect 28718 29696 28724 29708
rect 27856 29668 28724 29696
rect 27856 29656 27862 29668
rect 28718 29656 28724 29668
rect 28776 29696 28782 29708
rect 28813 29699 28871 29705
rect 28813 29696 28825 29699
rect 28776 29668 28825 29696
rect 28776 29656 28782 29668
rect 28813 29665 28825 29668
rect 28859 29665 28871 29699
rect 28813 29659 28871 29665
rect 29181 29699 29239 29705
rect 29181 29665 29193 29699
rect 29227 29696 29239 29699
rect 29564 29696 29592 29727
rect 30834 29724 30840 29736
rect 30892 29724 30898 29776
rect 35437 29767 35495 29773
rect 35437 29733 35449 29767
rect 35483 29764 35495 29767
rect 45278 29764 45284 29776
rect 35483 29736 45284 29764
rect 35483 29733 35495 29736
rect 35437 29727 35495 29733
rect 29227 29668 29592 29696
rect 35253 29699 35311 29705
rect 29227 29665 29239 29668
rect 29181 29659 29239 29665
rect 35253 29665 35265 29699
rect 35299 29696 35311 29699
rect 35452 29696 35480 29727
rect 45278 29724 45284 29736
rect 45336 29724 45342 29776
rect 45465 29767 45523 29773
rect 45465 29764 45477 29767
rect 45388 29736 45477 29764
rect 35299 29668 35480 29696
rect 36633 29699 36691 29705
rect 35299 29665 35311 29668
rect 35253 29659 35311 29665
rect 36633 29665 36645 29699
rect 36679 29696 36691 29699
rect 36909 29699 36967 29705
rect 36909 29696 36921 29699
rect 36679 29668 36921 29696
rect 36679 29665 36691 29668
rect 36633 29659 36691 29665
rect 36909 29665 36921 29668
rect 36955 29696 36967 29699
rect 36998 29696 37004 29708
rect 36955 29668 37004 29696
rect 36955 29665 36967 29668
rect 36909 29659 36967 29665
rect 26936 29600 27384 29628
rect 26936 29588 26942 29600
rect 28166 29588 28172 29640
rect 28224 29628 28230 29640
rect 36648 29628 36676 29659
rect 36998 29656 37004 29668
rect 37056 29656 37062 29708
rect 37274 29656 37280 29708
rect 37332 29696 37338 29708
rect 38286 29696 38292 29708
rect 37332 29668 38292 29696
rect 37332 29656 37338 29668
rect 38286 29656 38292 29668
rect 38344 29656 38350 29708
rect 40954 29656 40960 29708
rect 41012 29696 41018 29708
rect 41049 29699 41107 29705
rect 41049 29696 41061 29699
rect 41012 29668 41061 29696
rect 41012 29656 41018 29668
rect 41049 29665 41061 29668
rect 41095 29665 41107 29699
rect 41230 29696 41236 29708
rect 41191 29668 41236 29696
rect 41049 29659 41107 29665
rect 41230 29656 41236 29668
rect 41288 29656 41294 29708
rect 41782 29696 41788 29708
rect 41743 29668 41788 29696
rect 41782 29656 41788 29668
rect 41840 29656 41846 29708
rect 41969 29699 42027 29705
rect 41969 29665 41981 29699
rect 42015 29696 42027 29699
rect 42794 29696 42800 29708
rect 42015 29668 42800 29696
rect 42015 29665 42027 29668
rect 41969 29659 42027 29665
rect 42794 29656 42800 29668
rect 42852 29656 42858 29708
rect 44269 29699 44327 29705
rect 44269 29665 44281 29699
rect 44315 29665 44327 29699
rect 44269 29659 44327 29665
rect 28224 29600 36676 29628
rect 28224 29588 28230 29600
rect 42242 29588 42248 29640
rect 42300 29628 42306 29640
rect 42705 29631 42763 29637
rect 42705 29628 42717 29631
rect 42300 29600 42717 29628
rect 42300 29588 42306 29600
rect 42705 29597 42717 29600
rect 42751 29628 42763 29631
rect 44174 29628 44180 29640
rect 42751 29600 44180 29628
rect 42751 29597 42763 29600
rect 42705 29591 42763 29597
rect 44174 29588 44180 29600
rect 44232 29588 44238 29640
rect 44284 29628 44312 29659
rect 45388 29640 45416 29736
rect 45465 29733 45477 29736
rect 45511 29733 45523 29767
rect 45465 29727 45523 29733
rect 46842 29724 46848 29776
rect 46900 29764 46906 29776
rect 46900 29736 48360 29764
rect 46900 29724 46906 29736
rect 47026 29696 47032 29708
rect 46987 29668 47032 29696
rect 47026 29656 47032 29668
rect 47084 29656 47090 29708
rect 48225 29699 48283 29705
rect 48225 29665 48237 29699
rect 48271 29665 48283 29699
rect 48332 29696 48360 29736
rect 50982 29696 50988 29708
rect 48332 29668 50988 29696
rect 48225 29659 48283 29665
rect 44284 29600 45324 29628
rect 2774 29520 2780 29572
rect 2832 29560 2838 29572
rect 3234 29560 3240 29572
rect 2832 29532 3240 29560
rect 2832 29520 2838 29532
rect 3234 29520 3240 29532
rect 3292 29520 3298 29572
rect 17310 29520 17316 29572
rect 17368 29560 17374 29572
rect 17368 29532 18368 29560
rect 17368 29520 17374 29532
rect 4062 29452 4068 29504
rect 4120 29492 4126 29504
rect 6089 29495 6147 29501
rect 6089 29492 6101 29495
rect 4120 29464 6101 29492
rect 4120 29452 4126 29464
rect 6089 29461 6101 29464
rect 6135 29461 6147 29495
rect 6089 29455 6147 29461
rect 9493 29495 9551 29501
rect 9493 29461 9505 29495
rect 9539 29492 9551 29495
rect 9674 29492 9680 29504
rect 9539 29464 9680 29492
rect 9539 29461 9551 29464
rect 9493 29455 9551 29461
rect 9674 29452 9680 29464
rect 9732 29452 9738 29504
rect 18340 29501 18368 29532
rect 24578 29520 24584 29572
rect 24636 29560 24642 29572
rect 24636 29532 29408 29560
rect 24636 29520 24642 29532
rect 18325 29495 18383 29501
rect 18325 29461 18337 29495
rect 18371 29461 18383 29495
rect 18325 29455 18383 29461
rect 18690 29452 18696 29504
rect 18748 29492 18754 29504
rect 19705 29495 19763 29501
rect 19705 29492 19717 29495
rect 18748 29464 19717 29492
rect 18748 29452 18754 29464
rect 19705 29461 19717 29464
rect 19751 29461 19763 29495
rect 19705 29455 19763 29461
rect 24762 29452 24768 29504
rect 24820 29492 24826 29504
rect 25133 29495 25191 29501
rect 25133 29492 25145 29495
rect 24820 29464 25145 29492
rect 24820 29452 24826 29464
rect 25133 29461 25145 29464
rect 25179 29492 25191 29495
rect 26326 29492 26332 29504
rect 25179 29464 26332 29492
rect 25179 29461 25191 29464
rect 25133 29455 25191 29461
rect 26326 29452 26332 29464
rect 26384 29452 26390 29504
rect 26418 29452 26424 29504
rect 26476 29492 26482 29504
rect 29270 29492 29276 29504
rect 26476 29464 29276 29492
rect 26476 29452 26482 29464
rect 29270 29452 29276 29464
rect 29328 29452 29334 29504
rect 29380 29492 29408 29532
rect 29454 29520 29460 29572
rect 29512 29560 29518 29572
rect 40494 29560 40500 29572
rect 29512 29532 40500 29560
rect 29512 29520 29518 29532
rect 40494 29520 40500 29532
rect 40552 29520 40558 29572
rect 45296 29560 45324 29600
rect 45370 29588 45376 29640
rect 45428 29588 45434 29640
rect 45554 29588 45560 29640
rect 45612 29628 45618 29640
rect 47857 29631 47915 29637
rect 47857 29628 47869 29631
rect 45612 29600 47869 29628
rect 45612 29588 45618 29600
rect 47857 29597 47869 29600
rect 47903 29628 47915 29631
rect 48240 29628 48268 29659
rect 50982 29656 50988 29668
rect 51040 29656 51046 29708
rect 51261 29699 51319 29705
rect 51261 29665 51273 29699
rect 51307 29696 51319 29699
rect 51445 29699 51503 29705
rect 51445 29696 51457 29699
rect 51307 29668 51457 29696
rect 51307 29665 51319 29668
rect 51261 29659 51319 29665
rect 51445 29665 51457 29668
rect 51491 29696 51503 29699
rect 51629 29699 51687 29705
rect 51629 29696 51641 29699
rect 51491 29668 51641 29696
rect 51491 29665 51503 29668
rect 51445 29659 51503 29665
rect 51629 29665 51641 29668
rect 51675 29696 51687 29699
rect 52089 29699 52147 29705
rect 52089 29696 52101 29699
rect 51675 29668 52101 29696
rect 51675 29665 51687 29668
rect 51629 29659 51687 29665
rect 52089 29665 52101 29668
rect 52135 29696 52147 29699
rect 52641 29699 52699 29705
rect 52641 29696 52653 29699
rect 52135 29668 52653 29696
rect 52135 29665 52147 29668
rect 52089 29659 52147 29665
rect 52641 29665 52653 29668
rect 52687 29696 52699 29699
rect 52730 29696 52736 29708
rect 52687 29668 52736 29696
rect 52687 29665 52699 29668
rect 52641 29659 52699 29665
rect 52730 29656 52736 29668
rect 52788 29656 52794 29708
rect 52825 29699 52883 29705
rect 52825 29665 52837 29699
rect 52871 29696 52883 29699
rect 52871 29668 53052 29696
rect 52871 29665 52883 29668
rect 52825 29659 52883 29665
rect 47903 29600 48268 29628
rect 51813 29631 51871 29637
rect 47903 29597 47915 29600
rect 47857 29591 47915 29597
rect 51813 29597 51825 29631
rect 51859 29628 51871 29631
rect 51994 29628 52000 29640
rect 51859 29600 52000 29628
rect 51859 29597 51871 29600
rect 51813 29591 51871 29597
rect 51994 29588 52000 29600
rect 52052 29588 52058 29640
rect 53024 29628 53052 29668
rect 53098 29656 53104 29708
rect 53156 29696 53162 29708
rect 54680 29696 54708 29804
rect 60550 29792 60556 29804
rect 60608 29792 60614 29844
rect 67634 29792 67640 29844
rect 67692 29832 67698 29844
rect 69385 29835 69443 29841
rect 69385 29832 69397 29835
rect 67692 29804 69397 29832
rect 67692 29792 67698 29804
rect 69385 29801 69397 29804
rect 69431 29801 69443 29835
rect 69385 29795 69443 29801
rect 56413 29767 56471 29773
rect 56413 29764 56425 29767
rect 53156 29668 54708 29696
rect 55048 29736 56425 29764
rect 53156 29656 53162 29668
rect 53190 29628 53196 29640
rect 53024 29600 53196 29628
rect 53190 29588 53196 29600
rect 53248 29628 53254 29640
rect 53377 29631 53435 29637
rect 53377 29628 53389 29631
rect 53248 29600 53389 29628
rect 53248 29588 53254 29600
rect 53377 29597 53389 29600
rect 53423 29628 53435 29631
rect 54662 29628 54668 29640
rect 53423 29600 54668 29628
rect 53423 29597 53435 29600
rect 53377 29591 53435 29597
rect 54662 29588 54668 29600
rect 54720 29588 54726 29640
rect 48038 29560 48044 29572
rect 45296 29532 48044 29560
rect 48038 29520 48044 29532
rect 48096 29520 48102 29572
rect 48130 29520 48136 29572
rect 48188 29560 48194 29572
rect 55048 29560 55076 29736
rect 56413 29733 56425 29736
rect 56459 29764 56471 29767
rect 56597 29767 56655 29773
rect 56597 29764 56609 29767
rect 56459 29736 56609 29764
rect 56459 29733 56471 29736
rect 56413 29727 56471 29733
rect 56597 29733 56609 29736
rect 56643 29764 56655 29767
rect 58253 29767 58311 29773
rect 56643 29736 57192 29764
rect 56643 29733 56655 29736
rect 56597 29727 56655 29733
rect 55125 29699 55183 29705
rect 55125 29665 55137 29699
rect 55171 29696 55183 29699
rect 55490 29696 55496 29708
rect 55171 29668 55496 29696
rect 55171 29665 55183 29668
rect 55125 29659 55183 29665
rect 55490 29656 55496 29668
rect 55548 29656 55554 29708
rect 56778 29696 56784 29708
rect 56739 29668 56784 29696
rect 56778 29656 56784 29668
rect 56836 29696 56842 29708
rect 57164 29705 57192 29736
rect 58253 29733 58265 29767
rect 58299 29764 58311 29767
rect 58299 29736 60320 29764
rect 58299 29733 58311 29736
rect 58253 29727 58311 29733
rect 56965 29699 57023 29705
rect 56965 29696 56977 29699
rect 56836 29668 56977 29696
rect 56836 29656 56842 29668
rect 56965 29665 56977 29668
rect 57011 29665 57023 29699
rect 56965 29659 57023 29665
rect 57149 29699 57207 29705
rect 57149 29665 57161 29699
rect 57195 29696 57207 29699
rect 57701 29699 57759 29705
rect 57701 29696 57713 29699
rect 57195 29668 57713 29696
rect 57195 29665 57207 29668
rect 57149 29659 57207 29665
rect 57701 29665 57713 29668
rect 57747 29665 57759 29699
rect 57882 29696 57888 29708
rect 57843 29668 57888 29696
rect 57701 29659 57759 29665
rect 57882 29656 57888 29668
rect 57940 29696 57946 29708
rect 58434 29696 58440 29708
rect 57940 29668 58440 29696
rect 57940 29656 57946 29668
rect 58434 29656 58440 29668
rect 58492 29656 58498 29708
rect 60292 29696 60320 29736
rect 61286 29724 61292 29776
rect 61344 29764 61350 29776
rect 61933 29767 61991 29773
rect 61933 29764 61945 29767
rect 61344 29736 61945 29764
rect 61344 29724 61350 29736
rect 61933 29733 61945 29736
rect 61979 29733 61991 29767
rect 61933 29727 61991 29733
rect 60461 29699 60519 29705
rect 60461 29696 60473 29699
rect 60292 29668 60473 29696
rect 60461 29665 60473 29668
rect 60507 29665 60519 29699
rect 60461 29659 60519 29665
rect 60550 29656 60556 29708
rect 60608 29696 60614 29708
rect 67910 29696 67916 29708
rect 60608 29668 67772 29696
rect 67871 29668 67916 29696
rect 60608 29656 60614 29668
rect 59449 29631 59507 29637
rect 59449 29597 59461 29631
rect 59495 29628 59507 29631
rect 59630 29628 59636 29640
rect 59495 29600 59636 29628
rect 59495 29597 59507 29600
rect 59449 29591 59507 29597
rect 59630 29588 59636 29600
rect 59688 29588 59694 29640
rect 60182 29628 60188 29640
rect 60143 29600 60188 29628
rect 60182 29588 60188 29600
rect 60240 29588 60246 29640
rect 67634 29628 67640 29640
rect 67595 29600 67640 29628
rect 67634 29588 67640 29600
rect 67692 29588 67698 29640
rect 67744 29628 67772 29668
rect 67910 29656 67916 29668
rect 67968 29656 67974 29708
rect 69400 29696 69428 29795
rect 69474 29792 69480 29844
rect 69532 29832 69538 29844
rect 73154 29832 73160 29844
rect 69532 29804 73160 29832
rect 69532 29792 69538 29804
rect 72528 29705 72556 29804
rect 73154 29792 73160 29804
rect 73212 29792 73218 29844
rect 74350 29792 74356 29844
rect 74408 29832 74414 29844
rect 75181 29835 75239 29841
rect 75181 29832 75193 29835
rect 74408 29804 75193 29832
rect 74408 29792 74414 29804
rect 75181 29801 75193 29804
rect 75227 29801 75239 29835
rect 75181 29795 75239 29801
rect 79321 29835 79379 29841
rect 79321 29801 79333 29835
rect 79367 29832 79379 29835
rect 80054 29832 80060 29844
rect 79367 29804 80060 29832
rect 79367 29801 79379 29804
rect 79321 29795 79379 29801
rect 80054 29792 80060 29804
rect 80112 29792 80118 29844
rect 80609 29835 80667 29841
rect 80609 29801 80621 29835
rect 80655 29832 80667 29835
rect 80698 29832 80704 29844
rect 80655 29804 80704 29832
rect 80655 29801 80667 29804
rect 80609 29795 80667 29801
rect 80698 29792 80704 29804
rect 80756 29792 80762 29844
rect 72881 29767 72939 29773
rect 72881 29733 72893 29767
rect 72927 29733 72939 29767
rect 72881 29727 72939 29733
rect 71225 29699 71283 29705
rect 71225 29696 71237 29699
rect 69400 29668 71237 29696
rect 71225 29665 71237 29668
rect 71271 29665 71283 29699
rect 71777 29699 71835 29705
rect 71777 29696 71789 29699
rect 71225 29659 71283 29665
rect 71424 29668 71789 29696
rect 71424 29637 71452 29668
rect 71777 29665 71789 29668
rect 71823 29696 71835 29699
rect 72329 29699 72387 29705
rect 72329 29696 72341 29699
rect 71823 29668 72341 29696
rect 71823 29665 71835 29668
rect 71777 29659 71835 29665
rect 72329 29665 72341 29668
rect 72375 29665 72387 29699
rect 72329 29659 72387 29665
rect 72513 29699 72571 29705
rect 72513 29665 72525 29699
rect 72559 29665 72571 29699
rect 72896 29696 72924 29727
rect 74077 29699 74135 29705
rect 74077 29696 74089 29699
rect 72896 29668 74089 29696
rect 72513 29659 72571 29665
rect 74077 29665 74089 29668
rect 74123 29665 74135 29699
rect 79226 29696 79232 29708
rect 79187 29668 79232 29696
rect 74077 29659 74135 29665
rect 79226 29656 79232 29668
rect 79284 29656 79290 29708
rect 80514 29696 80520 29708
rect 80475 29668 80520 29696
rect 80514 29656 80520 29668
rect 80572 29656 80578 29708
rect 71041 29631 71099 29637
rect 71041 29628 71053 29631
rect 67744 29600 71053 29628
rect 71041 29597 71053 29600
rect 71087 29628 71099 29631
rect 71409 29631 71467 29637
rect 71409 29628 71421 29631
rect 71087 29600 71421 29628
rect 71087 29597 71099 29600
rect 71041 29591 71099 29597
rect 71409 29597 71421 29600
rect 71455 29597 71467 29631
rect 71590 29628 71596 29640
rect 71551 29600 71596 29628
rect 71409 29591 71467 29597
rect 71590 29588 71596 29600
rect 71648 29588 71654 29640
rect 73801 29631 73859 29637
rect 73801 29597 73813 29631
rect 73847 29628 73859 29631
rect 75549 29631 75607 29637
rect 75549 29628 75561 29631
rect 73847 29600 75561 29628
rect 73847 29597 73859 29600
rect 73801 29591 73859 29597
rect 75549 29597 75561 29600
rect 75595 29628 75607 29631
rect 75914 29628 75920 29640
rect 75595 29600 75920 29628
rect 75595 29597 75607 29600
rect 75549 29591 75607 29597
rect 48188 29532 55076 29560
rect 48188 29520 48194 29532
rect 55306 29520 55312 29572
rect 55364 29560 55370 29572
rect 59078 29560 59084 29572
rect 55364 29532 55409 29560
rect 59039 29532 59084 29560
rect 55364 29520 55370 29532
rect 59078 29520 59084 29532
rect 59136 29520 59142 29572
rect 59538 29560 59544 29572
rect 59499 29532 59544 29560
rect 59538 29520 59544 29532
rect 59596 29520 59602 29572
rect 35069 29495 35127 29501
rect 35069 29492 35081 29495
rect 29380 29464 35081 29492
rect 35069 29461 35081 29464
rect 35115 29461 35127 29495
rect 35069 29455 35127 29461
rect 35894 29452 35900 29504
rect 35952 29492 35958 29504
rect 41598 29492 41604 29504
rect 35952 29464 41604 29492
rect 35952 29452 35958 29464
rect 41598 29452 41604 29464
rect 41656 29492 41662 29504
rect 43346 29492 43352 29504
rect 41656 29464 43352 29492
rect 41656 29452 41662 29464
rect 43346 29452 43352 29464
rect 43404 29492 43410 29504
rect 44085 29495 44143 29501
rect 44085 29492 44097 29495
rect 43404 29464 44097 29492
rect 43404 29452 43410 29464
rect 44085 29461 44097 29464
rect 44131 29461 44143 29495
rect 45370 29492 45376 29504
rect 45331 29464 45376 29492
rect 44085 29455 44143 29461
rect 45370 29452 45376 29464
rect 45428 29452 45434 29504
rect 46198 29452 46204 29504
rect 46256 29492 46262 29504
rect 48866 29492 48872 29504
rect 46256 29464 48872 29492
rect 46256 29452 46262 29464
rect 48866 29452 48872 29464
rect 48924 29452 48930 29504
rect 48958 29452 48964 29504
rect 49016 29492 49022 29504
rect 51261 29495 51319 29501
rect 51261 29492 51273 29495
rect 49016 29464 51273 29492
rect 49016 29452 49022 29464
rect 51261 29461 51273 29464
rect 51307 29461 51319 29495
rect 51261 29455 51319 29461
rect 53558 29452 53564 29504
rect 53616 29492 53622 29504
rect 58710 29492 58716 29504
rect 53616 29464 58716 29492
rect 53616 29452 53622 29464
rect 58710 29452 58716 29464
rect 58768 29452 58774 29504
rect 58897 29495 58955 29501
rect 58897 29461 58909 29495
rect 58943 29492 58955 29495
rect 58986 29492 58992 29504
rect 58943 29464 58992 29492
rect 58943 29461 58955 29464
rect 58897 29455 58955 29461
rect 58986 29452 58992 29464
rect 59044 29452 59050 29504
rect 59170 29492 59176 29504
rect 59131 29464 59176 29492
rect 59170 29452 59176 29464
rect 59228 29452 59234 29504
rect 59722 29492 59728 29504
rect 59683 29464 59728 29492
rect 59722 29452 59728 29464
rect 59780 29452 59786 29504
rect 59906 29492 59912 29504
rect 59867 29464 59912 29492
rect 59906 29452 59912 29464
rect 59964 29452 59970 29504
rect 60200 29492 60228 29588
rect 71225 29563 71283 29569
rect 71225 29529 71237 29563
rect 71271 29560 71283 29563
rect 73816 29560 73844 29591
rect 75914 29588 75920 29600
rect 75972 29588 75978 29640
rect 71271 29532 73844 29560
rect 71271 29529 71283 29532
rect 71225 29523 71283 29529
rect 82906 29520 82912 29572
rect 82964 29560 82970 29572
rect 83918 29560 83924 29572
rect 82964 29532 83924 29560
rect 82964 29520 82970 29532
rect 83918 29520 83924 29532
rect 83976 29560 83982 29572
rect 86865 29563 86923 29569
rect 86865 29560 86877 29563
rect 83976 29532 86877 29560
rect 83976 29520 83982 29532
rect 86865 29529 86877 29532
rect 86911 29529 86923 29563
rect 87138 29560 87144 29572
rect 87099 29532 87144 29560
rect 86865 29523 86923 29529
rect 87138 29520 87144 29532
rect 87196 29520 87202 29572
rect 61286 29492 61292 29504
rect 60200 29464 61292 29492
rect 61286 29452 61292 29464
rect 61344 29452 61350 29504
rect 61562 29492 61568 29504
rect 61523 29464 61568 29492
rect 61562 29452 61568 29464
rect 61620 29452 61626 29504
rect 67910 29452 67916 29504
rect 67968 29492 67974 29504
rect 68830 29492 68836 29504
rect 67968 29464 68836 29492
rect 67968 29452 67974 29464
rect 68830 29452 68836 29464
rect 68888 29492 68894 29504
rect 69017 29495 69075 29501
rect 69017 29492 69029 29495
rect 68888 29464 69029 29492
rect 68888 29452 68894 29464
rect 69017 29461 69029 29464
rect 69063 29461 69075 29495
rect 86310 29492 86316 29504
rect 86271 29464 86316 29492
rect 69017 29455 69075 29461
rect 86310 29452 86316 29464
rect 86368 29452 86374 29504
rect 86494 29492 86500 29504
rect 86455 29464 86500 29492
rect 86494 29452 86500 29464
rect 86552 29452 86558 29504
rect 86586 29452 86592 29504
rect 86644 29492 86650 29504
rect 86681 29495 86739 29501
rect 86681 29492 86693 29495
rect 86644 29464 86693 29492
rect 86644 29452 86650 29464
rect 86681 29461 86693 29464
rect 86727 29461 86739 29495
rect 87230 29492 87236 29504
rect 87191 29464 87236 29492
rect 86681 29455 86739 29461
rect 87230 29452 87236 29464
rect 87288 29452 87294 29504
rect 87414 29492 87420 29504
rect 87375 29464 87420 29492
rect 87414 29452 87420 29464
rect 87472 29452 87478 29504
rect 87598 29492 87604 29504
rect 87559 29464 87604 29492
rect 87598 29452 87604 29464
rect 87656 29452 87662 29504
rect 1104 29402 108008 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 65686 29402
rect 65738 29350 65750 29402
rect 65802 29350 65814 29402
rect 65866 29350 65878 29402
rect 65930 29350 96406 29402
rect 96458 29350 96470 29402
rect 96522 29350 96534 29402
rect 96586 29350 96598 29402
rect 96650 29350 108008 29402
rect 1104 29328 108008 29350
rect 4617 29291 4675 29297
rect 4617 29288 4629 29291
rect 2792 29260 4629 29288
rect 2590 29112 2596 29164
rect 2648 29152 2654 29164
rect 2792 29161 2820 29260
rect 4617 29257 4629 29260
rect 4663 29288 4675 29291
rect 4706 29288 4712 29300
rect 4663 29260 4712 29288
rect 4663 29257 4675 29260
rect 4617 29251 4675 29257
rect 4706 29248 4712 29260
rect 4764 29288 4770 29300
rect 4890 29288 4896 29300
rect 4764 29260 4896 29288
rect 4764 29248 4770 29260
rect 4890 29248 4896 29260
rect 4948 29248 4954 29300
rect 13173 29291 13231 29297
rect 13173 29257 13185 29291
rect 13219 29288 13231 29291
rect 23014 29288 23020 29300
rect 13219 29260 23020 29288
rect 13219 29257 13231 29260
rect 13173 29251 13231 29257
rect 2777 29155 2835 29161
rect 2777 29152 2789 29155
rect 2648 29124 2789 29152
rect 2648 29112 2654 29124
rect 2777 29121 2789 29124
rect 2823 29121 2835 29155
rect 3050 29152 3056 29164
rect 3011 29124 3056 29152
rect 2777 29115 2835 29121
rect 3050 29112 3056 29124
rect 3108 29112 3114 29164
rect 3418 29112 3424 29164
rect 3476 29152 3482 29164
rect 4157 29155 4215 29161
rect 4157 29152 4169 29155
rect 3476 29124 4169 29152
rect 3476 29112 3482 29124
rect 4157 29121 4169 29124
rect 4203 29121 4215 29155
rect 4157 29115 4215 29121
rect 11882 29112 11888 29164
rect 11940 29152 11946 29164
rect 12437 29155 12495 29161
rect 12437 29152 12449 29155
rect 11940 29124 12449 29152
rect 11940 29112 11946 29124
rect 12437 29121 12449 29124
rect 12483 29152 12495 29155
rect 13188 29152 13216 29251
rect 23014 29248 23020 29260
rect 23072 29248 23078 29300
rect 23106 29248 23112 29300
rect 23164 29288 23170 29300
rect 46198 29288 46204 29300
rect 23164 29260 46204 29288
rect 23164 29248 23170 29260
rect 46198 29248 46204 29260
rect 46256 29248 46262 29300
rect 47026 29248 47032 29300
rect 47084 29288 47090 29300
rect 55490 29288 55496 29300
rect 47084 29260 55496 29288
rect 47084 29248 47090 29260
rect 55490 29248 55496 29260
rect 55548 29248 55554 29300
rect 56778 29248 56784 29300
rect 56836 29288 56842 29300
rect 66070 29288 66076 29300
rect 56836 29260 66076 29288
rect 56836 29248 56842 29260
rect 66070 29248 66076 29260
rect 66128 29248 66134 29300
rect 20898 29220 20904 29232
rect 15396 29192 20904 29220
rect 15396 29161 15424 29192
rect 20898 29180 20904 29192
rect 20956 29180 20962 29232
rect 21361 29223 21419 29229
rect 21361 29220 21373 29223
rect 21008 29192 21373 29220
rect 12483 29124 13216 29152
rect 15381 29155 15439 29161
rect 12483 29121 12495 29124
rect 12437 29115 12495 29121
rect 15381 29121 15393 29155
rect 15427 29121 15439 29155
rect 15381 29115 15439 29121
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29152 20499 29155
rect 20487 29124 20668 29152
rect 20487 29121 20499 29124
rect 20441 29115 20499 29121
rect 12342 29044 12348 29096
rect 12400 29084 12406 29096
rect 12529 29087 12587 29093
rect 12529 29084 12541 29087
rect 12400 29056 12541 29084
rect 12400 29044 12406 29056
rect 12529 29053 12541 29056
rect 12575 29053 12587 29087
rect 12529 29047 12587 29053
rect 14553 29087 14611 29093
rect 14553 29053 14565 29087
rect 14599 29084 14611 29087
rect 14918 29084 14924 29096
rect 14599 29056 14924 29084
rect 14599 29053 14611 29056
rect 14553 29047 14611 29053
rect 14918 29044 14924 29056
rect 14976 29084 14982 29096
rect 14976 29056 15056 29084
rect 14976 29044 14982 29056
rect 12989 29019 13047 29025
rect 12989 28985 13001 29019
rect 13035 29016 13047 29019
rect 13262 29016 13268 29028
rect 13035 28988 13268 29016
rect 13035 28985 13047 28988
rect 12989 28979 13047 28985
rect 13262 28976 13268 28988
rect 13320 28976 13326 29028
rect 13998 28976 14004 29028
rect 14056 29016 14062 29028
rect 15028 29025 15056 29056
rect 16574 29044 16580 29096
rect 16632 29084 16638 29096
rect 19334 29084 19340 29096
rect 16632 29056 19340 29084
rect 16632 29044 16638 29056
rect 19334 29044 19340 29056
rect 19392 29044 19398 29096
rect 20349 29087 20407 29093
rect 20349 29053 20361 29087
rect 20395 29084 20407 29087
rect 20553 29087 20611 29093
rect 20395 29056 20484 29084
rect 20395 29053 20407 29056
rect 20349 29047 20407 29053
rect 20456 29028 20484 29056
rect 20553 29053 20565 29087
rect 20599 29053 20611 29087
rect 20640 29084 20668 29124
rect 20714 29112 20720 29164
rect 20772 29152 20778 29164
rect 21008 29152 21036 29192
rect 21361 29189 21373 29192
rect 21407 29220 21419 29223
rect 24578 29220 24584 29232
rect 21407 29192 24584 29220
rect 21407 29189 21419 29192
rect 21361 29183 21419 29189
rect 24578 29180 24584 29192
rect 24636 29180 24642 29232
rect 25038 29180 25044 29232
rect 25096 29220 25102 29232
rect 25314 29220 25320 29232
rect 25096 29192 25320 29220
rect 25096 29180 25102 29192
rect 25314 29180 25320 29192
rect 25372 29180 25378 29232
rect 25498 29180 25504 29232
rect 25556 29220 25562 29232
rect 51994 29220 52000 29232
rect 25556 29192 52000 29220
rect 25556 29180 25562 29192
rect 51994 29180 52000 29192
rect 52052 29180 52058 29232
rect 52638 29180 52644 29232
rect 52696 29220 52702 29232
rect 59998 29220 60004 29232
rect 52696 29192 60004 29220
rect 52696 29180 52702 29192
rect 59998 29180 60004 29192
rect 60056 29180 60062 29232
rect 63494 29180 63500 29232
rect 63552 29220 63558 29232
rect 69474 29220 69480 29232
rect 63552 29192 69480 29220
rect 63552 29180 63558 29192
rect 69474 29180 69480 29192
rect 69532 29180 69538 29232
rect 20772 29124 21036 29152
rect 21177 29155 21235 29161
rect 20772 29112 20778 29124
rect 21177 29121 21189 29155
rect 21223 29152 21235 29155
rect 21223 29124 25360 29152
rect 21223 29121 21235 29124
rect 21177 29115 21235 29121
rect 21192 29084 21220 29115
rect 20640 29056 21220 29084
rect 23661 29087 23719 29093
rect 20553 29047 20611 29053
rect 23661 29053 23673 29087
rect 23707 29084 23719 29087
rect 25038 29084 25044 29096
rect 23707 29056 25044 29084
rect 23707 29053 23719 29056
rect 23661 29047 23719 29053
rect 14645 29019 14703 29025
rect 14645 29016 14657 29019
rect 14056 28988 14657 29016
rect 14056 28976 14062 28988
rect 14645 28985 14657 28988
rect 14691 28985 14703 29019
rect 14645 28979 14703 28985
rect 15013 29019 15071 29025
rect 15013 28985 15025 29019
rect 15059 28985 15071 29019
rect 15013 28979 15071 28985
rect 17494 28976 17500 29028
rect 17552 29016 17558 29028
rect 17552 28988 19932 29016
rect 17552 28976 17558 28988
rect 14826 28948 14832 28960
rect 14787 28920 14832 28948
rect 14826 28908 14832 28920
rect 14884 28908 14890 28960
rect 14918 28908 14924 28960
rect 14976 28948 14982 28960
rect 19904 28948 19932 28988
rect 20438 28976 20444 29028
rect 20496 28976 20502 29028
rect 20165 28951 20223 28957
rect 20165 28948 20177 28951
rect 14976 28920 15021 28948
rect 19904 28920 20177 28948
rect 14976 28908 14982 28920
rect 20165 28917 20177 28920
rect 20211 28917 20223 28951
rect 20568 28948 20596 29047
rect 25038 29044 25044 29056
rect 25096 29044 25102 29096
rect 25130 29044 25136 29096
rect 25188 29084 25194 29096
rect 25188 29044 25222 29084
rect 20898 28976 20904 29028
rect 20956 29016 20962 29028
rect 20993 29019 21051 29025
rect 20993 29016 21005 29019
rect 20956 28988 21005 29016
rect 20956 28976 20962 28988
rect 20993 28985 21005 28988
rect 21039 28985 21051 29019
rect 20993 28979 21051 28985
rect 20806 28948 20812 28960
rect 20568 28920 20812 28948
rect 20165 28911 20223 28917
rect 20806 28908 20812 28920
rect 20864 28908 20870 28960
rect 23290 28908 23296 28960
rect 23348 28948 23354 28960
rect 23845 28951 23903 28957
rect 23845 28948 23857 28951
rect 23348 28920 23857 28948
rect 23348 28908 23354 28920
rect 23845 28917 23857 28920
rect 23891 28917 23903 28951
rect 23845 28911 23903 28917
rect 23934 28908 23940 28960
rect 23992 28948 23998 28960
rect 25194 28948 25222 29044
rect 25332 29016 25360 29124
rect 25590 29112 25596 29164
rect 25648 29152 25654 29164
rect 25648 29124 33824 29152
rect 25648 29112 25654 29124
rect 25406 29044 25412 29096
rect 25464 29084 25470 29096
rect 29454 29084 29460 29096
rect 25464 29056 29460 29084
rect 25464 29044 25470 29056
rect 29454 29044 29460 29056
rect 29512 29044 29518 29096
rect 33796 29084 33824 29124
rect 35434 29112 35440 29164
rect 35492 29152 35498 29164
rect 42794 29152 42800 29164
rect 35492 29124 42800 29152
rect 35492 29112 35498 29124
rect 42794 29112 42800 29124
rect 42852 29112 42858 29164
rect 45370 29112 45376 29164
rect 45428 29152 45434 29164
rect 53834 29152 53840 29164
rect 45428 29124 53840 29152
rect 45428 29112 45434 29124
rect 53834 29112 53840 29124
rect 53892 29112 53898 29164
rect 59262 29112 59268 29164
rect 59320 29152 59326 29164
rect 61562 29152 61568 29164
rect 59320 29124 61568 29152
rect 59320 29112 59326 29124
rect 61562 29112 61568 29124
rect 61620 29112 61626 29164
rect 73614 29152 73620 29164
rect 67652 29124 73620 29152
rect 67652 29084 67680 29124
rect 73614 29112 73620 29124
rect 73672 29112 73678 29164
rect 33796 29056 67680 29084
rect 25332 28988 50936 29016
rect 23992 28920 25222 28948
rect 50908 28948 50936 28988
rect 50982 28976 50988 29028
rect 51040 29016 51046 29028
rect 57790 29016 57796 29028
rect 51040 28988 57796 29016
rect 51040 28976 51046 28988
rect 57790 28976 57796 28988
rect 57848 29016 57854 29028
rect 59722 29016 59728 29028
rect 57848 28988 59728 29016
rect 57848 28976 57854 28988
rect 59722 28976 59728 28988
rect 59780 28976 59786 29028
rect 53558 28948 53564 28960
rect 50908 28920 53564 28948
rect 23992 28908 23998 28920
rect 53558 28908 53564 28920
rect 53616 28908 53622 28960
rect 1104 28858 29256 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 29256 28858
rect 1104 28784 29256 28806
rect 4525 28747 4583 28753
rect 4525 28713 4537 28747
rect 4571 28744 4583 28747
rect 4614 28744 4620 28756
rect 4571 28716 4620 28744
rect 4571 28713 4583 28716
rect 4525 28707 4583 28713
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 9582 28704 9588 28756
rect 9640 28744 9646 28756
rect 13541 28747 13599 28753
rect 13541 28744 13553 28747
rect 9640 28716 13553 28744
rect 9640 28704 9646 28716
rect 13541 28713 13553 28716
rect 13587 28713 13599 28747
rect 15102 28744 15108 28756
rect 13541 28707 13599 28713
rect 13740 28716 15108 28744
rect 3970 28636 3976 28688
rect 4028 28676 4034 28688
rect 13740 28676 13768 28716
rect 15102 28704 15108 28716
rect 15160 28704 15166 28756
rect 15378 28744 15384 28756
rect 15339 28716 15384 28744
rect 15378 28704 15384 28716
rect 15436 28744 15442 28756
rect 15436 28716 15976 28744
rect 15436 28704 15442 28716
rect 15948 28685 15976 28716
rect 19334 28704 19340 28756
rect 19392 28744 19398 28756
rect 20898 28744 20904 28756
rect 19392 28716 20904 28744
rect 19392 28704 19398 28716
rect 20898 28704 20904 28716
rect 20956 28704 20962 28756
rect 4028 28648 13768 28676
rect 14001 28679 14059 28685
rect 4028 28636 4034 28648
rect 14001 28645 14013 28679
rect 14047 28676 14059 28679
rect 15289 28679 15347 28685
rect 14047 28648 14596 28676
rect 14047 28645 14059 28648
rect 14001 28639 14059 28645
rect 4065 28611 4123 28617
rect 4065 28577 4077 28611
rect 4111 28608 4123 28611
rect 4614 28608 4620 28620
rect 4111 28580 4620 28608
rect 4111 28577 4123 28580
rect 4065 28571 4123 28577
rect 4614 28568 4620 28580
rect 4672 28568 4678 28620
rect 8205 28611 8263 28617
rect 8205 28577 8217 28611
rect 8251 28577 8263 28611
rect 8205 28571 8263 28577
rect 2958 28500 2964 28552
rect 3016 28540 3022 28552
rect 5074 28540 5080 28552
rect 3016 28512 5080 28540
rect 3016 28500 3022 28512
rect 5074 28500 5080 28512
rect 5132 28500 5138 28552
rect 8220 28484 8248 28571
rect 8294 28568 8300 28620
rect 8352 28608 8358 28620
rect 9677 28611 9735 28617
rect 9677 28608 9689 28611
rect 8352 28580 9689 28608
rect 8352 28568 8358 28580
rect 9677 28577 9689 28580
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 10686 28568 10692 28620
rect 10744 28608 10750 28620
rect 11241 28611 11299 28617
rect 11241 28608 11253 28611
rect 10744 28580 11253 28608
rect 10744 28568 10750 28580
rect 11241 28577 11253 28580
rect 11287 28577 11299 28611
rect 13814 28608 13820 28620
rect 13775 28580 13820 28608
rect 11241 28571 11299 28577
rect 13814 28568 13820 28580
rect 13872 28568 13878 28620
rect 13906 28568 13912 28620
rect 13964 28608 13970 28620
rect 13964 28580 14009 28608
rect 13964 28568 13970 28580
rect 13633 28543 13691 28549
rect 13633 28509 13645 28543
rect 13679 28540 13691 28543
rect 13998 28540 14004 28552
rect 13679 28512 14004 28540
rect 13679 28509 13691 28512
rect 13633 28503 13691 28509
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 14090 28500 14096 28552
rect 14148 28540 14154 28552
rect 14369 28543 14427 28549
rect 14369 28540 14381 28543
rect 14148 28512 14381 28540
rect 14148 28500 14154 28512
rect 14369 28509 14381 28512
rect 14415 28509 14427 28543
rect 14369 28503 14427 28509
rect 8113 28475 8171 28481
rect 8113 28441 8125 28475
rect 8159 28472 8171 28475
rect 8202 28472 8208 28484
rect 8159 28444 8208 28472
rect 8159 28441 8171 28444
rect 8113 28435 8171 28441
rect 8202 28432 8208 28444
rect 8260 28432 8266 28484
rect 14568 28481 14596 28648
rect 15289 28645 15301 28679
rect 15335 28676 15347 28679
rect 15841 28679 15899 28685
rect 15841 28676 15853 28679
rect 15335 28648 15853 28676
rect 15335 28645 15347 28648
rect 15289 28639 15347 28645
rect 15841 28645 15853 28648
rect 15887 28645 15899 28679
rect 15841 28639 15899 28645
rect 15933 28679 15991 28685
rect 15933 28645 15945 28679
rect 15979 28645 15991 28679
rect 15933 28639 15991 28645
rect 14826 28568 14832 28620
rect 14884 28608 14890 28620
rect 15746 28608 15752 28620
rect 14884 28580 15752 28608
rect 14884 28568 14890 28580
rect 15746 28568 15752 28580
rect 15804 28568 15810 28620
rect 15856 28608 15884 28639
rect 17862 28608 17868 28620
rect 15856 28580 17868 28608
rect 17862 28568 17868 28580
rect 17920 28568 17926 28620
rect 15286 28500 15292 28552
rect 15344 28540 15350 28552
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 15344 28512 15577 28540
rect 15344 28500 15350 28512
rect 15565 28509 15577 28512
rect 15611 28509 15623 28543
rect 15565 28503 15623 28509
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28540 16359 28543
rect 23658 28540 23664 28552
rect 16347 28512 23664 28540
rect 16347 28509 16359 28512
rect 16301 28503 16359 28509
rect 23658 28500 23664 28512
rect 23716 28500 23722 28552
rect 14553 28475 14611 28481
rect 14553 28441 14565 28475
rect 14599 28472 14611 28475
rect 37918 28472 37924 28484
rect 14599 28444 37924 28472
rect 14599 28441 14611 28444
rect 14553 28435 14611 28441
rect 37918 28432 37924 28444
rect 37976 28432 37982 28484
rect 4249 28407 4307 28413
rect 4249 28373 4261 28407
rect 4295 28404 4307 28407
rect 4614 28404 4620 28416
rect 4295 28376 4620 28404
rect 4295 28373 4307 28376
rect 4249 28367 4307 28373
rect 4614 28364 4620 28376
rect 4672 28364 4678 28416
rect 8294 28404 8300 28416
rect 8255 28376 8300 28404
rect 8294 28364 8300 28376
rect 8352 28364 8358 28416
rect 9858 28404 9864 28416
rect 9819 28376 9864 28404
rect 9858 28364 9864 28376
rect 9916 28364 9922 28416
rect 11425 28407 11483 28413
rect 11425 28373 11437 28407
rect 11471 28404 11483 28407
rect 12710 28404 12716 28416
rect 11471 28376 12716 28404
rect 11471 28373 11483 28376
rect 11425 28367 11483 28373
rect 12710 28364 12716 28376
rect 12768 28364 12774 28416
rect 13541 28407 13599 28413
rect 13541 28373 13553 28407
rect 13587 28404 13599 28407
rect 15013 28407 15071 28413
rect 15013 28404 15025 28407
rect 13587 28376 15025 28404
rect 13587 28373 13599 28376
rect 13541 28367 13599 28373
rect 15013 28373 15025 28376
rect 15059 28404 15071 28407
rect 15289 28407 15347 28413
rect 15289 28404 15301 28407
rect 15059 28376 15301 28404
rect 15059 28373 15071 28376
rect 15013 28367 15071 28373
rect 15289 28373 15301 28376
rect 15335 28373 15347 28407
rect 15289 28367 15347 28373
rect 25222 28364 25228 28416
rect 25280 28404 25286 28416
rect 26234 28404 26240 28416
rect 25280 28376 26240 28404
rect 25280 28364 25286 28376
rect 26234 28364 26240 28376
rect 26292 28364 26298 28416
rect 1104 28314 29256 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 29256 28314
rect 1104 28240 29256 28262
rect 9582 28160 9588 28212
rect 9640 28200 9646 28212
rect 9769 28203 9827 28209
rect 9769 28200 9781 28203
rect 9640 28172 9781 28200
rect 9640 28160 9646 28172
rect 9769 28169 9781 28172
rect 9815 28169 9827 28203
rect 9769 28163 9827 28169
rect 2590 28064 2596 28076
rect 2551 28036 2596 28064
rect 2590 28024 2596 28036
rect 2648 28024 2654 28076
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28064 2927 28067
rect 3510 28064 3516 28076
rect 2915 28036 3516 28064
rect 2915 28033 2927 28036
rect 2869 28027 2927 28033
rect 3510 28024 3516 28036
rect 3568 28024 3574 28076
rect 8113 27999 8171 28005
rect 8113 27965 8125 27999
rect 8159 27965 8171 27999
rect 9784 27996 9812 28163
rect 11054 28160 11060 28212
rect 11112 28200 11118 28212
rect 16390 28200 16396 28212
rect 11112 28172 16396 28200
rect 11112 28160 11118 28172
rect 16390 28160 16396 28172
rect 16448 28160 16454 28212
rect 17862 28160 17868 28212
rect 17920 28200 17926 28212
rect 18417 28203 18475 28209
rect 18417 28200 18429 28203
rect 17920 28172 18429 28200
rect 17920 28160 17926 28172
rect 18417 28169 18429 28172
rect 18463 28169 18475 28203
rect 20254 28200 20260 28212
rect 20215 28172 20260 28200
rect 18417 28163 18475 28169
rect 20254 28160 20260 28172
rect 20312 28160 20318 28212
rect 21174 28200 21180 28212
rect 21135 28172 21180 28200
rect 21174 28160 21180 28172
rect 21232 28160 21238 28212
rect 24489 28203 24547 28209
rect 24489 28169 24501 28203
rect 24535 28200 24547 28203
rect 24946 28200 24952 28212
rect 24535 28172 24952 28200
rect 24535 28169 24547 28172
rect 24489 28163 24547 28169
rect 24946 28160 24952 28172
rect 25004 28200 25010 28212
rect 25590 28200 25596 28212
rect 25004 28172 25596 28200
rect 25004 28160 25010 28172
rect 25590 28160 25596 28172
rect 25648 28160 25654 28212
rect 9858 28092 9864 28144
rect 9916 28132 9922 28144
rect 10045 28135 10103 28141
rect 10045 28132 10057 28135
rect 9916 28104 10057 28132
rect 9916 28092 9922 28104
rect 10045 28101 10057 28104
rect 10091 28132 10103 28135
rect 13814 28132 13820 28144
rect 10091 28104 13820 28132
rect 10091 28101 10103 28104
rect 10045 28095 10103 28101
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 14918 28132 14924 28144
rect 14476 28104 14924 28132
rect 14476 28076 14504 28104
rect 14918 28092 14924 28104
rect 14976 28092 14982 28144
rect 15105 28135 15163 28141
rect 15105 28101 15117 28135
rect 15151 28132 15163 28135
rect 48314 28132 48320 28144
rect 15151 28104 48320 28132
rect 15151 28101 15163 28104
rect 15105 28095 15163 28101
rect 10686 28064 10692 28076
rect 10647 28036 10692 28064
rect 10686 28024 10692 28036
rect 10744 28024 10750 28076
rect 13906 28024 13912 28076
rect 13964 28064 13970 28076
rect 14458 28064 14464 28076
rect 13964 28036 14464 28064
rect 13964 28024 13970 28036
rect 14458 28024 14464 28036
rect 14516 28024 14522 28076
rect 9953 27999 10011 28005
rect 9953 27996 9965 27999
rect 9784 27968 9965 27996
rect 8113 27959 8171 27965
rect 9953 27965 9965 27968
rect 9999 27965 10011 27999
rect 9953 27959 10011 27965
rect 2958 27820 2964 27872
rect 3016 27860 3022 27872
rect 3973 27863 4031 27869
rect 3973 27860 3985 27863
rect 3016 27832 3985 27860
rect 3016 27820 3022 27832
rect 3973 27829 3985 27832
rect 4019 27829 4031 27863
rect 3973 27823 4031 27829
rect 4433 27863 4491 27869
rect 4433 27829 4445 27863
rect 4479 27860 4491 27863
rect 4890 27860 4896 27872
rect 4479 27832 4896 27860
rect 4479 27829 4491 27832
rect 4433 27823 4491 27829
rect 4890 27820 4896 27832
rect 4948 27820 4954 27872
rect 8021 27863 8079 27869
rect 8021 27829 8033 27863
rect 8067 27860 8079 27863
rect 8128 27860 8156 27959
rect 10134 27956 10140 28008
rect 10192 27996 10198 28008
rect 10229 27999 10287 28005
rect 10229 27996 10241 27999
rect 10192 27968 10241 27996
rect 10192 27956 10198 27968
rect 10229 27965 10241 27968
rect 10275 27965 10287 27999
rect 10229 27959 10287 27965
rect 14274 27956 14280 28008
rect 14332 27996 14338 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 14332 27968 14933 27996
rect 14332 27956 14338 27968
rect 14921 27965 14933 27968
rect 14967 27965 14979 27999
rect 14921 27959 14979 27965
rect 12618 27888 12624 27940
rect 12676 27928 12682 27940
rect 13998 27928 14004 27940
rect 12676 27900 14004 27928
rect 12676 27888 12682 27900
rect 13998 27888 14004 27900
rect 14056 27928 14062 27940
rect 14185 27931 14243 27937
rect 14185 27928 14197 27931
rect 14056 27900 14197 27928
rect 14056 27888 14062 27900
rect 14185 27897 14197 27900
rect 14231 27897 14243 27931
rect 14458 27928 14464 27940
rect 14419 27900 14464 27928
rect 14185 27891 14243 27897
rect 14458 27888 14464 27900
rect 14516 27888 14522 27940
rect 14553 27931 14611 27937
rect 14553 27897 14565 27931
rect 14599 27928 14611 27931
rect 15120 27928 15148 28095
rect 48314 28092 48320 28104
rect 48372 28092 48378 28144
rect 15194 28024 15200 28076
rect 15252 28064 15258 28076
rect 15749 28067 15807 28073
rect 15749 28064 15761 28067
rect 15252 28036 15761 28064
rect 15252 28024 15258 28036
rect 15749 28033 15761 28036
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 17862 28024 17868 28076
rect 17920 28064 17926 28076
rect 19889 28067 19947 28073
rect 17920 28036 19472 28064
rect 17920 28024 17926 28036
rect 19153 27999 19211 28005
rect 19153 27965 19165 27999
rect 19199 27965 19211 27999
rect 19334 27996 19340 28008
rect 19295 27968 19340 27996
rect 19153 27959 19211 27965
rect 14599 27900 15148 27928
rect 14599 27897 14611 27900
rect 14553 27891 14611 27897
rect 15746 27888 15752 27940
rect 15804 27928 15810 27940
rect 15933 27931 15991 27937
rect 15933 27928 15945 27931
rect 15804 27900 15945 27928
rect 15804 27888 15810 27900
rect 15933 27897 15945 27900
rect 15979 27897 15991 27931
rect 16114 27928 16120 27940
rect 16075 27900 16120 27928
rect 15933 27891 15991 27897
rect 16114 27888 16120 27900
rect 16172 27888 16178 27940
rect 16485 27931 16543 27937
rect 16485 27897 16497 27931
rect 16531 27928 16543 27931
rect 16758 27928 16764 27940
rect 16531 27900 16764 27928
rect 16531 27897 16543 27900
rect 16485 27891 16543 27897
rect 16758 27888 16764 27900
rect 16816 27888 16822 27940
rect 18138 27888 18144 27940
rect 18196 27928 18202 27940
rect 18601 27931 18659 27937
rect 18601 27928 18613 27931
rect 18196 27900 18613 27928
rect 18196 27888 18202 27900
rect 18601 27897 18613 27900
rect 18647 27897 18659 27931
rect 19168 27928 19196 27959
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 19444 28005 19472 28036
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20254 28064 20260 28076
rect 19935 28036 20260 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20901 28067 20959 28073
rect 20901 28033 20913 28067
rect 20947 28064 20959 28067
rect 24762 28064 24768 28076
rect 20947 28036 21680 28064
rect 24723 28036 24768 28064
rect 20947 28033 20959 28036
rect 20901 28027 20959 28033
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27965 19487 27999
rect 19978 27996 19984 28008
rect 19939 27968 19984 27996
rect 19429 27959 19487 27965
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 20806 27956 20812 28008
rect 20864 27996 20870 28008
rect 20993 27999 21051 28005
rect 20993 27996 21005 27999
rect 20864 27968 21005 27996
rect 20864 27956 20870 27968
rect 20993 27965 21005 27968
rect 21039 27965 21051 27999
rect 20993 27959 21051 27965
rect 19886 27928 19892 27940
rect 19168 27900 19892 27928
rect 18601 27891 18659 27897
rect 19886 27888 19892 27900
rect 19944 27928 19950 27940
rect 21652 27937 21680 28036
rect 24762 28024 24768 28036
rect 24820 28024 24826 28076
rect 25317 28067 25375 28073
rect 25317 28033 25329 28067
rect 25363 28064 25375 28067
rect 27522 28064 27528 28076
rect 25363 28036 27528 28064
rect 25363 28033 25375 28036
rect 25317 28027 25375 28033
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 25038 27956 25044 28008
rect 25096 27996 25102 28008
rect 25179 27999 25237 28005
rect 25179 27996 25191 27999
rect 25096 27968 25191 27996
rect 25096 27956 25102 27968
rect 25179 27965 25191 27968
rect 25225 27965 25237 27999
rect 25590 27996 25596 28008
rect 25551 27968 25596 27996
rect 25179 27959 25237 27965
rect 25590 27956 25596 27968
rect 25648 27956 25654 28008
rect 25777 27999 25835 28005
rect 25777 27965 25789 27999
rect 25823 27996 25835 27999
rect 27430 27996 27436 28008
rect 25823 27968 27436 27996
rect 25823 27965 25835 27968
rect 25777 27959 25835 27965
rect 27430 27956 27436 27968
rect 27488 27956 27494 28008
rect 20349 27931 20407 27937
rect 20349 27928 20361 27931
rect 19944 27900 20361 27928
rect 19944 27888 19950 27900
rect 20349 27897 20361 27900
rect 20395 27897 20407 27931
rect 20349 27891 20407 27897
rect 21637 27931 21695 27937
rect 21637 27897 21649 27931
rect 21683 27928 21695 27931
rect 67910 27928 67916 27940
rect 21683 27900 67916 27928
rect 21683 27897 21695 27900
rect 21637 27891 21695 27897
rect 67910 27888 67916 27900
rect 67968 27888 67974 27940
rect 8202 27860 8208 27872
rect 8067 27832 8208 27860
rect 8067 27829 8079 27832
rect 8021 27823 8079 27829
rect 8202 27820 8208 27832
rect 8260 27820 8266 27872
rect 8297 27863 8355 27869
rect 8297 27829 8309 27863
rect 8343 27860 8355 27863
rect 9674 27860 9680 27872
rect 8343 27832 9680 27860
rect 8343 27829 8355 27832
rect 8297 27823 8355 27829
rect 9674 27820 9680 27832
rect 9732 27820 9738 27872
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 14366 27860 14372 27872
rect 13872 27832 14372 27860
rect 13872 27820 13878 27832
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 14918 27820 14924 27872
rect 14976 27860 14982 27872
rect 16025 27863 16083 27869
rect 16025 27860 16037 27863
rect 14976 27832 16037 27860
rect 14976 27820 14982 27832
rect 16025 27829 16037 27832
rect 16071 27829 16083 27863
rect 16025 27823 16083 27829
rect 1104 27770 29256 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 29256 27770
rect 1104 27696 29256 27718
rect 13814 27656 13820 27668
rect 13775 27628 13820 27656
rect 13814 27616 13820 27628
rect 13872 27616 13878 27668
rect 13924 27628 14136 27656
rect 8757 27591 8815 27597
rect 8757 27557 8769 27591
rect 8803 27588 8815 27591
rect 13924 27588 13952 27628
rect 8803 27560 13952 27588
rect 14001 27591 14059 27597
rect 8803 27557 8815 27560
rect 8757 27551 8815 27557
rect 14001 27557 14013 27591
rect 14047 27557 14059 27591
rect 14108 27588 14136 27628
rect 14182 27616 14188 27668
rect 14240 27656 14246 27668
rect 16114 27656 16120 27668
rect 14240 27628 16120 27656
rect 14240 27616 14246 27628
rect 16114 27616 16120 27628
rect 16172 27616 16178 27668
rect 17862 27616 17868 27668
rect 17920 27656 17926 27668
rect 18233 27659 18291 27665
rect 18233 27656 18245 27659
rect 17920 27628 18245 27656
rect 17920 27616 17926 27628
rect 18233 27625 18245 27628
rect 18279 27656 18291 27659
rect 22741 27659 22799 27665
rect 18279 27628 19380 27656
rect 18279 27625 18291 27628
rect 18233 27619 18291 27625
rect 14108 27560 19104 27588
rect 14001 27551 14059 27557
rect 6917 27523 6975 27529
rect 6917 27489 6929 27523
rect 6963 27520 6975 27523
rect 7282 27520 7288 27532
rect 6963 27492 7288 27520
rect 6963 27489 6975 27492
rect 6917 27483 6975 27489
rect 7282 27480 7288 27492
rect 7340 27520 7346 27532
rect 8021 27523 8079 27529
rect 8021 27520 8033 27523
rect 7340 27492 8033 27520
rect 7340 27480 7346 27492
rect 8021 27489 8033 27492
rect 8067 27489 8079 27523
rect 8021 27483 8079 27489
rect 8297 27523 8355 27529
rect 8297 27489 8309 27523
rect 8343 27489 8355 27523
rect 8297 27483 8355 27489
rect 9677 27523 9735 27529
rect 9677 27489 9689 27523
rect 9723 27520 9735 27523
rect 9858 27520 9864 27532
rect 9723 27492 9864 27520
rect 9723 27489 9735 27492
rect 9677 27483 9735 27489
rect 8312 27452 8340 27483
rect 9858 27480 9864 27492
rect 9916 27480 9922 27532
rect 9953 27523 10011 27529
rect 9953 27489 9965 27523
rect 9999 27520 10011 27523
rect 9999 27492 10180 27520
rect 9999 27489 10011 27492
rect 9953 27483 10011 27489
rect 8386 27452 8392 27464
rect 8299 27424 8392 27452
rect 8386 27412 8392 27424
rect 8444 27452 8450 27464
rect 10152 27452 10180 27492
rect 10226 27480 10232 27532
rect 10284 27520 10290 27532
rect 11241 27523 11299 27529
rect 11241 27520 11253 27523
rect 10284 27492 11253 27520
rect 10284 27480 10290 27492
rect 11241 27489 11253 27492
rect 11287 27489 11299 27523
rect 12526 27520 12532 27532
rect 12487 27492 12532 27520
rect 11241 27483 11299 27489
rect 12526 27480 12532 27492
rect 12584 27480 12590 27532
rect 13630 27520 13636 27532
rect 13591 27492 13636 27520
rect 13630 27480 13636 27492
rect 13688 27480 13694 27532
rect 13906 27520 13912 27532
rect 13867 27492 13912 27520
rect 13906 27480 13912 27492
rect 13964 27480 13970 27532
rect 14016 27520 14044 27551
rect 14182 27520 14188 27532
rect 14016 27492 14188 27520
rect 14182 27480 14188 27492
rect 14240 27480 14246 27532
rect 14458 27480 14464 27532
rect 14516 27520 14522 27532
rect 15381 27523 15439 27529
rect 15381 27520 15393 27523
rect 14516 27492 15393 27520
rect 14516 27480 14522 27492
rect 15381 27489 15393 27492
rect 15427 27489 15439 27523
rect 15381 27483 15439 27489
rect 18969 27523 19027 27529
rect 18969 27489 18981 27523
rect 19015 27489 19027 27523
rect 18969 27483 19027 27489
rect 8444 27424 10180 27452
rect 8444 27412 8450 27424
rect 7929 27387 7987 27393
rect 7929 27353 7941 27387
rect 7975 27384 7987 27387
rect 8113 27387 8171 27393
rect 8113 27384 8125 27387
rect 7975 27356 8125 27384
rect 7975 27353 7987 27356
rect 7929 27347 7987 27353
rect 8113 27353 8125 27356
rect 8159 27384 8171 27387
rect 8202 27384 8208 27396
rect 8159 27356 8208 27384
rect 8159 27353 8171 27356
rect 8113 27347 8171 27353
rect 8202 27344 8208 27356
rect 8260 27344 8266 27396
rect 9766 27384 9772 27396
rect 9727 27356 9772 27384
rect 9766 27344 9772 27356
rect 9824 27344 9830 27396
rect 10152 27384 10180 27424
rect 10413 27455 10471 27461
rect 10413 27421 10425 27455
rect 10459 27452 10471 27455
rect 10686 27452 10692 27464
rect 10459 27424 10692 27452
rect 10459 27421 10471 27424
rect 10413 27415 10471 27421
rect 10686 27412 10692 27424
rect 10744 27412 10750 27464
rect 13648 27384 13676 27480
rect 14366 27452 14372 27464
rect 14327 27424 14372 27452
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 15286 27452 15292 27464
rect 15247 27424 15292 27452
rect 15286 27412 15292 27424
rect 15344 27412 15350 27464
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 15841 27455 15899 27461
rect 15841 27452 15853 27455
rect 15804 27424 15853 27452
rect 15804 27412 15810 27424
rect 15841 27421 15853 27424
rect 15887 27421 15899 27455
rect 15841 27415 15899 27421
rect 16298 27412 16304 27464
rect 16356 27452 16362 27464
rect 18417 27455 18475 27461
rect 18417 27452 18429 27455
rect 16356 27424 18429 27452
rect 16356 27412 16362 27424
rect 18417 27421 18429 27424
rect 18463 27421 18475 27455
rect 18417 27415 18475 27421
rect 10152 27356 13676 27384
rect 13722 27344 13728 27396
rect 13780 27384 13786 27396
rect 15654 27384 15660 27396
rect 13780 27356 15660 27384
rect 13780 27344 13786 27356
rect 15654 27344 15660 27356
rect 15712 27344 15718 27396
rect 7101 27319 7159 27325
rect 7101 27285 7113 27319
rect 7147 27316 7159 27319
rect 9582 27316 9588 27328
rect 7147 27288 9588 27316
rect 7147 27285 7159 27288
rect 7101 27279 7159 27285
rect 9582 27276 9588 27288
rect 9640 27276 9646 27328
rect 11425 27319 11483 27325
rect 11425 27285 11437 27319
rect 11471 27316 11483 27319
rect 12618 27316 12624 27328
rect 11471 27288 12624 27316
rect 11471 27285 11483 27288
rect 11425 27279 11483 27285
rect 12618 27276 12624 27288
rect 12676 27276 12682 27328
rect 12713 27319 12771 27325
rect 12713 27285 12725 27319
rect 12759 27316 12771 27319
rect 13906 27316 13912 27328
rect 12759 27288 13912 27316
rect 12759 27285 12771 27288
rect 12713 27279 12771 27285
rect 13906 27276 13912 27288
rect 13964 27276 13970 27328
rect 18984 27316 19012 27483
rect 19076 27384 19104 27560
rect 19153 27523 19211 27529
rect 19153 27489 19165 27523
rect 19199 27489 19211 27523
rect 19153 27483 19211 27489
rect 19245 27523 19303 27529
rect 19245 27489 19257 27523
rect 19291 27520 19303 27523
rect 19352 27520 19380 27628
rect 22741 27625 22753 27659
rect 22787 27625 22799 27659
rect 22741 27619 22799 27625
rect 22756 27588 22784 27619
rect 25038 27588 25044 27600
rect 22756 27560 25044 27588
rect 25038 27548 25044 27560
rect 25096 27548 25102 27600
rect 25685 27591 25743 27597
rect 25685 27588 25697 27591
rect 25516 27560 25697 27588
rect 19889 27523 19947 27529
rect 19291 27492 19380 27520
rect 19628 27492 19840 27520
rect 19291 27489 19303 27492
rect 19245 27483 19303 27489
rect 19168 27452 19196 27483
rect 19334 27452 19340 27464
rect 19168 27424 19340 27452
rect 19334 27412 19340 27424
rect 19392 27412 19398 27464
rect 19628 27384 19656 27492
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19812 27452 19840 27492
rect 19889 27489 19901 27523
rect 19935 27520 19947 27523
rect 20806 27520 20812 27532
rect 19935 27492 20812 27520
rect 19935 27489 19947 27492
rect 19889 27483 19947 27489
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 22563 27523 22621 27529
rect 22563 27489 22575 27523
rect 22609 27489 22621 27523
rect 22563 27483 22621 27489
rect 22572 27452 22600 27483
rect 23382 27480 23388 27532
rect 23440 27520 23446 27532
rect 24213 27523 24271 27529
rect 24213 27520 24225 27523
rect 23440 27492 24225 27520
rect 23440 27480 23446 27492
rect 24213 27489 24225 27492
rect 24259 27520 24271 27523
rect 24946 27520 24952 27532
rect 24259 27492 24952 27520
rect 24259 27489 24271 27492
rect 24213 27483 24271 27489
rect 24946 27480 24952 27492
rect 25004 27480 25010 27532
rect 25056 27520 25084 27548
rect 25314 27520 25320 27532
rect 25056 27492 25320 27520
rect 25314 27480 25320 27492
rect 25372 27480 25378 27532
rect 25516 27529 25544 27560
rect 25685 27557 25697 27560
rect 25731 27588 25743 27591
rect 35434 27588 35440 27600
rect 25731 27560 35440 27588
rect 25731 27557 25743 27560
rect 25685 27551 25743 27557
rect 35434 27548 35440 27560
rect 35492 27548 35498 27600
rect 25501 27523 25559 27529
rect 25501 27489 25513 27523
rect 25547 27489 25559 27523
rect 25501 27483 25559 27489
rect 26694 27480 26700 27532
rect 26752 27520 26758 27532
rect 27249 27523 27307 27529
rect 27249 27520 27261 27523
rect 26752 27492 27261 27520
rect 26752 27480 26758 27492
rect 27249 27489 27261 27492
rect 27295 27489 27307 27523
rect 27430 27520 27436 27532
rect 27391 27492 27436 27520
rect 27249 27483 27307 27489
rect 27430 27480 27436 27492
rect 27488 27480 27494 27532
rect 19812 27424 22600 27452
rect 19705 27415 19763 27421
rect 19076 27356 19656 27384
rect 19720 27384 19748 27415
rect 23474 27412 23480 27464
rect 23532 27452 23538 27464
rect 24305 27455 24363 27461
rect 24305 27452 24317 27455
rect 23532 27424 24317 27452
rect 23532 27412 23538 27424
rect 24305 27421 24317 27424
rect 24351 27421 24363 27455
rect 24305 27415 24363 27421
rect 25041 27455 25099 27461
rect 25041 27421 25053 27455
rect 25087 27452 25099 27455
rect 25866 27452 25872 27464
rect 25087 27424 25872 27452
rect 25087 27421 25099 27424
rect 25041 27415 25099 27421
rect 25866 27412 25872 27424
rect 25924 27412 25930 27464
rect 26234 27412 26240 27464
rect 26292 27452 26298 27464
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 26292 27424 26525 27452
rect 26292 27412 26298 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 20073 27387 20131 27393
rect 20073 27384 20085 27387
rect 19720 27356 20085 27384
rect 20073 27353 20085 27356
rect 20119 27384 20131 27387
rect 50154 27384 50160 27396
rect 20119 27356 50160 27384
rect 20119 27353 20131 27356
rect 20073 27347 20131 27353
rect 50154 27344 50160 27356
rect 50212 27344 50218 27396
rect 20162 27316 20168 27328
rect 18984 27288 20168 27316
rect 20162 27276 20168 27288
rect 20220 27276 20226 27328
rect 25866 27316 25872 27328
rect 25827 27288 25872 27316
rect 25866 27276 25872 27288
rect 25924 27276 25930 27328
rect 26234 27316 26240 27328
rect 26195 27288 26240 27316
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 26786 27276 26792 27328
rect 26844 27316 26850 27328
rect 27709 27319 27767 27325
rect 27709 27316 27721 27319
rect 26844 27288 27721 27316
rect 26844 27276 26850 27288
rect 27709 27285 27721 27288
rect 27755 27285 27767 27319
rect 27709 27279 27767 27285
rect 1104 27226 29256 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 29256 27226
rect 1104 27152 29256 27174
rect 4709 27115 4767 27121
rect 4709 27081 4721 27115
rect 4755 27112 4767 27115
rect 4982 27112 4988 27124
rect 4755 27084 4988 27112
rect 4755 27081 4767 27084
rect 4709 27075 4767 27081
rect 3973 26911 4031 26917
rect 3973 26877 3985 26911
rect 4019 26908 4031 26911
rect 4724 26908 4752 27075
rect 4982 27072 4988 27084
rect 5040 27072 5046 27124
rect 7282 27112 7288 27124
rect 7243 27084 7288 27112
rect 7282 27072 7288 27084
rect 7340 27072 7346 27124
rect 9858 27072 9864 27124
rect 9916 27112 9922 27124
rect 9916 27084 10640 27112
rect 9916 27072 9922 27084
rect 8294 27044 8300 27056
rect 8255 27016 8300 27044
rect 8294 27004 8300 27016
rect 8352 27044 8358 27056
rect 9953 27047 10011 27053
rect 9953 27044 9965 27047
rect 8352 27016 9965 27044
rect 8352 27004 8358 27016
rect 9953 27013 9965 27016
rect 9999 27013 10011 27047
rect 9953 27007 10011 27013
rect 8941 26979 8999 26985
rect 8941 26945 8953 26979
rect 8987 26976 8999 26979
rect 10612 26976 10640 27084
rect 10686 27072 10692 27124
rect 10744 27112 10750 27124
rect 15930 27112 15936 27124
rect 10744 27084 15936 27112
rect 10744 27072 10750 27084
rect 15930 27072 15936 27084
rect 15988 27072 15994 27124
rect 23845 27115 23903 27121
rect 23845 27081 23857 27115
rect 23891 27112 23903 27115
rect 23934 27112 23940 27124
rect 23891 27084 23940 27112
rect 23891 27081 23903 27084
rect 23845 27075 23903 27081
rect 23934 27072 23940 27084
rect 23992 27112 23998 27124
rect 24578 27112 24584 27124
rect 23992 27084 24584 27112
rect 23992 27072 23998 27084
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 25866 27072 25872 27124
rect 25924 27112 25930 27124
rect 41874 27112 41880 27124
rect 25924 27084 41880 27112
rect 25924 27072 25930 27084
rect 41874 27072 41880 27084
rect 41932 27072 41938 27124
rect 14093 27047 14151 27053
rect 14093 27013 14105 27047
rect 14139 27044 14151 27047
rect 18598 27044 18604 27056
rect 14139 27016 18604 27044
rect 14139 27013 14151 27016
rect 14093 27007 14151 27013
rect 18598 27004 18604 27016
rect 18656 27004 18662 27056
rect 26142 27004 26148 27056
rect 26200 27044 26206 27056
rect 26329 27047 26387 27053
rect 26329 27044 26341 27047
rect 26200 27016 26341 27044
rect 26200 27004 26206 27016
rect 26329 27013 26341 27016
rect 26375 27044 26387 27047
rect 26375 27016 26556 27044
rect 26375 27013 26387 27016
rect 26329 27007 26387 27013
rect 12526 26976 12532 26988
rect 8987 26948 10548 26976
rect 10612 26948 12532 26976
rect 8987 26945 8999 26948
rect 8941 26939 8999 26945
rect 4019 26880 4752 26908
rect 7101 26911 7159 26917
rect 4019 26877 4031 26880
rect 3973 26871 4031 26877
rect 7101 26877 7113 26911
rect 7147 26908 7159 26911
rect 7193 26911 7251 26917
rect 7193 26908 7205 26911
rect 7147 26880 7205 26908
rect 7147 26877 7159 26880
rect 7101 26871 7159 26877
rect 7193 26877 7205 26880
rect 7239 26908 7251 26911
rect 8205 26911 8263 26917
rect 8205 26908 8217 26911
rect 7239 26880 8217 26908
rect 7239 26877 7251 26880
rect 7193 26871 7251 26877
rect 3789 26843 3847 26849
rect 3789 26809 3801 26843
rect 3835 26809 3847 26843
rect 3789 26803 3847 26809
rect 3418 26732 3424 26784
rect 3476 26772 3482 26784
rect 3694 26772 3700 26784
rect 3476 26744 3700 26772
rect 3476 26732 3482 26744
rect 3694 26732 3700 26744
rect 3752 26732 3758 26784
rect 3804 26772 3832 26803
rect 4246 26800 4252 26852
rect 4304 26840 4310 26852
rect 4341 26843 4399 26849
rect 4341 26840 4353 26843
rect 4304 26812 4353 26840
rect 4304 26800 4310 26812
rect 4341 26809 4353 26812
rect 4387 26809 4399 26843
rect 4341 26803 4399 26809
rect 7944 26784 7972 26880
rect 8205 26877 8217 26880
rect 8251 26877 8263 26911
rect 8481 26911 8539 26917
rect 8481 26908 8493 26911
rect 8205 26871 8263 26877
rect 8312 26880 8493 26908
rect 8312 26784 8340 26880
rect 8481 26877 8493 26880
rect 8527 26877 8539 26911
rect 9858 26908 9864 26920
rect 9819 26880 9864 26908
rect 8481 26871 8539 26877
rect 9858 26868 9864 26880
rect 9916 26868 9922 26920
rect 10134 26908 10140 26920
rect 10095 26880 10140 26908
rect 10134 26868 10140 26880
rect 10192 26868 10198 26920
rect 10520 26908 10548 26948
rect 12526 26936 12532 26948
rect 12584 26976 12590 26988
rect 26528 26985 26556 27016
rect 15289 26979 15347 26985
rect 15289 26976 15301 26979
rect 12584 26948 15301 26976
rect 12584 26936 12590 26948
rect 13722 26908 13728 26920
rect 10520 26880 13728 26908
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 13998 26868 14004 26920
rect 14056 26908 14062 26920
rect 14752 26917 14780 26948
rect 15289 26945 15301 26948
rect 15335 26945 15347 26979
rect 15289 26939 15347 26945
rect 26513 26979 26571 26985
rect 26513 26945 26525 26979
rect 26559 26945 26571 26979
rect 26786 26976 26792 26988
rect 26747 26948 26792 26976
rect 26513 26939 26571 26945
rect 26786 26936 26792 26948
rect 26844 26936 26850 26988
rect 14737 26911 14795 26917
rect 14056 26880 14688 26908
rect 14056 26868 14062 26880
rect 10597 26843 10655 26849
rect 10597 26809 10609 26843
rect 10643 26840 10655 26843
rect 10686 26840 10692 26852
rect 10643 26812 10692 26840
rect 10643 26809 10655 26812
rect 10597 26803 10655 26809
rect 10686 26800 10692 26812
rect 10744 26800 10750 26852
rect 14093 26843 14151 26849
rect 14093 26809 14105 26843
rect 14139 26840 14151 26843
rect 14185 26843 14243 26849
rect 14185 26840 14197 26843
rect 14139 26812 14197 26840
rect 14139 26809 14151 26812
rect 14093 26803 14151 26809
rect 14185 26809 14197 26812
rect 14231 26809 14243 26843
rect 14660 26840 14688 26880
rect 14737 26877 14749 26911
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 14826 26868 14832 26920
rect 14884 26908 14890 26920
rect 15013 26911 15071 26917
rect 14884 26880 14929 26908
rect 14884 26868 14890 26880
rect 15013 26877 15025 26911
rect 15059 26908 15071 26911
rect 15102 26908 15108 26920
rect 15059 26880 15108 26908
rect 15059 26877 15071 26880
rect 15013 26871 15071 26877
rect 15028 26840 15056 26871
rect 15102 26868 15108 26880
rect 15160 26868 15166 26920
rect 15657 26911 15715 26917
rect 15657 26877 15669 26911
rect 15703 26908 15715 26911
rect 15746 26908 15752 26920
rect 15703 26880 15752 26908
rect 15703 26877 15715 26880
rect 15657 26871 15715 26877
rect 15746 26868 15752 26880
rect 15804 26868 15810 26920
rect 23658 26908 23664 26920
rect 23619 26880 23664 26908
rect 23658 26868 23664 26880
rect 23716 26908 23722 26920
rect 24765 26911 24823 26917
rect 24765 26908 24777 26911
rect 23716 26880 24777 26908
rect 23716 26868 23722 26880
rect 24765 26877 24777 26880
rect 24811 26877 24823 26911
rect 24765 26871 24823 26877
rect 14660 26812 15056 26840
rect 14185 26803 14243 26809
rect 4522 26772 4528 26784
rect 3804 26744 4528 26772
rect 4522 26732 4528 26744
rect 4580 26732 4586 26784
rect 7926 26772 7932 26784
rect 7887 26744 7932 26772
rect 7926 26732 7932 26744
rect 7984 26732 7990 26784
rect 8018 26732 8024 26784
rect 8076 26772 8082 26784
rect 8294 26772 8300 26784
rect 8076 26744 8300 26772
rect 8076 26732 8082 26744
rect 8294 26732 8300 26744
rect 8352 26732 8358 26784
rect 9766 26732 9772 26784
rect 9824 26772 9830 26784
rect 14826 26772 14832 26784
rect 9824 26744 14832 26772
rect 9824 26732 9830 26744
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 24854 26732 24860 26784
rect 24912 26772 24918 26784
rect 24949 26775 25007 26781
rect 24949 26772 24961 26775
rect 24912 26744 24961 26772
rect 24912 26732 24918 26744
rect 24949 26741 24961 26744
rect 24995 26741 25007 26775
rect 28074 26772 28080 26784
rect 28035 26744 28080 26772
rect 24949 26735 25007 26741
rect 28074 26732 28080 26744
rect 28132 26732 28138 26784
rect 1104 26682 29256 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 29256 26682
rect 1104 26608 29256 26630
rect 5810 26528 5816 26580
rect 5868 26568 5874 26580
rect 6546 26568 6552 26580
rect 5868 26540 6552 26568
rect 5868 26528 5874 26540
rect 6546 26528 6552 26540
rect 6604 26528 6610 26580
rect 8386 26568 8392 26580
rect 8347 26540 8392 26568
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 9769 26571 9827 26577
rect 9769 26537 9781 26571
rect 9815 26568 9827 26571
rect 10134 26568 10140 26580
rect 9815 26540 10140 26568
rect 9815 26537 9827 26540
rect 9769 26531 9827 26537
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 24213 26571 24271 26577
rect 24213 26568 24225 26571
rect 23768 26540 24225 26568
rect 4246 26500 4252 26512
rect 4207 26472 4252 26500
rect 4246 26460 4252 26472
rect 4304 26460 4310 26512
rect 4522 26460 4528 26512
rect 4580 26500 4586 26512
rect 5629 26503 5687 26509
rect 5629 26500 5641 26503
rect 4580 26472 5641 26500
rect 4580 26460 4586 26472
rect 5629 26469 5641 26472
rect 5675 26500 5687 26503
rect 6365 26503 6423 26509
rect 6365 26500 6377 26503
rect 5675 26472 6377 26500
rect 5675 26469 5687 26472
rect 5629 26463 5687 26469
rect 6365 26469 6377 26472
rect 6411 26500 6423 26503
rect 10594 26500 10600 26512
rect 6411 26472 10600 26500
rect 6411 26469 6423 26472
rect 6365 26463 6423 26469
rect 10594 26460 10600 26472
rect 10652 26460 10658 26512
rect 15746 26460 15752 26512
rect 15804 26500 15810 26512
rect 19334 26500 19340 26512
rect 15804 26472 19340 26500
rect 15804 26460 15810 26472
rect 4157 26435 4215 26441
rect 4157 26401 4169 26435
rect 4203 26401 4215 26435
rect 4157 26395 4215 26401
rect 4341 26435 4399 26441
rect 4341 26401 4353 26435
rect 4387 26432 4399 26435
rect 5166 26432 5172 26444
rect 4387 26404 5172 26432
rect 4387 26401 4399 26404
rect 4341 26395 4399 26401
rect 4172 26364 4200 26395
rect 5166 26392 5172 26404
rect 5224 26392 5230 26444
rect 5810 26432 5816 26444
rect 5771 26404 5816 26432
rect 5810 26392 5816 26404
rect 5868 26392 5874 26444
rect 8205 26435 8263 26441
rect 8205 26401 8217 26435
rect 8251 26432 8263 26435
rect 8294 26432 8300 26444
rect 8251 26404 8300 26432
rect 8251 26401 8263 26404
rect 8205 26395 8263 26401
rect 8294 26392 8300 26404
rect 8352 26432 8358 26444
rect 9677 26435 9735 26441
rect 9677 26432 9689 26435
rect 8352 26404 9689 26432
rect 8352 26392 8358 26404
rect 9677 26401 9689 26404
rect 9723 26432 9735 26435
rect 9953 26435 10011 26441
rect 9953 26432 9965 26435
rect 9723 26404 9965 26432
rect 9723 26401 9735 26404
rect 9677 26395 9735 26401
rect 9953 26401 9965 26404
rect 9999 26401 10011 26435
rect 10686 26432 10692 26444
rect 10647 26404 10692 26432
rect 9953 26395 10011 26401
rect 10686 26392 10692 26404
rect 10744 26392 10750 26444
rect 17328 26441 17356 26472
rect 19334 26460 19340 26472
rect 19392 26460 19398 26512
rect 22830 26460 22836 26512
rect 22888 26500 22894 26512
rect 23290 26500 23296 26512
rect 22888 26472 23296 26500
rect 22888 26460 22894 26472
rect 23290 26460 23296 26472
rect 23348 26500 23354 26512
rect 23768 26500 23796 26540
rect 24213 26537 24225 26540
rect 24259 26537 24271 26571
rect 24213 26531 24271 26537
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 28077 26571 28135 26577
rect 28077 26568 28089 26571
rect 27488 26540 28089 26568
rect 27488 26528 27494 26540
rect 28077 26537 28089 26540
rect 28123 26537 28135 26571
rect 28077 26531 28135 26537
rect 28166 26528 28172 26580
rect 28224 26568 28230 26580
rect 28224 26540 31708 26568
rect 28224 26528 28230 26540
rect 24121 26503 24179 26509
rect 24121 26500 24133 26503
rect 23348 26472 23796 26500
rect 23348 26460 23354 26472
rect 17313 26435 17371 26441
rect 17313 26401 17325 26435
rect 17359 26401 17371 26435
rect 17313 26395 17371 26401
rect 17402 26392 17408 26444
rect 17460 26432 17466 26444
rect 18601 26435 18659 26441
rect 18601 26432 18613 26435
rect 17460 26404 18613 26432
rect 17460 26392 17466 26404
rect 18601 26401 18613 26404
rect 18647 26401 18659 26435
rect 18601 26395 18659 26401
rect 22370 26392 22376 26444
rect 22428 26432 22434 26444
rect 22649 26435 22707 26441
rect 22649 26432 22661 26435
rect 22428 26404 22661 26432
rect 22428 26392 22434 26404
rect 22649 26401 22661 26404
rect 22695 26432 22707 26435
rect 23382 26432 23388 26444
rect 22695 26404 23388 26432
rect 22695 26401 22707 26404
rect 22649 26395 22707 26401
rect 23382 26392 23388 26404
rect 23440 26392 23446 26444
rect 23768 26441 23796 26472
rect 23952 26472 24133 26500
rect 23952 26441 23980 26472
rect 24121 26469 24133 26472
rect 24167 26500 24179 26503
rect 31680 26500 31708 26540
rect 63494 26528 63500 26580
rect 63552 26528 63558 26580
rect 57882 26500 57888 26512
rect 24167 26472 28488 26500
rect 31680 26472 57888 26500
rect 24167 26469 24179 26472
rect 24121 26463 24179 26469
rect 23753 26435 23811 26441
rect 23753 26401 23765 26435
rect 23799 26401 23811 26435
rect 23753 26395 23811 26401
rect 23937 26435 23995 26441
rect 23937 26401 23949 26435
rect 23983 26401 23995 26435
rect 24762 26432 24768 26444
rect 24723 26404 24768 26432
rect 23937 26395 23995 26401
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 27985 26435 28043 26441
rect 27985 26401 27997 26435
rect 28031 26432 28043 26435
rect 28074 26432 28080 26444
rect 28031 26404 28080 26432
rect 28031 26401 28043 26404
rect 27985 26395 28043 26401
rect 28074 26392 28080 26404
rect 28132 26432 28138 26444
rect 28132 26404 28396 26432
rect 28132 26392 28138 26404
rect 4614 26364 4620 26376
rect 4172 26336 4620 26364
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 4706 26324 4712 26376
rect 4764 26364 4770 26376
rect 4801 26367 4859 26373
rect 4801 26364 4813 26367
rect 4764 26336 4813 26364
rect 4764 26324 4770 26336
rect 4801 26333 4813 26336
rect 4847 26333 4859 26367
rect 4801 26327 4859 26333
rect 5350 26324 5356 26376
rect 5408 26364 5414 26376
rect 6089 26367 6147 26373
rect 6089 26364 6101 26367
rect 5408 26336 6101 26364
rect 5408 26324 5414 26336
rect 6089 26333 6101 26336
rect 6135 26333 6147 26367
rect 6089 26327 6147 26333
rect 17129 26367 17187 26373
rect 17129 26333 17141 26367
rect 17175 26364 17187 26367
rect 17221 26367 17279 26373
rect 17221 26364 17233 26367
rect 17175 26336 17233 26364
rect 17175 26333 17187 26336
rect 17129 26327 17187 26333
rect 17221 26333 17233 26336
rect 17267 26364 17279 26367
rect 17862 26364 17868 26376
rect 17267 26336 17868 26364
rect 17267 26333 17279 26336
rect 17221 26327 17279 26333
rect 17862 26324 17868 26336
rect 17920 26324 17926 26376
rect 18782 26373 18788 26376
rect 18748 26367 18788 26373
rect 18748 26333 18760 26367
rect 18748 26327 18788 26333
rect 18782 26324 18788 26327
rect 18840 26324 18846 26376
rect 18969 26367 19027 26373
rect 18969 26333 18981 26367
rect 19015 26364 19027 26367
rect 19426 26364 19432 26376
rect 19015 26336 19432 26364
rect 19015 26333 19027 26336
rect 18969 26327 19027 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 22738 26364 22744 26376
rect 22699 26336 22744 26364
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 24489 26367 24547 26373
rect 24489 26364 24501 26367
rect 23523 26336 24501 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 24489 26333 24501 26336
rect 24535 26364 24547 26367
rect 28166 26364 28172 26376
rect 24535 26336 28172 26364
rect 24535 26333 24547 26336
rect 24489 26327 24547 26333
rect 28166 26324 28172 26336
rect 28224 26324 28230 26376
rect 4632 26296 4660 26324
rect 4982 26296 4988 26308
rect 4632 26268 4988 26296
rect 4982 26256 4988 26268
rect 5040 26256 5046 26308
rect 10873 26299 10931 26305
rect 10873 26265 10885 26299
rect 10919 26296 10931 26299
rect 11606 26296 11612 26308
rect 10919 26268 11612 26296
rect 10919 26265 10931 26268
rect 10873 26259 10931 26265
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 28368 26305 28396 26404
rect 28460 26364 28488 26472
rect 57882 26460 57888 26472
rect 57940 26460 57946 26512
rect 63512 26364 63540 26528
rect 28460 26336 63540 26364
rect 18877 26299 18935 26305
rect 14384 26268 18828 26296
rect 5166 26228 5172 26240
rect 5127 26200 5172 26228
rect 5166 26188 5172 26200
rect 5224 26188 5230 26240
rect 8018 26228 8024 26240
rect 7979 26200 8024 26228
rect 8018 26188 8024 26200
rect 8076 26188 8082 26240
rect 8294 26188 8300 26240
rect 8352 26228 8358 26240
rect 14384 26228 14412 26268
rect 17494 26228 17500 26240
rect 8352 26200 14412 26228
rect 17455 26200 17500 26228
rect 8352 26188 8358 26200
rect 17494 26188 17500 26200
rect 17552 26188 17558 26240
rect 18800 26228 18828 26268
rect 18877 26265 18889 26299
rect 18923 26296 18935 26299
rect 24857 26299 24915 26305
rect 24857 26296 24869 26299
rect 18923 26268 24869 26296
rect 18923 26265 18935 26268
rect 18877 26259 18935 26265
rect 24857 26265 24869 26268
rect 24903 26265 24915 26299
rect 24857 26259 24915 26265
rect 28353 26299 28411 26305
rect 28353 26265 28365 26299
rect 28399 26296 28411 26299
rect 56686 26296 56692 26308
rect 28399 26268 56692 26296
rect 28399 26265 28411 26268
rect 28353 26259 28411 26265
rect 56686 26256 56692 26268
rect 56744 26256 56750 26308
rect 19061 26231 19119 26237
rect 19061 26228 19073 26231
rect 18800 26200 19073 26228
rect 19061 26197 19073 26200
rect 19107 26197 19119 26231
rect 19061 26191 19119 26197
rect 55122 26188 55128 26240
rect 55180 26228 55186 26240
rect 56594 26228 56600 26240
rect 55180 26200 56600 26228
rect 55180 26188 55186 26200
rect 56594 26188 56600 26200
rect 56652 26188 56658 26240
rect 1104 26138 29256 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 29256 26138
rect 1104 26064 29256 26086
rect 8297 26027 8355 26033
rect 8297 25993 8309 26027
rect 8343 26024 8355 26027
rect 9858 26024 9864 26036
rect 8343 25996 9864 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 9858 25984 9864 25996
rect 9916 25984 9922 26036
rect 15930 26024 15936 26036
rect 15891 25996 15936 26024
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 18414 26024 18420 26036
rect 18375 25996 18420 26024
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 18782 26024 18788 26036
rect 18743 25996 18788 26024
rect 18782 25984 18788 25996
rect 18840 25984 18846 26036
rect 3878 25916 3884 25968
rect 3936 25956 3942 25968
rect 9950 25956 9956 25968
rect 3936 25928 9956 25956
rect 3936 25916 3942 25928
rect 9950 25916 9956 25928
rect 10008 25916 10014 25968
rect 12710 25916 12716 25968
rect 12768 25956 12774 25968
rect 14921 25959 14979 25965
rect 14921 25956 14933 25959
rect 12768 25928 14933 25956
rect 12768 25916 12774 25928
rect 14921 25925 14933 25928
rect 14967 25925 14979 25959
rect 14921 25919 14979 25925
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25888 2927 25891
rect 4798 25888 4804 25900
rect 2915 25860 4804 25888
rect 2915 25857 2927 25860
rect 2869 25851 2927 25857
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 2593 25823 2651 25829
rect 2593 25789 2605 25823
rect 2639 25789 2651 25823
rect 8113 25823 8171 25829
rect 8113 25820 8125 25823
rect 2593 25783 2651 25789
rect 7944 25792 8125 25820
rect 2608 25684 2636 25783
rect 3528 25724 4476 25752
rect 3528 25684 3556 25724
rect 4448 25696 4476 25724
rect 7944 25696 7972 25792
rect 8113 25789 8125 25792
rect 8159 25789 8171 25823
rect 14936 25820 14964 25919
rect 18432 25888 18460 25984
rect 18509 25891 18567 25897
rect 18509 25888 18521 25891
rect 18432 25860 18521 25888
rect 18509 25857 18521 25860
rect 18555 25857 18567 25891
rect 18509 25851 18567 25857
rect 15105 25823 15163 25829
rect 15105 25820 15117 25823
rect 14936 25792 15117 25820
rect 8113 25783 8171 25789
rect 15105 25789 15117 25792
rect 15151 25789 15163 25823
rect 15105 25783 15163 25789
rect 15930 25780 15936 25832
rect 15988 25820 15994 25832
rect 16117 25823 16175 25829
rect 16117 25820 16129 25823
rect 15988 25792 16129 25820
rect 15988 25780 15994 25792
rect 16117 25789 16129 25792
rect 16163 25789 16175 25823
rect 18598 25820 18604 25832
rect 18559 25792 18604 25820
rect 16117 25783 16175 25789
rect 18598 25780 18604 25792
rect 18656 25820 18662 25832
rect 18966 25820 18972 25832
rect 18656 25792 18972 25820
rect 18656 25780 18662 25792
rect 18966 25780 18972 25792
rect 19024 25780 19030 25832
rect 2608 25656 3556 25684
rect 3786 25644 3792 25696
rect 3844 25684 3850 25696
rect 3973 25687 4031 25693
rect 3973 25684 3985 25687
rect 3844 25656 3985 25684
rect 3844 25644 3850 25656
rect 3973 25653 3985 25656
rect 4019 25653 4031 25687
rect 4430 25684 4436 25696
rect 4391 25656 4436 25684
rect 3973 25647 4031 25653
rect 4430 25644 4436 25656
rect 4488 25644 4494 25696
rect 7926 25684 7932 25696
rect 7887 25656 7932 25684
rect 7926 25644 7932 25656
rect 7984 25644 7990 25696
rect 15197 25687 15255 25693
rect 15197 25653 15209 25687
rect 15243 25684 15255 25687
rect 15838 25684 15844 25696
rect 15243 25656 15844 25684
rect 15243 25653 15255 25656
rect 15197 25647 15255 25653
rect 15838 25644 15844 25656
rect 15896 25644 15902 25696
rect 16206 25684 16212 25696
rect 16167 25656 16212 25684
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 1104 25594 29256 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 29256 25594
rect 1104 25520 29256 25542
rect 11606 25440 11612 25492
rect 11664 25480 11670 25492
rect 13081 25483 13139 25489
rect 13081 25480 13093 25483
rect 11664 25452 13093 25480
rect 11664 25440 11670 25452
rect 13081 25449 13093 25452
rect 13127 25480 13139 25483
rect 21637 25483 21695 25489
rect 21637 25480 21649 25483
rect 13127 25452 21649 25480
rect 13127 25449 13139 25452
rect 13081 25443 13139 25449
rect 12158 25412 12164 25424
rect 11716 25384 12164 25412
rect 4430 25304 4436 25356
rect 4488 25344 4494 25356
rect 4890 25344 4896 25356
rect 4488 25316 4896 25344
rect 4488 25304 4494 25316
rect 4890 25304 4896 25316
rect 4948 25344 4954 25356
rect 11716 25353 11744 25384
rect 12158 25372 12164 25384
rect 12216 25372 12222 25424
rect 5629 25347 5687 25353
rect 5629 25344 5641 25347
rect 4948 25316 5641 25344
rect 4948 25304 4954 25316
rect 5629 25313 5641 25316
rect 5675 25344 5687 25347
rect 7377 25347 7435 25353
rect 7377 25344 7389 25347
rect 5675 25316 7389 25344
rect 5675 25313 5687 25316
rect 5629 25307 5687 25313
rect 7377 25313 7389 25316
rect 7423 25313 7435 25347
rect 7377 25307 7435 25313
rect 11149 25347 11207 25353
rect 11149 25313 11161 25347
rect 11195 25344 11207 25347
rect 11701 25347 11759 25353
rect 11701 25344 11713 25347
rect 11195 25316 11713 25344
rect 11195 25313 11207 25316
rect 11149 25307 11207 25313
rect 11701 25313 11713 25316
rect 11747 25313 11759 25347
rect 11701 25307 11759 25313
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25344 11943 25347
rect 12802 25344 12808 25356
rect 11931 25316 12808 25344
rect 11931 25313 11943 25316
rect 11885 25307 11943 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 13188 25353 13216 25452
rect 21637 25449 21649 25452
rect 21683 25480 21695 25483
rect 22370 25480 22376 25492
rect 21683 25452 22376 25480
rect 21683 25449 21695 25452
rect 21637 25443 21695 25449
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 23106 25480 23112 25492
rect 23067 25452 23112 25480
rect 23106 25440 23112 25452
rect 23164 25440 23170 25492
rect 24121 25483 24179 25489
rect 24121 25449 24133 25483
rect 24167 25480 24179 25483
rect 24302 25480 24308 25492
rect 24167 25452 24308 25480
rect 24167 25449 24179 25452
rect 24121 25443 24179 25449
rect 24302 25440 24308 25452
rect 24360 25440 24366 25492
rect 24762 25480 24768 25492
rect 24412 25452 24768 25480
rect 15289 25415 15347 25421
rect 15289 25381 15301 25415
rect 15335 25412 15347 25415
rect 17402 25412 17408 25424
rect 15335 25384 17408 25412
rect 15335 25381 15347 25384
rect 15289 25375 15347 25381
rect 17402 25372 17408 25384
rect 17460 25372 17466 25424
rect 13173 25347 13231 25353
rect 13173 25313 13185 25347
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 15933 25347 15991 25353
rect 15933 25313 15945 25347
rect 15979 25344 15991 25347
rect 16206 25344 16212 25356
rect 15979 25316 16212 25344
rect 15979 25313 15991 25316
rect 15933 25307 15991 25313
rect 16206 25304 16212 25316
rect 16264 25304 16270 25356
rect 16301 25347 16359 25353
rect 16301 25313 16313 25347
rect 16347 25313 16359 25347
rect 16301 25307 16359 25313
rect 16485 25347 16543 25353
rect 16485 25313 16497 25347
rect 16531 25344 16543 25347
rect 17494 25344 17500 25356
rect 16531 25316 17500 25344
rect 16531 25313 16543 25316
rect 16485 25307 16543 25313
rect 5905 25279 5963 25285
rect 5905 25245 5917 25279
rect 5951 25276 5963 25279
rect 6086 25276 6092 25288
rect 5951 25248 6092 25276
rect 5951 25245 5963 25248
rect 5905 25239 5963 25245
rect 6086 25236 6092 25248
rect 6144 25236 6150 25288
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25276 10931 25279
rect 11054 25276 11060 25288
rect 10919 25248 11060 25276
rect 10919 25245 10931 25248
rect 10873 25239 10931 25245
rect 11054 25236 11060 25248
rect 11112 25236 11118 25288
rect 15838 25276 15844 25288
rect 15799 25248 15844 25276
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 11514 25168 11520 25220
rect 11572 25208 11578 25220
rect 12069 25211 12127 25217
rect 12069 25208 12081 25211
rect 11572 25180 12081 25208
rect 11572 25168 11578 25180
rect 12069 25177 12081 25180
rect 12115 25177 12127 25211
rect 12069 25171 12127 25177
rect 14734 25168 14740 25220
rect 14792 25208 14798 25220
rect 16316 25208 16344 25307
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 18969 25347 19027 25353
rect 18969 25313 18981 25347
rect 19015 25344 19027 25347
rect 19058 25344 19064 25356
rect 19015 25316 19064 25344
rect 19015 25313 19027 25316
rect 18969 25307 19027 25313
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 19199 25347 19257 25353
rect 19199 25313 19211 25347
rect 19245 25344 19257 25347
rect 20990 25344 20996 25356
rect 19245 25316 20996 25344
rect 19245 25313 19257 25316
rect 19199 25307 19257 25313
rect 20990 25304 20996 25316
rect 21048 25304 21054 25356
rect 22370 25344 22376 25356
rect 22331 25316 22376 25344
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 22741 25347 22799 25353
rect 22741 25313 22753 25347
rect 22787 25344 22799 25347
rect 22830 25344 22836 25356
rect 22787 25316 22836 25344
rect 22787 25313 22799 25316
rect 22741 25307 22799 25313
rect 22830 25304 22836 25316
rect 22888 25304 22894 25356
rect 22925 25347 22983 25353
rect 22925 25313 22937 25347
rect 22971 25344 22983 25347
rect 23124 25344 23152 25440
rect 22971 25316 23152 25344
rect 22971 25313 22983 25316
rect 22925 25307 22983 25313
rect 24118 25304 24124 25356
rect 24176 25344 24182 25356
rect 24412 25353 24440 25452
rect 24762 25440 24768 25452
rect 24820 25480 24826 25492
rect 26694 25480 26700 25492
rect 24820 25452 26700 25480
rect 24820 25440 24826 25452
rect 25685 25415 25743 25421
rect 25685 25412 25697 25415
rect 24964 25384 25697 25412
rect 24397 25347 24455 25353
rect 24397 25344 24409 25347
rect 24176 25316 24409 25344
rect 24176 25304 24182 25316
rect 24397 25313 24409 25316
rect 24443 25313 24455 25347
rect 24397 25307 24455 25313
rect 24762 25304 24768 25356
rect 24820 25344 24826 25356
rect 24964 25353 24992 25384
rect 25685 25381 25697 25384
rect 25731 25381 25743 25415
rect 25685 25375 25743 25381
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 24820 25316 24961 25344
rect 24820 25304 24826 25316
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 25130 25344 25136 25356
rect 25091 25316 25136 25344
rect 24949 25307 25007 25313
rect 25130 25304 25136 25316
rect 25188 25304 25194 25356
rect 26528 25353 26556 25452
rect 26694 25440 26700 25452
rect 26752 25440 26758 25492
rect 26513 25347 26571 25353
rect 26513 25313 26525 25347
rect 26559 25313 26571 25347
rect 26513 25307 26571 25313
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25276 19395 25279
rect 19426 25276 19432 25288
rect 19383 25248 19432 25276
rect 19383 25245 19395 25248
rect 19337 25239 19395 25245
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 21726 25276 21732 25288
rect 21687 25248 21732 25276
rect 21726 25236 21732 25248
rect 21784 25236 21790 25288
rect 22462 25276 22468 25288
rect 22423 25248 22468 25276
rect 22462 25236 22468 25248
rect 22520 25236 22526 25288
rect 22848 25276 22876 25304
rect 23201 25279 23259 25285
rect 23201 25276 23213 25279
rect 22848 25248 23213 25276
rect 23201 25245 23213 25248
rect 23247 25245 23259 25279
rect 23201 25239 23259 25245
rect 24026 25236 24032 25288
rect 24084 25276 24090 25288
rect 24302 25276 24308 25288
rect 24084 25248 24308 25276
rect 24084 25236 24090 25248
rect 24302 25236 24308 25248
rect 24360 25236 24366 25288
rect 14792 25180 16344 25208
rect 19134 25211 19192 25217
rect 14792 25168 14798 25180
rect 19134 25177 19146 25211
rect 19180 25208 19192 25211
rect 19180 25180 19380 25208
rect 19180 25177 19192 25180
rect 19134 25171 19192 25177
rect 19352 25152 19380 25180
rect 24688 25180 25544 25208
rect 24688 25152 24716 25180
rect 7190 25140 7196 25152
rect 7151 25112 7196 25140
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 12158 25100 12164 25152
rect 12216 25140 12222 25152
rect 12529 25143 12587 25149
rect 12529 25140 12541 25143
rect 12216 25112 12541 25140
rect 12216 25100 12222 25112
rect 12529 25109 12541 25112
rect 12575 25140 12587 25143
rect 12710 25140 12716 25152
rect 12575 25112 12716 25140
rect 12575 25109 12587 25112
rect 12529 25103 12587 25109
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 13357 25143 13415 25149
rect 13357 25109 13369 25143
rect 13403 25140 13415 25143
rect 13538 25140 13544 25152
rect 13403 25112 13544 25140
rect 13403 25109 13415 25112
rect 13357 25103 13415 25109
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 19334 25100 19340 25152
rect 19392 25100 19398 25152
rect 19610 25140 19616 25152
rect 19571 25112 19616 25140
rect 19610 25100 19616 25112
rect 19668 25100 19674 25152
rect 24670 25100 24676 25152
rect 24728 25100 24734 25152
rect 25406 25140 25412 25152
rect 25367 25112 25412 25140
rect 25406 25100 25412 25112
rect 25464 25100 25470 25152
rect 25516 25140 25544 25180
rect 25958 25168 25964 25220
rect 26016 25208 26022 25220
rect 31754 25208 31760 25220
rect 26016 25180 31760 25208
rect 26016 25168 26022 25180
rect 31754 25168 31760 25180
rect 31812 25168 31818 25220
rect 26697 25143 26755 25149
rect 26697 25140 26709 25143
rect 25516 25112 26709 25140
rect 26697 25109 26709 25112
rect 26743 25109 26755 25143
rect 26697 25103 26755 25109
rect 1104 25050 29256 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 29256 25050
rect 1104 24976 29256 24998
rect 12710 24896 12716 24948
rect 12768 24936 12774 24948
rect 24305 24939 24363 24945
rect 24305 24936 24317 24939
rect 12768 24908 24317 24936
rect 12768 24896 12774 24908
rect 24305 24905 24317 24908
rect 24351 24936 24363 24939
rect 24762 24936 24768 24948
rect 24351 24908 24768 24936
rect 24351 24905 24363 24908
rect 24305 24899 24363 24905
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 31570 24936 31576 24948
rect 25240 24908 31576 24936
rect 7190 24868 7196 24880
rect 7103 24840 7196 24868
rect 7190 24828 7196 24840
rect 7248 24868 7254 24880
rect 18414 24868 18420 24880
rect 7248 24840 18420 24868
rect 7248 24828 7254 24840
rect 18414 24828 18420 24840
rect 18472 24828 18478 24880
rect 19058 24868 19064 24880
rect 19019 24840 19064 24868
rect 19058 24828 19064 24840
rect 19116 24828 19122 24880
rect 21542 24828 21548 24880
rect 21600 24868 21606 24880
rect 25240 24868 25268 24908
rect 31570 24896 31576 24908
rect 31628 24896 31634 24948
rect 21600 24840 25268 24868
rect 21600 24828 21606 24840
rect 26510 24828 26516 24880
rect 26568 24868 26574 24880
rect 31662 24868 31668 24880
rect 26568 24840 31668 24868
rect 26568 24828 26574 24840
rect 31662 24828 31668 24840
rect 31720 24828 31726 24880
rect 6089 24803 6147 24809
rect 6089 24800 6101 24803
rect 5460 24772 6101 24800
rect 4982 24692 4988 24744
rect 5040 24732 5046 24744
rect 5169 24735 5227 24741
rect 5169 24732 5181 24735
rect 5040 24704 5181 24732
rect 5040 24692 5046 24704
rect 5169 24701 5181 24704
rect 5215 24701 5227 24735
rect 5350 24732 5356 24744
rect 5311 24704 5356 24732
rect 5169 24695 5227 24701
rect 5077 24599 5135 24605
rect 5077 24565 5089 24599
rect 5123 24596 5135 24599
rect 5184 24596 5212 24695
rect 5350 24692 5356 24704
rect 5408 24692 5414 24744
rect 5460 24741 5488 24772
rect 6089 24769 6101 24772
rect 6135 24800 6147 24803
rect 19610 24800 19616 24812
rect 6135 24772 19616 24800
rect 6135 24769 6147 24772
rect 6089 24763 6147 24769
rect 19610 24760 19616 24772
rect 19668 24760 19674 24812
rect 25406 24760 25412 24812
rect 25464 24800 25470 24812
rect 25501 24803 25559 24809
rect 25501 24800 25513 24803
rect 25464 24772 25513 24800
rect 25464 24760 25470 24772
rect 25501 24769 25513 24772
rect 25547 24769 25559 24803
rect 25501 24763 25559 24769
rect 5445 24735 5503 24741
rect 5445 24701 5457 24735
rect 5491 24701 5503 24735
rect 5445 24695 5503 24701
rect 6825 24735 6883 24741
rect 6825 24701 6837 24735
rect 6871 24732 6883 24735
rect 7190 24732 7196 24744
rect 6871 24704 7196 24732
rect 6871 24701 6883 24704
rect 6825 24695 6883 24701
rect 7190 24692 7196 24704
rect 7248 24692 7254 24744
rect 12618 24732 12624 24744
rect 12579 24704 12624 24732
rect 12618 24692 12624 24704
rect 12676 24692 12682 24744
rect 12802 24732 12808 24744
rect 12763 24704 12808 24732
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 13357 24735 13415 24741
rect 13357 24701 13369 24735
rect 13403 24732 13415 24735
rect 13538 24732 13544 24744
rect 13403 24704 13544 24732
rect 13403 24701 13415 24704
rect 13357 24695 13415 24701
rect 13538 24692 13544 24704
rect 13596 24692 13602 24744
rect 13633 24735 13691 24741
rect 13633 24701 13645 24735
rect 13679 24701 13691 24735
rect 13633 24695 13691 24701
rect 5902 24664 5908 24676
rect 5863 24636 5908 24664
rect 5902 24624 5908 24636
rect 5960 24624 5966 24676
rect 12636 24664 12664 24692
rect 13648 24664 13676 24695
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 15988 24704 18061 24732
rect 15988 24692 15994 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18414 24732 18420 24744
rect 18375 24704 18420 24732
rect 18049 24695 18107 24701
rect 12636 24636 13676 24664
rect 13909 24667 13967 24673
rect 13909 24633 13921 24667
rect 13955 24664 13967 24667
rect 14458 24664 14464 24676
rect 13955 24636 14464 24664
rect 13955 24633 13967 24636
rect 13909 24627 13967 24633
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 18064 24664 18092 24695
rect 18414 24692 18420 24704
rect 18472 24692 18478 24744
rect 18782 24732 18788 24744
rect 18743 24704 18788 24732
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 19061 24735 19119 24741
rect 19061 24701 19073 24735
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 20257 24735 20315 24741
rect 20257 24701 20269 24735
rect 20303 24732 20315 24735
rect 22738 24732 22744 24744
rect 20303 24704 22744 24732
rect 20303 24701 20315 24704
rect 20257 24695 20315 24701
rect 19076 24664 19104 24695
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 24118 24732 24124 24744
rect 24079 24704 24124 24732
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24732 25191 24735
rect 25225 24735 25283 24741
rect 25225 24732 25237 24735
rect 25179 24704 25237 24732
rect 25179 24701 25191 24704
rect 25133 24695 25191 24701
rect 25225 24701 25237 24704
rect 25271 24732 25283 24735
rect 26142 24732 26148 24744
rect 25271 24704 26148 24732
rect 25271 24701 25283 24704
rect 25225 24695 25283 24701
rect 26142 24692 26148 24704
rect 26200 24692 26206 24744
rect 26878 24664 26884 24676
rect 18064 24636 19104 24664
rect 26839 24636 26884 24664
rect 26878 24624 26884 24636
rect 26936 24624 26942 24676
rect 6178 24596 6184 24608
rect 5123 24568 6184 24596
rect 5123 24565 5135 24568
rect 5077 24559 5135 24565
rect 6178 24556 6184 24568
rect 6236 24556 6242 24608
rect 6914 24596 6920 24608
rect 6875 24568 6920 24596
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 18598 24556 18604 24608
rect 18656 24596 18662 24608
rect 20349 24599 20407 24605
rect 20349 24596 20361 24599
rect 18656 24568 20361 24596
rect 18656 24556 18662 24568
rect 20349 24565 20361 24568
rect 20395 24565 20407 24599
rect 20349 24559 20407 24565
rect 23198 24556 23204 24608
rect 23256 24596 23262 24608
rect 24946 24596 24952 24608
rect 23256 24568 24952 24596
rect 23256 24556 23262 24568
rect 24946 24556 24952 24568
rect 25004 24596 25010 24608
rect 25498 24596 25504 24608
rect 25004 24568 25504 24596
rect 25004 24556 25010 24568
rect 25498 24556 25504 24568
rect 25556 24556 25562 24608
rect 1104 24506 29256 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 29256 24506
rect 1104 24432 29256 24454
rect 6086 24352 6092 24404
rect 6144 24392 6150 24404
rect 6181 24395 6239 24401
rect 6181 24392 6193 24395
rect 6144 24364 6193 24392
rect 6144 24352 6150 24364
rect 6181 24361 6193 24364
rect 6227 24361 6239 24395
rect 6181 24355 6239 24361
rect 18414 24352 18420 24404
rect 18472 24392 18478 24404
rect 25130 24392 25136 24404
rect 18472 24364 25136 24392
rect 18472 24352 18478 24364
rect 25130 24352 25136 24364
rect 25188 24392 25194 24404
rect 26605 24395 26663 24401
rect 26605 24392 26617 24395
rect 25188 24364 26617 24392
rect 25188 24352 25194 24364
rect 26605 24361 26617 24364
rect 26651 24361 26663 24395
rect 26605 24355 26663 24361
rect 18693 24327 18751 24333
rect 18693 24293 18705 24327
rect 18739 24324 18751 24327
rect 19426 24324 19432 24336
rect 18739 24296 19432 24324
rect 18739 24293 18751 24296
rect 18693 24287 18751 24293
rect 19426 24284 19432 24296
rect 19484 24284 19490 24336
rect 22462 24284 22468 24336
rect 22520 24324 22526 24336
rect 24670 24324 24676 24336
rect 22520 24296 23888 24324
rect 22520 24284 22526 24296
rect 5169 24259 5227 24265
rect 5169 24225 5181 24259
rect 5215 24256 5227 24259
rect 5626 24256 5632 24268
rect 5215 24228 5632 24256
rect 5215 24225 5227 24228
rect 5169 24219 5227 24225
rect 5626 24216 5632 24228
rect 5684 24256 5690 24268
rect 5721 24259 5779 24265
rect 5721 24256 5733 24259
rect 5684 24228 5733 24256
rect 5684 24216 5690 24228
rect 5721 24225 5733 24228
rect 5767 24225 5779 24259
rect 5721 24219 5779 24225
rect 5905 24259 5963 24265
rect 5905 24225 5917 24259
rect 5951 24256 5963 24259
rect 6914 24256 6920 24268
rect 5951 24228 6920 24256
rect 5951 24225 5963 24228
rect 5905 24219 5963 24225
rect 6914 24216 6920 24228
rect 6972 24216 6978 24268
rect 11514 24256 11520 24268
rect 11475 24228 11520 24256
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 17494 24216 17500 24268
rect 17552 24256 17558 24268
rect 18233 24259 18291 24265
rect 18233 24256 18245 24259
rect 17552 24228 18245 24256
rect 17552 24216 17558 24228
rect 18233 24225 18245 24228
rect 18279 24225 18291 24259
rect 18233 24219 18291 24225
rect 23109 24259 23167 24265
rect 23109 24225 23121 24259
rect 23155 24256 23167 24259
rect 23198 24256 23204 24268
rect 23155 24228 23204 24256
rect 23155 24225 23167 24228
rect 23109 24219 23167 24225
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 23860 24265 23888 24296
rect 23952 24296 24676 24324
rect 23952 24268 23980 24296
rect 24670 24284 24676 24296
rect 24728 24284 24734 24336
rect 23385 24259 23443 24265
rect 23385 24225 23397 24259
rect 23431 24256 23443 24259
rect 23845 24259 23903 24265
rect 23431 24228 23612 24256
rect 23431 24225 23443 24228
rect 23385 24219 23443 24225
rect 3326 24148 3332 24200
rect 3384 24188 3390 24200
rect 4062 24188 4068 24200
rect 3384 24160 4068 24188
rect 3384 24148 3390 24160
rect 4062 24148 4068 24160
rect 4120 24148 4126 24200
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4816 24160 4997 24188
rect 4816 24064 4844 24160
rect 4985 24157 4997 24160
rect 5031 24157 5043 24191
rect 11241 24191 11299 24197
rect 11241 24188 11253 24191
rect 4985 24151 5043 24157
rect 11164 24160 11253 24188
rect 11164 24064 11192 24160
rect 11241 24157 11253 24160
rect 11287 24157 11299 24191
rect 11241 24151 11299 24157
rect 18046 24148 18052 24200
rect 18104 24188 18110 24200
rect 18141 24191 18199 24197
rect 18141 24188 18153 24191
rect 18104 24160 18153 24188
rect 18104 24148 18110 24160
rect 18141 24157 18153 24160
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19426 24188 19432 24200
rect 18840 24160 19432 24188
rect 18840 24148 18846 24160
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 13538 24080 13544 24132
rect 13596 24120 13602 24132
rect 18800 24120 18828 24148
rect 13596 24092 18828 24120
rect 13596 24080 13602 24092
rect 4798 24052 4804 24064
rect 4759 24024 4804 24052
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 11146 24052 11152 24064
rect 11107 24024 11152 24052
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 12710 24012 12716 24064
rect 12768 24052 12774 24064
rect 12805 24055 12863 24061
rect 12805 24052 12817 24055
rect 12768 24024 12817 24052
rect 12768 24012 12774 24024
rect 12805 24021 12817 24024
rect 12851 24021 12863 24055
rect 23584 24052 23612 24228
rect 23845 24225 23857 24259
rect 23891 24225 23903 24259
rect 23845 24219 23903 24225
rect 23934 24216 23940 24268
rect 23992 24256 23998 24268
rect 23992 24228 24085 24256
rect 23992 24216 23998 24228
rect 24578 24216 24584 24268
rect 24636 24256 24642 24268
rect 24857 24259 24915 24265
rect 24857 24256 24869 24259
rect 24636 24228 24869 24256
rect 24636 24216 24642 24228
rect 24857 24225 24869 24228
rect 24903 24225 24915 24259
rect 24857 24219 24915 24225
rect 26513 24259 26571 24265
rect 26513 24225 26525 24259
rect 26559 24256 26571 24259
rect 26878 24256 26884 24268
rect 26559 24228 26884 24256
rect 26559 24225 26571 24228
rect 26513 24219 26571 24225
rect 26878 24216 26884 24228
rect 26936 24216 26942 24268
rect 24118 24080 24124 24132
rect 24176 24120 24182 24132
rect 24305 24123 24363 24129
rect 24305 24120 24317 24123
rect 24176 24092 24317 24120
rect 24176 24080 24182 24092
rect 24305 24089 24317 24092
rect 24351 24089 24363 24123
rect 24305 24083 24363 24089
rect 24578 24052 24584 24064
rect 23584 24024 24584 24052
rect 12805 24015 12863 24021
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 26878 24052 26884 24064
rect 26839 24024 26884 24052
rect 26878 24012 26884 24024
rect 26936 24012 26942 24064
rect 27430 24012 27436 24064
rect 27488 24052 27494 24064
rect 28905 24055 28963 24061
rect 28905 24052 28917 24055
rect 27488 24024 28917 24052
rect 27488 24012 27494 24024
rect 28905 24021 28917 24024
rect 28951 24052 28963 24055
rect 31570 24052 31576 24064
rect 28951 24024 31576 24052
rect 28951 24021 28963 24024
rect 28905 24015 28963 24021
rect 31570 24012 31576 24024
rect 31628 24012 31634 24064
rect 1104 23962 29256 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 29256 23962
rect 1104 23888 29256 23910
rect 4062 23808 4068 23860
rect 4120 23848 4126 23860
rect 32214 23848 32220 23860
rect 4120 23820 32220 23848
rect 4120 23808 4126 23820
rect 32214 23808 32220 23820
rect 32272 23808 32278 23860
rect 12802 23740 12808 23792
rect 12860 23780 12866 23792
rect 12897 23783 12955 23789
rect 12897 23780 12909 23783
rect 12860 23752 12909 23780
rect 12860 23740 12866 23752
rect 12897 23749 12909 23752
rect 12943 23749 12955 23783
rect 12897 23743 12955 23749
rect 13906 23740 13912 23792
rect 13964 23780 13970 23792
rect 16298 23780 16304 23792
rect 13964 23752 16304 23780
rect 13964 23740 13970 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 4249 23715 4307 23721
rect 4249 23681 4261 23715
rect 4295 23712 4307 23715
rect 4890 23712 4896 23724
rect 4295 23684 4896 23712
rect 4295 23681 4307 23684
rect 4249 23675 4307 23681
rect 4890 23672 4896 23684
rect 4948 23712 4954 23724
rect 5997 23715 6055 23721
rect 5997 23712 6009 23715
rect 4948 23684 6009 23712
rect 4948 23672 4954 23684
rect 5997 23681 6009 23684
rect 6043 23681 6055 23715
rect 15194 23712 15200 23724
rect 15155 23684 15200 23712
rect 5997 23675 6055 23681
rect 15194 23672 15200 23684
rect 15252 23672 15258 23724
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 19429 23715 19487 23721
rect 19429 23712 19441 23715
rect 19392 23684 19441 23712
rect 19392 23672 19398 23684
rect 19429 23681 19441 23684
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23712 25835 23715
rect 26510 23712 26516 23724
rect 25823 23684 26516 23712
rect 25823 23681 25835 23684
rect 25777 23675 25835 23681
rect 26510 23672 26516 23684
rect 26568 23672 26574 23724
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 4062 23644 4068 23656
rect 3476 23616 4068 23644
rect 3476 23604 3482 23616
rect 4062 23604 4068 23616
rect 4120 23604 4126 23656
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23644 4583 23647
rect 5534 23644 5540 23656
rect 4571 23616 5540 23644
rect 4571 23613 4583 23616
rect 4525 23607 4583 23613
rect 5534 23604 5540 23616
rect 5592 23604 5598 23656
rect 5905 23647 5963 23653
rect 5905 23613 5917 23647
rect 5951 23644 5963 23647
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 5951 23616 6837 23644
rect 5951 23613 5963 23616
rect 5905 23607 5963 23613
rect 6825 23613 6837 23616
rect 6871 23644 6883 23647
rect 6871 23616 7236 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 7208 23585 7236 23616
rect 12710 23604 12716 23656
rect 12768 23644 12774 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12768 23616 12817 23644
rect 12768 23604 12774 23616
rect 12805 23613 12817 23616
rect 12851 23613 12863 23647
rect 13906 23644 13912 23656
rect 13867 23616 13912 23644
rect 12805 23607 12863 23613
rect 13906 23604 13912 23616
rect 13964 23604 13970 23656
rect 14274 23644 14280 23656
rect 14235 23616 14280 23644
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 14458 23644 14464 23656
rect 14419 23616 14464 23644
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 14737 23647 14795 23653
rect 14737 23613 14749 23647
rect 14783 23644 14795 23647
rect 14826 23644 14832 23656
rect 14783 23616 14832 23644
rect 14783 23613 14795 23616
rect 14737 23607 14795 23613
rect 7193 23579 7251 23585
rect 7193 23545 7205 23579
rect 7239 23576 7251 23579
rect 13814 23576 13820 23588
rect 7239 23548 13676 23576
rect 13727 23548 13820 23576
rect 7239 23545 7251 23548
rect 7193 23539 7251 23545
rect 3050 23468 3056 23520
rect 3108 23508 3114 23520
rect 3694 23508 3700 23520
rect 3108 23480 3700 23508
rect 3108 23468 3114 23480
rect 3694 23468 3700 23480
rect 3752 23468 3758 23520
rect 6086 23468 6092 23520
rect 6144 23508 6150 23520
rect 6917 23511 6975 23517
rect 6917 23508 6929 23511
rect 6144 23480 6929 23508
rect 6144 23468 6150 23480
rect 6917 23477 6929 23480
rect 6963 23477 6975 23511
rect 12710 23508 12716 23520
rect 12671 23480 12716 23508
rect 6917 23471 6975 23477
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 13648 23508 13676 23548
rect 13814 23536 13820 23548
rect 13872 23576 13878 23588
rect 14752 23576 14780 23607
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 14921 23647 14979 23653
rect 14921 23613 14933 23647
rect 14967 23644 14979 23647
rect 15102 23644 15108 23656
rect 14967 23616 15108 23644
rect 14967 23613 14979 23616
rect 14921 23607 14979 23613
rect 15102 23604 15108 23616
rect 15160 23604 15166 23656
rect 18877 23647 18935 23653
rect 18877 23644 18889 23647
rect 18708 23616 18889 23644
rect 13872 23548 14780 23576
rect 13872 23536 13878 23548
rect 18708 23517 18736 23616
rect 18877 23613 18889 23616
rect 18923 23613 18935 23647
rect 18877 23607 18935 23613
rect 18966 23604 18972 23656
rect 19024 23644 19030 23656
rect 24121 23647 24179 23653
rect 19024 23616 19069 23644
rect 19024 23604 19030 23616
rect 24121 23613 24133 23647
rect 24167 23613 24179 23647
rect 24394 23644 24400 23656
rect 24355 23616 24400 23644
rect 24121 23607 24179 23613
rect 18693 23511 18751 23517
rect 18693 23508 18705 23511
rect 13648 23480 18705 23508
rect 18693 23477 18705 23480
rect 18739 23508 18751 23511
rect 18782 23508 18788 23520
rect 18739 23480 18788 23508
rect 18739 23477 18751 23480
rect 18693 23471 18751 23477
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 24029 23511 24087 23517
rect 24029 23477 24041 23511
rect 24075 23508 24087 23511
rect 24136 23508 24164 23607
rect 24394 23604 24400 23616
rect 24452 23604 24458 23656
rect 24210 23508 24216 23520
rect 24075 23480 24216 23508
rect 24075 23477 24087 23480
rect 24029 23471 24087 23477
rect 24210 23468 24216 23480
rect 24268 23468 24274 23520
rect 1104 23418 29256 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 29256 23418
rect 1104 23344 29256 23366
rect 4798 23264 4804 23316
rect 4856 23304 4862 23316
rect 4856 23276 6224 23304
rect 4856 23264 4862 23276
rect 5626 23236 5632 23248
rect 4540 23208 5632 23236
rect 4540 23177 4568 23208
rect 5626 23196 5632 23208
rect 5684 23196 5690 23248
rect 4510 23171 4568 23177
rect 4510 23137 4522 23171
rect 4556 23137 4568 23171
rect 5074 23168 5080 23180
rect 5035 23140 5080 23168
rect 4510 23131 4568 23137
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 5261 23171 5319 23177
rect 5261 23137 5273 23171
rect 5307 23168 5319 23171
rect 6086 23168 6092 23180
rect 5307 23140 6092 23168
rect 5307 23137 5319 23140
rect 5261 23131 5319 23137
rect 6086 23128 6092 23140
rect 6144 23128 6150 23180
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 5534 23100 5540 23112
rect 5495 23072 5540 23100
rect 4341 23063 4399 23069
rect 3418 22924 3424 22976
rect 3476 22964 3482 22976
rect 4249 22967 4307 22973
rect 4249 22964 4261 22967
rect 3476 22936 4261 22964
rect 3476 22924 3482 22936
rect 4249 22933 4261 22936
rect 4295 22964 4307 22967
rect 4356 22964 4384 23063
rect 5534 23060 5540 23072
rect 5592 23060 5598 23112
rect 6196 23032 6224 23276
rect 12618 23264 12624 23316
rect 12676 23304 12682 23316
rect 12805 23307 12863 23313
rect 12805 23304 12817 23307
rect 12676 23276 12817 23304
rect 12676 23264 12682 23276
rect 12805 23273 12817 23276
rect 12851 23304 12863 23307
rect 13722 23304 13728 23316
rect 12851 23276 13728 23304
rect 12851 23273 12863 23276
rect 12805 23267 12863 23273
rect 13722 23264 13728 23276
rect 13780 23264 13786 23316
rect 22462 23264 22468 23316
rect 22520 23304 22526 23316
rect 22649 23307 22707 23313
rect 22649 23304 22661 23307
rect 22520 23276 22661 23304
rect 22520 23264 22526 23276
rect 22649 23273 22661 23276
rect 22695 23273 22707 23307
rect 22649 23267 22707 23273
rect 24394 23264 24400 23316
rect 24452 23304 24458 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24452 23276 24777 23304
rect 24452 23264 24458 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 9493 23239 9551 23245
rect 9493 23205 9505 23239
rect 9539 23236 9551 23239
rect 24026 23236 24032 23248
rect 9539 23208 24032 23236
rect 9539 23205 9551 23208
rect 9493 23199 9551 23205
rect 24026 23196 24032 23208
rect 24084 23196 24090 23248
rect 26605 23239 26663 23245
rect 26605 23236 26617 23239
rect 24504 23208 26617 23236
rect 13538 23168 13544 23180
rect 13499 23140 13544 23168
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 13722 23128 13728 23180
rect 13780 23168 13786 23180
rect 13817 23171 13875 23177
rect 13817 23168 13829 23171
rect 13780 23140 13829 23168
rect 13780 23128 13786 23140
rect 13817 23137 13829 23140
rect 13863 23137 13875 23171
rect 13817 23131 13875 23137
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23168 14151 23171
rect 14274 23168 14280 23180
rect 14139 23140 14280 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 17494 23128 17500 23180
rect 17552 23168 17558 23180
rect 17681 23171 17739 23177
rect 17681 23168 17693 23171
rect 17552 23140 17693 23168
rect 17552 23128 17558 23140
rect 17681 23137 17693 23140
rect 17727 23137 17739 23171
rect 17681 23131 17739 23137
rect 22557 23171 22615 23177
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 22925 23171 22983 23177
rect 22925 23168 22937 23171
rect 22603 23140 22937 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 22925 23137 22937 23140
rect 22971 23168 22983 23171
rect 23753 23171 23811 23177
rect 22971 23140 23704 23168
rect 22971 23137 22983 23140
rect 22925 23131 22983 23137
rect 13170 23100 13176 23112
rect 13131 23072 13176 23100
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 13832 23072 23397 23100
rect 13832 23032 13860 23072
rect 23385 23069 23397 23072
rect 23431 23100 23443 23103
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 23431 23072 23581 23100
rect 23431 23069 23443 23072
rect 23385 23063 23443 23069
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 6196 23004 13860 23032
rect 13906 22992 13912 23044
rect 13964 23032 13970 23044
rect 18138 23032 18144 23044
rect 13964 23004 18144 23032
rect 13964 22992 13970 23004
rect 18138 22992 18144 23004
rect 18196 22992 18202 23044
rect 9493 22967 9551 22973
rect 9493 22964 9505 22967
rect 4295 22936 9505 22964
rect 4295 22933 4307 22936
rect 4249 22927 4307 22933
rect 9493 22933 9505 22936
rect 9539 22933 9551 22967
rect 17862 22964 17868 22976
rect 17823 22936 17868 22964
rect 9493 22927 9551 22933
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 23584 22964 23612 23063
rect 23676 23032 23704 23140
rect 23753 23137 23765 23171
rect 23799 23168 23811 23171
rect 24302 23168 24308 23180
rect 23799 23140 24308 23168
rect 23799 23137 23811 23140
rect 23753 23131 23811 23137
rect 24302 23128 24308 23140
rect 24360 23128 24366 23180
rect 24504 23177 24532 23208
rect 26605 23205 26617 23208
rect 26651 23205 26663 23239
rect 26605 23199 26663 23205
rect 24489 23171 24547 23177
rect 24489 23137 24501 23171
rect 24535 23137 24547 23171
rect 26510 23168 26516 23180
rect 26471 23140 26516 23168
rect 24489 23131 24547 23137
rect 26510 23128 26516 23140
rect 26568 23128 26574 23180
rect 25406 23032 25412 23044
rect 23676 23004 25412 23032
rect 25406 22992 25412 23004
rect 25464 22992 25470 23044
rect 26234 22964 26240 22976
rect 23584 22936 26240 22964
rect 26234 22924 26240 22936
rect 26292 22924 26298 22976
rect 1104 22874 29256 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 29256 22874
rect 1104 22800 29256 22822
rect 8478 22720 8484 22772
rect 8536 22760 8542 22772
rect 8849 22763 8907 22769
rect 8849 22760 8861 22763
rect 8536 22732 8861 22760
rect 8536 22720 8542 22732
rect 8849 22729 8861 22732
rect 8895 22760 8907 22763
rect 9306 22760 9312 22772
rect 8895 22732 9312 22760
rect 8895 22729 8907 22732
rect 8849 22723 8907 22729
rect 9306 22720 9312 22732
rect 9364 22760 9370 22772
rect 13814 22760 13820 22772
rect 9364 22732 13820 22760
rect 9364 22720 9370 22732
rect 13814 22720 13820 22732
rect 13872 22720 13878 22772
rect 17862 22760 17868 22772
rect 17823 22732 17868 22760
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 20625 22763 20683 22769
rect 20625 22760 20637 22763
rect 18248 22732 20637 22760
rect 5074 22692 5080 22704
rect 3068 22664 5080 22692
rect 2593 22627 2651 22633
rect 2593 22593 2605 22627
rect 2639 22624 2651 22627
rect 2777 22627 2835 22633
rect 2777 22624 2789 22627
rect 2639 22596 2789 22624
rect 2639 22593 2651 22596
rect 2593 22587 2651 22593
rect 2777 22593 2789 22596
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 2792 22488 2820 22587
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 3068 22556 3096 22664
rect 5074 22652 5080 22664
rect 5132 22652 5138 22704
rect 8386 22652 8392 22704
rect 8444 22692 8450 22704
rect 15105 22695 15163 22701
rect 15105 22692 15117 22695
rect 8444 22664 15117 22692
rect 8444 22652 8450 22664
rect 15105 22661 15117 22664
rect 15151 22661 15163 22695
rect 15105 22655 15163 22661
rect 13538 22584 13544 22636
rect 13596 22624 13602 22636
rect 18248 22633 18276 22732
rect 20625 22729 20637 22732
rect 20671 22729 20683 22763
rect 20625 22723 20683 22729
rect 13633 22627 13691 22633
rect 13633 22624 13645 22627
rect 13596 22596 13645 22624
rect 13596 22584 13602 22596
rect 13633 22593 13645 22596
rect 13679 22624 13691 22627
rect 18233 22627 18291 22633
rect 13679 22596 14596 22624
rect 13679 22593 13691 22596
rect 13633 22587 13691 22593
rect 14568 22568 14596 22596
rect 18233 22593 18245 22627
rect 18279 22593 18291 22627
rect 23385 22627 23443 22633
rect 18233 22587 18291 22593
rect 18524 22596 18828 22624
rect 3421 22559 3479 22565
rect 3421 22556 3433 22559
rect 2915 22528 3433 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 3421 22525 3433 22528
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22556 3663 22559
rect 4154 22556 4160 22568
rect 3651 22528 4160 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 4154 22516 4160 22528
rect 4212 22516 4218 22568
rect 8478 22556 8484 22568
rect 8439 22528 8484 22556
rect 8478 22516 8484 22528
rect 8536 22516 8542 22568
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22556 13783 22559
rect 13906 22556 13912 22568
rect 13771 22528 13912 22556
rect 13771 22525 13783 22528
rect 13725 22519 13783 22525
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 14090 22556 14096 22568
rect 14051 22528 14096 22556
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 14274 22556 14280 22568
rect 14235 22528 14280 22556
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 14550 22556 14556 22568
rect 14511 22528 14556 22556
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 14737 22559 14795 22565
rect 14737 22525 14749 22559
rect 14783 22556 14795 22559
rect 15102 22556 15108 22568
rect 14783 22528 15108 22556
rect 14783 22525 14795 22528
rect 14737 22519 14795 22525
rect 15102 22516 15108 22528
rect 15160 22516 15166 22568
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18524 22556 18552 22596
rect 17920 22528 18552 22556
rect 18601 22559 18659 22565
rect 17920 22516 17926 22528
rect 18601 22525 18613 22559
rect 18647 22556 18659 22559
rect 18690 22556 18696 22568
rect 18647 22528 18696 22556
rect 18647 22525 18659 22528
rect 18601 22519 18659 22525
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 18800 22565 18828 22596
rect 23385 22593 23397 22627
rect 23431 22624 23443 22627
rect 23431 22596 24072 22624
rect 23431 22593 23443 22596
rect 23385 22587 23443 22593
rect 24044 22568 24072 22596
rect 18785 22559 18843 22565
rect 18785 22525 18797 22559
rect 18831 22525 18843 22559
rect 18966 22556 18972 22568
rect 18927 22528 18972 22556
rect 18785 22519 18843 22525
rect 18966 22516 18972 22528
rect 19024 22516 19030 22568
rect 19058 22516 19064 22568
rect 19116 22556 19122 22568
rect 19153 22559 19211 22565
rect 19153 22556 19165 22559
rect 19116 22528 19165 22556
rect 19116 22516 19122 22528
rect 19153 22525 19165 22528
rect 19199 22525 19211 22559
rect 19153 22519 19211 22525
rect 20533 22559 20591 22565
rect 20533 22525 20545 22559
rect 20579 22556 20591 22559
rect 23474 22556 23480 22568
rect 20579 22528 23480 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 23474 22516 23480 22528
rect 23532 22516 23538 22568
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 23937 22559 23995 22565
rect 23937 22556 23949 22559
rect 23900 22528 23949 22556
rect 23900 22516 23906 22528
rect 23937 22525 23949 22528
rect 23983 22525 23995 22559
rect 23937 22519 23995 22525
rect 3786 22488 3792 22500
rect 2792 22460 3792 22488
rect 3786 22448 3792 22460
rect 3844 22448 3850 22500
rect 8754 22448 8760 22500
rect 8812 22488 8818 22500
rect 19705 22491 19763 22497
rect 19705 22488 19717 22491
rect 8812 22460 19717 22488
rect 8812 22448 8818 22460
rect 19705 22457 19717 22460
rect 19751 22457 19763 22491
rect 23952 22488 23980 22519
rect 24026 22516 24032 22568
rect 24084 22556 24090 22568
rect 24489 22559 24547 22565
rect 24084 22528 24129 22556
rect 24084 22516 24090 22528
rect 24489 22525 24501 22559
rect 24535 22525 24547 22559
rect 24489 22519 24547 22525
rect 24673 22559 24731 22565
rect 24673 22525 24685 22559
rect 24719 22525 24731 22559
rect 25958 22556 25964 22568
rect 25919 22528 25964 22556
rect 24673 22519 24731 22525
rect 24302 22488 24308 22500
rect 23952 22460 24308 22488
rect 19705 22451 19763 22457
rect 24302 22448 24308 22460
rect 24360 22488 24366 22500
rect 24504 22488 24532 22519
rect 24360 22460 24532 22488
rect 24688 22488 24716 22519
rect 25958 22516 25964 22528
rect 26016 22516 26022 22568
rect 26053 22491 26111 22497
rect 26053 22488 26065 22491
rect 24688 22460 26065 22488
rect 24360 22448 24366 22460
rect 26053 22457 26065 22460
rect 26099 22457 26111 22491
rect 26053 22451 26111 22457
rect 3878 22420 3884 22432
rect 3839 22392 3884 22420
rect 3878 22380 3884 22392
rect 3936 22380 3942 22432
rect 8570 22420 8576 22432
rect 8531 22392 8576 22420
rect 8570 22380 8576 22392
rect 8628 22380 8634 22432
rect 18141 22423 18199 22429
rect 18141 22389 18153 22423
rect 18187 22420 18199 22423
rect 18966 22420 18972 22432
rect 18187 22392 18972 22420
rect 18187 22389 18199 22392
rect 18141 22383 18199 22389
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 24949 22423 25007 22429
rect 24949 22420 24961 22423
rect 24912 22392 24961 22420
rect 24912 22380 24918 22392
rect 24949 22389 24961 22392
rect 24995 22389 25007 22423
rect 24949 22383 25007 22389
rect 1104 22330 29256 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 29256 22330
rect 1104 22256 29256 22278
rect 8018 22216 8024 22228
rect 7979 22188 8024 22216
rect 8018 22176 8024 22188
rect 8076 22176 8082 22228
rect 13081 22219 13139 22225
rect 13081 22216 13093 22219
rect 12912 22188 13093 22216
rect 12912 22157 12940 22188
rect 13081 22185 13093 22188
rect 13127 22185 13139 22219
rect 19058 22216 19064 22228
rect 13081 22179 13139 22185
rect 18248 22188 19064 22216
rect 12897 22151 12955 22157
rect 12897 22148 12909 22151
rect 12268 22120 12909 22148
rect 4065 22083 4123 22089
rect 4065 22049 4077 22083
rect 4111 22049 4123 22083
rect 4065 22043 4123 22049
rect 4080 22012 4108 22043
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 4212 22052 4257 22080
rect 4212 22040 4218 22052
rect 5074 22040 5080 22092
rect 5132 22080 5138 22092
rect 7009 22083 7067 22089
rect 7009 22080 7021 22083
rect 5132 22052 7021 22080
rect 5132 22040 5138 22052
rect 7009 22049 7021 22052
rect 7055 22080 7067 22083
rect 7561 22083 7619 22089
rect 7561 22080 7573 22083
rect 7055 22052 7573 22080
rect 7055 22049 7067 22052
rect 7009 22043 7067 22049
rect 7561 22049 7573 22052
rect 7607 22049 7619 22083
rect 7561 22043 7619 22049
rect 7745 22083 7803 22089
rect 7745 22049 7757 22083
rect 7791 22080 7803 22083
rect 8570 22080 8576 22092
rect 7791 22052 8576 22080
rect 7791 22049 7803 22052
rect 7745 22043 7803 22049
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 11609 22083 11667 22089
rect 11609 22049 11621 22083
rect 11655 22080 11667 22083
rect 12158 22080 12164 22092
rect 11655 22052 12164 22080
rect 11655 22049 11667 22052
rect 11609 22043 11667 22049
rect 12158 22040 12164 22052
rect 12216 22080 12222 22092
rect 12268 22080 12296 22120
rect 12897 22117 12909 22120
rect 12943 22117 12955 22151
rect 13170 22148 13176 22160
rect 12897 22111 12955 22117
rect 13096 22120 13176 22148
rect 12216 22052 12296 22080
rect 12345 22083 12403 22089
rect 12216 22040 12222 22052
rect 12345 22049 12357 22083
rect 12391 22080 12403 22083
rect 13096 22080 13124 22120
rect 13170 22108 13176 22120
rect 13228 22148 13234 22160
rect 13725 22151 13783 22157
rect 13725 22148 13737 22151
rect 13228 22120 13737 22148
rect 13228 22108 13234 22120
rect 13725 22117 13737 22120
rect 13771 22117 13783 22151
rect 13725 22111 13783 22117
rect 12391 22052 13124 22080
rect 13633 22083 13691 22089
rect 12391 22049 12403 22052
rect 12345 22043 12403 22049
rect 13633 22049 13645 22083
rect 13679 22080 13691 22083
rect 14090 22080 14096 22092
rect 13679 22052 14096 22080
rect 13679 22049 13691 22052
rect 13633 22043 13691 22049
rect 14090 22040 14096 22052
rect 14148 22040 14154 22092
rect 15565 22083 15623 22089
rect 15565 22049 15577 22083
rect 15611 22080 15623 22083
rect 18248 22080 18276 22188
rect 19058 22176 19064 22188
rect 19116 22216 19122 22228
rect 19116 22188 19288 22216
rect 19116 22176 19122 22188
rect 18800 22120 19012 22148
rect 15611 22052 18276 22080
rect 18325 22083 18383 22089
rect 15611 22049 15623 22052
rect 15565 22043 15623 22049
rect 18325 22049 18337 22083
rect 18371 22080 18383 22083
rect 18598 22080 18604 22092
rect 18371 22052 18604 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 18800 22080 18828 22120
rect 18739 22052 18828 22080
rect 18877 22083 18935 22089
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 18877 22049 18889 22083
rect 18923 22049 18935 22083
rect 18877 22043 18935 22049
rect 6825 22015 6883 22021
rect 6825 22012 6837 22015
rect 4080 21984 4476 22012
rect 4448 21885 4476 21984
rect 6656 21984 6837 22012
rect 6656 21944 6684 21984
rect 6825 21981 6837 21984
rect 6871 21981 6883 22015
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 6825 21975 6883 21981
rect 11256 21984 11437 22012
rect 11054 21944 11060 21956
rect 6656 21916 11060 21944
rect 4433 21879 4491 21885
rect 4433 21845 4445 21879
rect 4479 21876 4491 21879
rect 4614 21876 4620 21888
rect 4479 21848 4620 21876
rect 4479 21845 4491 21848
rect 4433 21839 4491 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 6656 21885 6684 21916
rect 11054 21904 11060 21916
rect 11112 21904 11118 21956
rect 11256 21944 11284 21984
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 18892 22012 18920 22043
rect 17920 21984 18920 22012
rect 18984 22012 19012 22120
rect 19150 22080 19156 22092
rect 19111 22052 19156 22080
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19260 22089 19288 22188
rect 23658 22176 23664 22228
rect 23716 22216 23722 22228
rect 31570 22216 31576 22228
rect 23716 22188 31576 22216
rect 23716 22176 23722 22188
rect 31570 22176 31576 22188
rect 31628 22176 31634 22228
rect 19245 22083 19303 22089
rect 19245 22049 19257 22083
rect 19291 22049 19303 22083
rect 24118 22080 24124 22092
rect 24079 22052 24124 22080
rect 19245 22043 19303 22049
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 21174 22012 21180 22024
rect 18984 21984 21180 22012
rect 17920 21972 17926 21984
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 17954 21944 17960 21956
rect 11256 21916 17960 21944
rect 6641 21879 6699 21885
rect 6641 21876 6653 21879
rect 6604 21848 6653 21876
rect 6604 21836 6610 21848
rect 6641 21845 6653 21848
rect 6687 21845 6699 21879
rect 6641 21839 6699 21845
rect 7466 21836 7472 21888
rect 7524 21876 7530 21888
rect 11256 21885 11284 21916
rect 17954 21904 17960 21916
rect 18012 21904 18018 21956
rect 18049 21947 18107 21953
rect 18049 21913 18061 21947
rect 18095 21944 18107 21947
rect 19150 21944 19156 21956
rect 18095 21916 19156 21944
rect 18095 21913 18107 21916
rect 18049 21907 18107 21913
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 11241 21879 11299 21885
rect 11241 21876 11253 21879
rect 7524 21848 11253 21876
rect 7524 21836 7530 21848
rect 11241 21845 11253 21848
rect 11287 21845 11299 21879
rect 11241 21839 11299 21845
rect 12621 21879 12679 21885
rect 12621 21845 12633 21879
rect 12667 21876 12679 21879
rect 12710 21876 12716 21888
rect 12667 21848 12716 21876
rect 12667 21845 12679 21848
rect 12621 21839 12679 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 14001 21879 14059 21885
rect 14001 21845 14013 21879
rect 14047 21876 14059 21879
rect 14090 21876 14096 21888
rect 14047 21848 14096 21876
rect 14047 21845 14059 21848
rect 14001 21839 14059 21845
rect 14090 21836 14096 21848
rect 14148 21836 14154 21888
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 15749 21879 15807 21885
rect 15749 21876 15761 21879
rect 15160 21848 15761 21876
rect 15160 21836 15166 21848
rect 15749 21845 15761 21848
rect 15795 21845 15807 21879
rect 15749 21839 15807 21845
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 18141 21879 18199 21885
rect 18141 21876 18153 21879
rect 17920 21848 18153 21876
rect 17920 21836 17926 21848
rect 18141 21845 18153 21848
rect 18187 21845 18199 21879
rect 18141 21839 18199 21845
rect 18230 21836 18236 21888
rect 18288 21876 18294 21888
rect 19705 21879 19763 21885
rect 19705 21876 19717 21879
rect 18288 21848 19717 21876
rect 18288 21836 18294 21848
rect 19705 21845 19717 21848
rect 19751 21845 19763 21879
rect 19705 21839 19763 21845
rect 23753 21879 23811 21885
rect 23753 21845 23765 21879
rect 23799 21876 23811 21879
rect 23860 21876 23888 21975
rect 24210 21876 24216 21888
rect 23799 21848 24216 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 24210 21836 24216 21848
rect 24268 21836 24274 21888
rect 25406 21876 25412 21888
rect 25367 21848 25412 21876
rect 25406 21836 25412 21848
rect 25464 21836 25470 21888
rect 1104 21786 29256 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 29256 21786
rect 1104 21712 29256 21734
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5813 21675 5871 21681
rect 5813 21672 5825 21675
rect 5132 21644 5825 21672
rect 5132 21632 5138 21644
rect 5813 21641 5825 21644
rect 5859 21641 5871 21675
rect 9306 21672 9312 21684
rect 5813 21635 5871 21641
rect 6288 21644 8800 21672
rect 9267 21644 9312 21672
rect 4341 21607 4399 21613
rect 4341 21573 4353 21607
rect 4387 21604 4399 21607
rect 4614 21604 4620 21616
rect 4387 21576 4620 21604
rect 4387 21573 4399 21576
rect 4341 21567 4399 21573
rect 4614 21564 4620 21576
rect 4672 21604 4678 21616
rect 6288 21604 6316 21644
rect 4672 21576 6316 21604
rect 8772 21604 8800 21644
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 13538 21672 13544 21684
rect 9416 21644 13544 21672
rect 9416 21604 9444 21644
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 21358 21672 21364 21684
rect 18012 21644 21364 21672
rect 18012 21632 18018 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 25958 21672 25964 21684
rect 25919 21644 25964 21672
rect 25958 21632 25964 21644
rect 26016 21632 26022 21684
rect 8772 21576 9444 21604
rect 4672 21564 4678 21576
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 3878 21536 3884 21548
rect 3099 21508 3884 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 7745 21539 7803 21545
rect 7745 21536 7757 21539
rect 4908 21508 7757 21536
rect 4908 21480 4936 21508
rect 7745 21505 7757 21508
rect 7791 21505 7803 21539
rect 8018 21536 8024 21548
rect 7979 21508 8024 21536
rect 7745 21499 7803 21505
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 4890 21468 4896 21480
rect 2823 21440 4896 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 4632 21344 4660 21440
rect 4890 21428 4896 21440
rect 4948 21428 4954 21480
rect 5626 21468 5632 21480
rect 5587 21440 5632 21468
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 7760 21468 7788 21499
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 12710 21536 12716 21548
rect 12671 21508 12716 21536
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 24673 21539 24731 21545
rect 24673 21505 24685 21539
rect 24719 21536 24731 21539
rect 24854 21536 24860 21548
rect 24719 21508 24860 21536
rect 24719 21505 24731 21508
rect 24673 21499 24731 21505
rect 24854 21496 24860 21508
rect 24912 21496 24918 21548
rect 9493 21471 9551 21477
rect 9493 21468 9505 21471
rect 7760 21440 9505 21468
rect 9493 21437 9505 21440
rect 9539 21468 9551 21471
rect 11146 21468 11152 21480
rect 9539 21440 11152 21468
rect 9539 21437 9551 21440
rect 9493 21431 9551 21437
rect 11146 21428 11152 21440
rect 11204 21468 11210 21480
rect 12161 21471 12219 21477
rect 12161 21468 12173 21471
rect 11204 21440 12173 21468
rect 11204 21428 11210 21440
rect 12161 21437 12173 21440
rect 12207 21468 12219 21471
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 12207 21440 12449 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 15657 21471 15715 21477
rect 15657 21437 15669 21471
rect 15703 21468 15715 21471
rect 21726 21468 21732 21480
rect 15703 21440 21732 21468
rect 15703 21437 15715 21440
rect 15657 21431 15715 21437
rect 21726 21428 21732 21440
rect 21784 21428 21790 21480
rect 24397 21471 24455 21477
rect 24397 21468 24409 21471
rect 24228 21440 24409 21468
rect 14090 21400 14096 21412
rect 14051 21372 14096 21400
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 24228 21344 24256 21440
rect 24397 21437 24409 21440
rect 24443 21437 24455 21471
rect 24397 21431 24455 21437
rect 4614 21332 4620 21344
rect 4575 21304 4620 21332
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 10502 21292 10508 21344
rect 10560 21332 10566 21344
rect 15194 21332 15200 21344
rect 10560 21304 15200 21332
rect 10560 21292 10566 21304
rect 15194 21292 15200 21304
rect 15252 21292 15258 21344
rect 15746 21332 15752 21344
rect 15707 21304 15752 21332
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 24210 21332 24216 21344
rect 24171 21304 24216 21332
rect 24210 21292 24216 21304
rect 24268 21292 24274 21344
rect 1104 21242 29256 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 29256 21242
rect 1104 21168 29256 21190
rect 3786 21088 3792 21140
rect 3844 21128 3850 21140
rect 7466 21128 7472 21140
rect 3844 21100 7472 21128
rect 3844 21088 3850 21100
rect 7466 21088 7472 21100
rect 7524 21088 7530 21140
rect 7558 21088 7564 21140
rect 7616 21128 7622 21140
rect 18230 21128 18236 21140
rect 7616 21100 18236 21128
rect 7616 21088 7622 21100
rect 18230 21088 18236 21100
rect 18288 21088 18294 21140
rect 23658 21060 23664 21072
rect 23619 21032 23664 21060
rect 23658 21020 23664 21032
rect 23716 21020 23722 21072
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20893 22063 20927
rect 22278 20924 22284 20936
rect 22239 20896 22284 20924
rect 22005 20887 22063 20893
rect 11054 20816 11060 20868
rect 11112 20856 11118 20868
rect 16206 20856 16212 20868
rect 11112 20828 16212 20856
rect 11112 20816 11118 20828
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 22020 20788 22048 20887
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 23845 20791 23903 20797
rect 23845 20788 23857 20791
rect 22020 20760 23857 20788
rect 23845 20757 23857 20760
rect 23891 20788 23903 20791
rect 24210 20788 24216 20800
rect 23891 20760 24216 20788
rect 23891 20757 23903 20760
rect 23845 20751 23903 20757
rect 24210 20748 24216 20760
rect 24268 20788 24274 20800
rect 24762 20788 24768 20800
rect 24268 20760 24768 20788
rect 24268 20748 24274 20760
rect 24762 20748 24768 20760
rect 24820 20748 24826 20800
rect 26418 20748 26424 20800
rect 26476 20788 26482 20800
rect 28994 20788 29000 20800
rect 26476 20760 29000 20788
rect 26476 20748 26482 20760
rect 28994 20748 29000 20760
rect 29052 20748 29058 20800
rect 59354 20748 59360 20800
rect 59412 20788 59418 20800
rect 59906 20788 59912 20800
rect 59412 20760 59912 20788
rect 59412 20748 59418 20760
rect 59906 20748 59912 20760
rect 59964 20748 59970 20800
rect 1104 20698 29256 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 29256 20698
rect 1104 20624 29256 20646
rect 4433 20587 4491 20593
rect 4433 20553 4445 20587
rect 4479 20584 4491 20587
rect 5258 20584 5264 20596
rect 4479 20556 5264 20584
rect 4479 20553 4491 20556
rect 4433 20547 4491 20553
rect 3970 20516 3976 20528
rect 3931 20488 3976 20516
rect 3970 20476 3976 20488
rect 4028 20476 4034 20528
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 4448 20448 4476 20547
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 16301 20587 16359 20593
rect 16301 20584 16313 20587
rect 15252 20556 16313 20584
rect 15252 20544 15258 20556
rect 16301 20553 16313 20556
rect 16347 20553 16359 20587
rect 16574 20584 16580 20596
rect 16535 20556 16580 20584
rect 16301 20547 16359 20553
rect 14458 20476 14464 20528
rect 14516 20516 14522 20528
rect 15102 20516 15108 20528
rect 14516 20488 15108 20516
rect 14516 20476 14522 20488
rect 15102 20476 15108 20488
rect 15160 20516 15166 20528
rect 16316 20516 16344 20547
rect 16574 20544 16580 20556
rect 16632 20544 16638 20596
rect 23842 20584 23848 20596
rect 23803 20556 23848 20584
rect 23842 20544 23848 20556
rect 23900 20544 23906 20596
rect 17862 20516 17868 20528
rect 15160 20488 15884 20516
rect 16316 20488 17868 20516
rect 15160 20476 15166 20488
rect 14366 20448 14372 20460
rect 2915 20420 4476 20448
rect 10612 20420 14372 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 2590 20380 2596 20392
rect 2551 20352 2596 20380
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 5626 20340 5632 20392
rect 5684 20380 5690 20392
rect 10612 20389 10640 20420
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20448 14795 20451
rect 15746 20448 15752 20460
rect 14783 20420 15752 20448
rect 14783 20417 14795 20420
rect 14737 20411 14795 20417
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 5684 20352 6837 20380
rect 5684 20340 5690 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 8159 20352 10609 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 10597 20349 10609 20352
rect 10643 20349 10655 20383
rect 10597 20343 10655 20349
rect 15105 20383 15163 20389
rect 15105 20349 15117 20383
rect 15151 20349 15163 20383
rect 15105 20343 15163 20349
rect 6840 20312 6868 20343
rect 15120 20312 15148 20343
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15289 20383 15347 20389
rect 15289 20380 15301 20383
rect 15252 20352 15301 20380
rect 15252 20340 15258 20352
rect 15289 20349 15301 20352
rect 15335 20349 15347 20383
rect 15562 20380 15568 20392
rect 15523 20352 15568 20380
rect 15289 20343 15347 20349
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 15657 20383 15715 20389
rect 15657 20349 15669 20383
rect 15703 20380 15715 20383
rect 15856 20380 15884 20488
rect 17862 20476 17868 20488
rect 17920 20476 17926 20528
rect 18417 20451 18475 20457
rect 18417 20448 18429 20451
rect 18064 20420 18429 20448
rect 15703 20352 15884 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18064 20389 18092 20420
rect 18417 20417 18429 20420
rect 18463 20448 18475 20451
rect 27430 20448 27436 20460
rect 18463 20420 27436 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 18012 20352 18061 20380
rect 18012 20340 18018 20352
rect 18049 20349 18061 20352
rect 18095 20349 18107 20383
rect 18049 20343 18107 20349
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20380 22615 20383
rect 23474 20380 23480 20392
rect 22603 20352 23480 20380
rect 22603 20349 22615 20352
rect 22557 20343 22615 20349
rect 23474 20340 23480 20352
rect 23532 20340 23538 20392
rect 23658 20380 23664 20392
rect 23716 20389 23722 20392
rect 23625 20352 23664 20380
rect 23658 20340 23664 20352
rect 23716 20343 23725 20389
rect 26329 20383 26387 20389
rect 26329 20349 26341 20383
rect 26375 20380 26387 20383
rect 26418 20380 26424 20392
rect 26375 20352 26424 20380
rect 26375 20349 26387 20352
rect 26329 20343 26387 20349
rect 23716 20340 23722 20343
rect 26418 20340 26424 20352
rect 26476 20340 26482 20392
rect 16574 20312 16580 20324
rect 6840 20284 8340 20312
rect 15120 20284 16580 20312
rect 4614 20244 4620 20256
rect 4575 20216 4620 20244
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 7006 20244 7012 20256
rect 6052 20216 7012 20244
rect 6052 20204 6058 20216
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 8312 20253 8340 20284
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 16758 20272 16764 20324
rect 16816 20312 16822 20324
rect 16816 20284 23520 20312
rect 16816 20272 16822 20284
rect 8297 20247 8355 20253
rect 8297 20213 8309 20247
rect 8343 20213 8355 20247
rect 8297 20207 8355 20213
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 10781 20247 10839 20253
rect 10781 20244 10793 20247
rect 8444 20216 10793 20244
rect 8444 20204 8450 20216
rect 10781 20213 10793 20216
rect 10827 20244 10839 20247
rect 11422 20244 11428 20256
rect 10827 20216 11428 20244
rect 10827 20213 10839 20216
rect 10781 20207 10839 20213
rect 11422 20204 11428 20216
rect 11480 20204 11486 20256
rect 14642 20244 14648 20256
rect 14555 20216 14648 20244
rect 14642 20204 14648 20216
rect 14700 20244 14706 20256
rect 15562 20244 15568 20256
rect 14700 20216 15568 20244
rect 14700 20204 14706 20216
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16114 20244 16120 20256
rect 16075 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 18138 20244 18144 20256
rect 18099 20216 18144 20244
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 22649 20247 22707 20253
rect 22649 20244 22661 20247
rect 22428 20216 22661 20244
rect 22428 20204 22434 20216
rect 22649 20213 22661 20216
rect 22695 20213 22707 20247
rect 23492 20244 23520 20284
rect 23658 20244 23664 20256
rect 23492 20216 23664 20244
rect 22649 20207 22707 20213
rect 23658 20204 23664 20216
rect 23716 20244 23722 20256
rect 24029 20247 24087 20253
rect 24029 20244 24041 20247
rect 23716 20216 24041 20244
rect 23716 20204 23722 20216
rect 24029 20213 24041 20216
rect 24075 20213 24087 20247
rect 24029 20207 24087 20213
rect 26421 20247 26479 20253
rect 26421 20213 26433 20247
rect 26467 20244 26479 20247
rect 27154 20244 27160 20256
rect 26467 20216 27160 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 27154 20204 27160 20216
rect 27212 20204 27218 20256
rect 1104 20154 29256 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 29256 20154
rect 1104 20080 29256 20102
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 16114 20040 16120 20052
rect 9180 20012 16120 20040
rect 9180 20000 9186 20012
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 17954 20040 17960 20052
rect 17915 20012 17960 20040
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 20438 20040 20444 20052
rect 20399 20012 20444 20040
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20040 21422 20052
rect 21416 20012 21496 20040
rect 21416 20000 21422 20012
rect 8294 19972 8300 19984
rect 5368 19944 8300 19972
rect 5368 19913 5396 19944
rect 8294 19932 8300 19944
rect 8352 19932 8358 19984
rect 5353 19907 5411 19913
rect 5353 19873 5365 19907
rect 5399 19873 5411 19907
rect 5353 19867 5411 19873
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19904 5963 19907
rect 5994 19904 6000 19916
rect 5951 19876 6000 19904
rect 5951 19873 5963 19876
rect 5905 19867 5963 19873
rect 5994 19864 6000 19876
rect 6052 19864 6058 19916
rect 6089 19907 6147 19913
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6914 19904 6920 19916
rect 6135 19876 6920 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 11422 19904 11428 19916
rect 11383 19876 11428 19904
rect 11422 19864 11428 19876
rect 11480 19904 11486 19916
rect 11977 19907 12035 19913
rect 11977 19904 11989 19907
rect 11480 19876 11989 19904
rect 11480 19864 11486 19876
rect 11977 19873 11989 19876
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 12161 19907 12219 19913
rect 12161 19873 12173 19907
rect 12207 19904 12219 19907
rect 12986 19904 12992 19916
rect 12207 19876 12992 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 20349 19907 20407 19913
rect 20349 19873 20361 19907
rect 20395 19904 20407 19907
rect 20456 19904 20484 20000
rect 21468 19913 21496 20012
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 22649 20043 22707 20049
rect 22649 20040 22661 20043
rect 22336 20012 22661 20040
rect 22336 20000 22342 20012
rect 22649 20009 22661 20012
rect 22695 20009 22707 20043
rect 22649 20003 22707 20009
rect 20395 19876 20484 19904
rect 21453 19907 21511 19913
rect 20395 19873 20407 19876
rect 20349 19867 20407 19873
rect 21453 19873 21465 19907
rect 21499 19873 21511 19907
rect 21453 19867 21511 19873
rect 21637 19907 21695 19913
rect 21637 19873 21649 19907
rect 21683 19904 21695 19907
rect 22002 19904 22008 19916
rect 21683 19876 22008 19904
rect 21683 19873 21695 19876
rect 21637 19867 21695 19873
rect 22002 19864 22008 19876
rect 22060 19904 22066 19916
rect 22189 19907 22247 19913
rect 22189 19904 22201 19907
rect 22060 19876 22201 19904
rect 22060 19864 22066 19876
rect 22189 19873 22201 19876
rect 22235 19873 22247 19907
rect 22370 19904 22376 19916
rect 22331 19876 22376 19904
rect 22189 19867 22247 19873
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 23842 19864 23848 19916
rect 23900 19904 23906 19916
rect 24857 19907 24915 19913
rect 24857 19904 24869 19907
rect 23900 19876 24869 19904
rect 23900 19864 23906 19876
rect 24857 19873 24869 19876
rect 24903 19873 24915 19907
rect 24857 19867 24915 19873
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 26513 19907 26571 19913
rect 26513 19904 26525 19907
rect 26292 19876 26525 19904
rect 26292 19864 26298 19876
rect 26513 19873 26525 19876
rect 26559 19904 26571 19907
rect 28994 19904 29000 19916
rect 26559 19876 29000 19904
rect 26559 19873 26571 19876
rect 26513 19867 26571 19873
rect 28994 19864 29000 19876
rect 29052 19864 29058 19916
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 5000 19808 5181 19836
rect 5000 19712 5028 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19805 11299 19839
rect 11241 19799 11299 19805
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19805 16635 19839
rect 16850 19836 16856 19848
rect 16811 19808 16856 19836
rect 16577 19799 16635 19805
rect 6270 19768 6276 19780
rect 6231 19740 6276 19768
rect 6270 19728 6276 19740
rect 6328 19728 6334 19780
rect 11256 19712 11284 19799
rect 12158 19728 12164 19780
rect 12216 19768 12222 19780
rect 16393 19771 16451 19777
rect 16393 19768 16405 19771
rect 12216 19740 16405 19768
rect 12216 19728 12222 19740
rect 16393 19737 16405 19740
rect 16439 19768 16451 19771
rect 16592 19768 16620 19799
rect 16850 19796 16856 19808
rect 16908 19796 16914 19848
rect 16439 19740 16620 19768
rect 16439 19737 16451 19740
rect 16393 19731 16451 19737
rect 4982 19700 4988 19712
rect 4943 19672 4988 19700
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 11149 19703 11207 19709
rect 11149 19669 11161 19703
rect 11195 19700 11207 19703
rect 11238 19700 11244 19712
rect 11195 19672 11244 19700
rect 11195 19669 11207 19672
rect 11149 19663 11207 19669
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 20162 19700 20168 19712
rect 12492 19672 12537 19700
rect 20123 19672 20168 19700
rect 12492 19660 12498 19672
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 24946 19660 24952 19712
rect 25004 19700 25010 19712
rect 25041 19703 25099 19709
rect 25041 19700 25053 19703
rect 25004 19672 25053 19700
rect 25004 19660 25010 19672
rect 25041 19669 25053 19672
rect 25087 19669 25099 19703
rect 26602 19700 26608 19712
rect 26563 19672 26608 19700
rect 25041 19663 25099 19669
rect 26602 19660 26608 19672
rect 26660 19660 26666 19712
rect 1104 19610 29256 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 29256 19610
rect 86678 19592 86684 19644
rect 86736 19632 86742 19644
rect 87230 19632 87236 19644
rect 86736 19604 87236 19632
rect 86736 19592 86742 19604
rect 87230 19592 87236 19604
rect 87288 19592 87294 19644
rect 1104 19536 29256 19558
rect 4982 19456 4988 19508
rect 5040 19496 5046 19508
rect 24854 19496 24860 19508
rect 5040 19468 24860 19496
rect 5040 19456 5046 19468
rect 24854 19456 24860 19468
rect 24912 19496 24918 19508
rect 24912 19468 25176 19496
rect 24912 19456 24918 19468
rect 12986 19428 12992 19440
rect 12947 19400 12992 19428
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 9950 19360 9956 19372
rect 9447 19332 9956 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 25148 19360 25176 19468
rect 26510 19456 26516 19508
rect 26568 19496 26574 19508
rect 26973 19499 27031 19505
rect 26973 19496 26985 19499
rect 26568 19468 26985 19496
rect 26568 19456 26574 19468
rect 26973 19465 26985 19468
rect 27019 19465 27031 19499
rect 26973 19459 27031 19465
rect 26510 19360 26516 19372
rect 25148 19332 26516 19360
rect 26510 19320 26516 19332
rect 26568 19320 26574 19372
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 6840 19224 6868 19255
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 6972 19264 7017 19292
rect 7944 19264 8125 19292
rect 6972 19252 6978 19264
rect 6840 19196 7236 19224
rect 7208 19168 7236 19196
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 7944 19165 7972 19264
rect 8113 19261 8125 19264
rect 8159 19261 8171 19295
rect 8294 19292 8300 19304
rect 8255 19264 8300 19292
rect 8113 19255 8171 19261
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19261 8907 19295
rect 8849 19255 8907 19261
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 10321 19295 10379 19301
rect 10321 19261 10333 19295
rect 10367 19292 10379 19295
rect 10686 19292 10692 19304
rect 10367 19264 10692 19292
rect 10367 19261 10379 19264
rect 10321 19255 10379 19261
rect 8312 19224 8340 19252
rect 8864 19224 8892 19255
rect 8312 19196 8892 19224
rect 9048 19224 9076 19255
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12851 19264 12909 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 16758 19292 16764 19304
rect 16719 19264 16764 19292
rect 12897 19255 12955 19261
rect 16758 19252 16764 19264
rect 16816 19292 16822 19304
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 16816 19264 16865 19292
rect 16816 19252 16822 19264
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 24854 19252 24860 19304
rect 24912 19292 24918 19304
rect 25409 19295 25467 19301
rect 25409 19292 25421 19295
rect 24912 19264 25421 19292
rect 24912 19252 24918 19264
rect 25409 19261 25421 19264
rect 25455 19292 25467 19295
rect 25593 19295 25651 19301
rect 25593 19292 25605 19295
rect 25455 19264 25605 19292
rect 25455 19261 25467 19264
rect 25409 19255 25467 19261
rect 25593 19261 25605 19264
rect 25639 19261 25651 19295
rect 25593 19255 25651 19261
rect 25869 19295 25927 19301
rect 25869 19261 25881 19295
rect 25915 19292 25927 19295
rect 27706 19292 27712 19304
rect 25915 19264 27712 19292
rect 25915 19261 25927 19264
rect 25869 19255 25927 19261
rect 27706 19252 27712 19264
rect 27764 19252 27770 19304
rect 10413 19227 10471 19233
rect 10413 19224 10425 19227
rect 9048 19196 10425 19224
rect 10413 19193 10425 19196
rect 10459 19193 10471 19227
rect 17678 19224 17684 19236
rect 10413 19187 10471 19193
rect 10520 19196 17684 19224
rect 7929 19159 7987 19165
rect 7929 19156 7941 19159
rect 7892 19128 7941 19156
rect 7892 19116 7898 19128
rect 7929 19125 7941 19128
rect 7975 19156 7987 19159
rect 10520 19156 10548 19196
rect 17678 19184 17684 19196
rect 17736 19224 17742 19236
rect 25682 19224 25688 19236
rect 17736 19196 25688 19224
rect 17736 19184 17742 19196
rect 25682 19184 25688 19196
rect 25740 19184 25746 19236
rect 10686 19156 10692 19168
rect 7975 19128 10548 19156
rect 10647 19128 10692 19156
rect 7975 19125 7987 19128
rect 7929 19119 7987 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 12805 19159 12863 19165
rect 12805 19125 12817 19159
rect 12851 19156 12863 19159
rect 13265 19159 13323 19165
rect 13265 19156 13277 19159
rect 12851 19128 13277 19156
rect 12851 19125 12863 19128
rect 12805 19119 12863 19125
rect 13265 19125 13277 19128
rect 13311 19156 13323 19159
rect 13722 19156 13728 19168
rect 13311 19128 13728 19156
rect 13311 19125 13323 19128
rect 13265 19119 13323 19125
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 17034 19156 17040 19168
rect 16947 19128 17040 19156
rect 17034 19116 17040 19128
rect 17092 19156 17098 19168
rect 22002 19156 22008 19168
rect 17092 19128 22008 19156
rect 17092 19116 17098 19128
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 23566 19116 23572 19168
rect 23624 19156 23630 19168
rect 27246 19156 27252 19168
rect 23624 19128 27252 19156
rect 23624 19116 23630 19128
rect 27246 19116 27252 19128
rect 27304 19116 27310 19168
rect 1104 19066 29256 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 29256 19066
rect 1104 18992 29256 19014
rect 6273 18955 6331 18961
rect 6273 18921 6285 18955
rect 6319 18952 6331 18955
rect 7190 18952 7196 18964
rect 6319 18924 7196 18952
rect 6319 18921 6331 18924
rect 6273 18915 6331 18921
rect 7190 18912 7196 18924
rect 7248 18952 7254 18964
rect 14642 18952 14648 18964
rect 7248 18924 14648 18952
rect 7248 18912 7254 18924
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 16206 18952 16212 18964
rect 16167 18924 16212 18952
rect 16206 18912 16212 18924
rect 16264 18952 16270 18964
rect 16264 18924 16344 18952
rect 16264 18912 16270 18924
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 6270 18816 6276 18828
rect 5031 18788 6276 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 9950 18816 9956 18828
rect 9911 18788 9956 18816
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 16316 18825 16344 18924
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 17497 18955 17555 18961
rect 17497 18952 17509 18955
rect 16908 18924 17509 18952
rect 16908 18912 16914 18924
rect 17497 18921 17509 18924
rect 17543 18921 17555 18955
rect 17497 18915 17555 18921
rect 20349 18955 20407 18961
rect 20349 18921 20361 18955
rect 20395 18952 20407 18955
rect 23566 18952 23572 18964
rect 20395 18924 23572 18952
rect 20395 18921 20407 18924
rect 20349 18915 20407 18921
rect 18966 18884 18972 18896
rect 16408 18856 18972 18884
rect 16301 18819 16359 18825
rect 12492 18788 12537 18816
rect 12492 18776 12498 18788
rect 16301 18785 16313 18819
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 4614 18708 4620 18760
rect 4672 18748 4678 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4672 18720 4721 18748
rect 4672 18708 4678 18720
rect 4709 18717 4721 18720
rect 4755 18748 4767 18751
rect 6457 18751 6515 18757
rect 6457 18748 6469 18751
rect 4755 18720 6469 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 6457 18717 6469 18720
rect 6503 18717 6515 18751
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 6457 18711 6515 18717
rect 9674 18708 9680 18720
rect 9732 18748 9738 18760
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 9732 18720 11437 18748
rect 9732 18708 9738 18720
rect 11425 18717 11437 18720
rect 11471 18748 11483 18751
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 11471 18720 11989 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 11977 18717 11989 18720
rect 12023 18748 12035 18751
rect 12158 18748 12164 18760
rect 12023 18720 12164 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 16408 18748 16436 18856
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 17034 18816 17040 18828
rect 16531 18788 17040 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 17221 18819 17279 18825
rect 17221 18785 17233 18819
rect 17267 18816 17279 18819
rect 18138 18816 18144 18828
rect 17267 18788 18144 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 19426 18816 19432 18828
rect 19387 18788 19432 18816
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 19981 18819 20039 18825
rect 19981 18785 19993 18819
rect 20027 18816 20039 18819
rect 20364 18816 20392 18915
rect 23566 18912 23572 18924
rect 23624 18912 23630 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 23937 18955 23995 18961
rect 23937 18952 23949 18955
rect 23808 18924 23949 18952
rect 23808 18912 23814 18924
rect 23937 18921 23949 18924
rect 23983 18952 23995 18955
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 23983 18924 24041 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 26237 18955 26295 18961
rect 26237 18952 26249 18955
rect 25740 18924 26249 18952
rect 25740 18912 25746 18924
rect 26237 18921 26249 18924
rect 26283 18952 26295 18955
rect 27706 18952 27712 18964
rect 26283 18924 26832 18952
rect 27667 18924 27712 18952
rect 26283 18921 26295 18924
rect 26237 18915 26295 18921
rect 22002 18844 22008 18896
rect 22060 18884 22066 18896
rect 22060 18856 26740 18884
rect 22060 18844 22066 18856
rect 20027 18788 20392 18816
rect 23937 18819 23995 18825
rect 20027 18785 20039 18788
rect 19981 18779 20039 18785
rect 23937 18785 23949 18819
rect 23983 18816 23995 18819
rect 24213 18819 24271 18825
rect 24213 18816 24225 18819
rect 23983 18788 24225 18816
rect 23983 18785 23995 18788
rect 23937 18779 23995 18785
rect 24213 18785 24225 18788
rect 24259 18785 24271 18819
rect 24213 18779 24271 18785
rect 24397 18819 24455 18825
rect 24397 18785 24409 18819
rect 24443 18816 24455 18819
rect 24946 18816 24952 18828
rect 24443 18788 24952 18816
rect 24443 18785 24455 18788
rect 24397 18779 24455 18785
rect 18782 18748 18788 18760
rect 13556 18720 16436 18748
rect 18743 18720 18788 18748
rect 10686 18572 10692 18624
rect 10744 18612 10750 18624
rect 11241 18615 11299 18621
rect 11241 18612 11253 18615
rect 10744 18584 11253 18612
rect 10744 18572 10750 18584
rect 11241 18581 11253 18584
rect 11287 18612 11299 18615
rect 13556 18612 13584 18720
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19334 18748 19340 18760
rect 19295 18720 19340 18748
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19812 18748 19840 18779
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19812 18720 20177 18748
rect 20165 18717 20177 18720
rect 20211 18748 20223 18751
rect 20254 18748 20260 18760
rect 20211 18720 20260 18748
rect 20211 18717 20223 18720
rect 20165 18711 20223 18717
rect 20254 18708 20260 18720
rect 20312 18748 20318 18760
rect 22830 18748 22836 18760
rect 20312 18720 22836 18748
rect 20312 18708 20318 18720
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 23952 18680 23980 18779
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 25133 18819 25191 18825
rect 25133 18785 25145 18819
rect 25179 18816 25191 18819
rect 26602 18816 26608 18828
rect 25179 18788 26608 18816
rect 25179 18785 25191 18788
rect 25133 18779 25191 18785
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 26712 18825 26740 18856
rect 26804 18825 26832 18924
rect 27706 18912 27712 18924
rect 27764 18912 27770 18964
rect 26697 18819 26755 18825
rect 26697 18785 26709 18819
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 26789 18819 26847 18825
rect 26789 18785 26801 18819
rect 26835 18785 26847 18819
rect 27154 18816 27160 18828
rect 27115 18788 27160 18816
rect 26789 18779 26847 18785
rect 27154 18776 27160 18788
rect 27212 18776 27218 18828
rect 27246 18776 27252 18828
rect 27304 18816 27310 18828
rect 27304 18788 27349 18816
rect 27304 18776 27310 18788
rect 17276 18652 23980 18680
rect 17276 18640 17282 18652
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25317 18683 25375 18689
rect 25317 18680 25329 18683
rect 25188 18652 25329 18680
rect 25188 18640 25194 18652
rect 25317 18649 25329 18652
rect 25363 18649 25375 18683
rect 25317 18643 25375 18649
rect 13722 18612 13728 18624
rect 11287 18584 13584 18612
rect 13635 18584 13728 18612
rect 11287 18581 11299 18584
rect 11241 18575 11299 18581
rect 13722 18572 13728 18584
rect 13780 18612 13786 18624
rect 19150 18612 19156 18624
rect 13780 18584 19156 18612
rect 13780 18572 13786 18584
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 24946 18572 24952 18624
rect 25004 18612 25010 18624
rect 27246 18612 27252 18624
rect 25004 18584 27252 18612
rect 25004 18572 25010 18584
rect 27246 18572 27252 18584
rect 27304 18572 27310 18624
rect 1104 18522 29256 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 29256 18522
rect 1104 18448 29256 18470
rect 4433 18411 4491 18417
rect 4433 18377 4445 18411
rect 4479 18408 4491 18411
rect 9214 18408 9220 18420
rect 4479 18380 9220 18408
rect 4479 18377 4491 18380
rect 4433 18371 4491 18377
rect 2590 18272 2596 18284
rect 2551 18244 2596 18272
rect 2590 18232 2596 18244
rect 2648 18232 2654 18284
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 4448 18272 4476 18371
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 17218 18408 17224 18420
rect 11296 18380 17224 18408
rect 11296 18368 11302 18380
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 20254 18408 20260 18420
rect 20215 18380 20260 18408
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 26234 18408 26240 18420
rect 26195 18380 26240 18408
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 20272 18340 20300 18368
rect 2915 18244 4476 18272
rect 19352 18312 20300 18340
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 9858 18204 9864 18216
rect 9819 18176 9864 18204
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 14185 18207 14243 18213
rect 14185 18173 14197 18207
rect 14231 18204 14243 18207
rect 18782 18204 18788 18216
rect 14231 18176 18788 18204
rect 14231 18173 14243 18176
rect 14185 18167 14243 18173
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 19352 18213 19380 18312
rect 25130 18272 25136 18284
rect 25091 18244 25136 18272
rect 25130 18232 25136 18244
rect 25188 18232 25194 18284
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 18693 18139 18751 18145
rect 18693 18136 18705 18139
rect 18012 18108 18705 18136
rect 18012 18096 18018 18108
rect 18693 18105 18705 18108
rect 18739 18105 18751 18139
rect 19168 18136 19196 18167
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 19705 18207 19763 18213
rect 19705 18204 19717 18207
rect 19484 18176 19717 18204
rect 19484 18164 19490 18176
rect 19705 18173 19717 18176
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 20990 18204 20996 18216
rect 19935 18176 20996 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 20990 18164 20996 18176
rect 21048 18164 21054 18216
rect 24854 18204 24860 18216
rect 24815 18176 24860 18204
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 26786 18204 26792 18216
rect 24964 18176 26792 18204
rect 20073 18139 20131 18145
rect 20073 18136 20085 18139
rect 19168 18108 20085 18136
rect 18693 18099 18751 18105
rect 20073 18105 20085 18108
rect 20119 18136 20131 18139
rect 24964 18136 24992 18176
rect 26786 18164 26792 18176
rect 26844 18164 26850 18216
rect 20119 18108 24992 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 4154 18068 4160 18080
rect 4115 18040 4160 18068
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4614 18068 4620 18080
rect 4575 18040 4620 18068
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14277 18071 14335 18077
rect 14277 18068 14289 18071
rect 13872 18040 14289 18068
rect 13872 18028 13878 18040
rect 14277 18037 14289 18040
rect 14323 18037 14335 18071
rect 14277 18031 14335 18037
rect 24765 18071 24823 18077
rect 24765 18037 24777 18071
rect 24811 18068 24823 18071
rect 24854 18068 24860 18080
rect 24811 18040 24860 18068
rect 24811 18037 24823 18040
rect 24765 18031 24823 18037
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 1104 17978 29256 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 29256 17978
rect 1104 17904 29256 17926
rect 20073 17867 20131 17873
rect 20073 17864 20085 17867
rect 19260 17836 20085 17864
rect 8018 17756 8024 17808
rect 8076 17796 8082 17808
rect 8202 17796 8208 17808
rect 8076 17768 8208 17796
rect 8076 17756 8082 17768
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 7837 17731 7895 17737
rect 7837 17697 7849 17731
rect 7883 17728 7895 17731
rect 14093 17731 14151 17737
rect 7883 17700 8248 17728
rect 7883 17697 7895 17700
rect 7837 17691 7895 17697
rect 8110 17620 8116 17672
rect 8168 17620 8174 17672
rect 8128 17536 8156 17620
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 7929 17527 7987 17533
rect 7929 17524 7941 17527
rect 7800 17496 7941 17524
rect 7800 17484 7806 17496
rect 7929 17493 7941 17496
rect 7975 17493 7987 17527
rect 7929 17487 7987 17493
rect 8110 17484 8116 17536
rect 8168 17484 8174 17536
rect 8220 17533 8248 17700
rect 14093 17697 14105 17731
rect 14139 17728 14151 17731
rect 17954 17728 17960 17740
rect 14139 17700 17960 17728
rect 14139 17697 14151 17700
rect 14093 17691 14151 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 18230 17688 18236 17740
rect 18288 17728 18294 17740
rect 19260 17737 19288 17836
rect 20073 17833 20085 17836
rect 20119 17864 20131 17867
rect 20162 17864 20168 17876
rect 20119 17836 20168 17864
rect 20119 17833 20131 17836
rect 20073 17827 20131 17833
rect 20162 17824 20168 17836
rect 20220 17864 20226 17876
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 20220 17836 20269 17864
rect 20220 17824 20226 17836
rect 20257 17833 20269 17836
rect 20303 17864 20315 17867
rect 23934 17864 23940 17876
rect 20303 17836 23940 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 23934 17824 23940 17836
rect 23992 17824 23998 17876
rect 19334 17756 19340 17808
rect 19392 17796 19398 17808
rect 20993 17799 21051 17805
rect 20993 17796 21005 17799
rect 19392 17768 21005 17796
rect 19392 17756 19398 17768
rect 19444 17737 19472 17768
rect 20993 17765 21005 17768
rect 21039 17765 21051 17799
rect 20993 17759 21051 17765
rect 86678 17756 86684 17808
rect 86736 17796 86742 17808
rect 87598 17796 87604 17808
rect 86736 17768 87604 17796
rect 86736 17756 86742 17768
rect 87598 17756 87604 17768
rect 87656 17756 87662 17808
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 18288 17700 18429 17728
rect 18288 17688 18294 17700
rect 18417 17697 18429 17700
rect 18463 17728 18475 17731
rect 18693 17731 18751 17737
rect 18463 17700 18644 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 18616 17672 18644 17700
rect 18693 17697 18705 17731
rect 18739 17728 18751 17731
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18739 17700 19257 17728
rect 18739 17697 18751 17700
rect 18693 17691 18751 17697
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 27985 17731 28043 17737
rect 27985 17697 27997 17731
rect 28031 17728 28043 17731
rect 28074 17728 28080 17740
rect 28031 17700 28080 17728
rect 28031 17697 28043 17700
rect 27985 17691 28043 17697
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 13412 17632 13553 17660
rect 13412 17620 13418 17632
rect 13541 17629 13553 17632
rect 13587 17660 13599 17663
rect 18598 17660 18604 17672
rect 13587 17632 18460 17660
rect 18559 17632 18604 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 13078 17552 13084 17604
rect 13136 17592 13142 17604
rect 14185 17595 14243 17601
rect 14185 17592 14197 17595
rect 13136 17564 14197 17592
rect 13136 17552 13142 17564
rect 14185 17561 14197 17564
rect 14231 17561 14243 17595
rect 14185 17555 14243 17561
rect 8205 17527 8263 17533
rect 8205 17493 8217 17527
rect 8251 17524 8263 17527
rect 8570 17524 8576 17536
rect 8251 17496 8576 17524
rect 8251 17493 8263 17496
rect 8205 17487 8263 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 18230 17524 18236 17536
rect 13596 17496 18236 17524
rect 13596 17484 13602 17496
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18432 17524 18460 17632
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19613 17595 19671 17601
rect 19613 17592 19625 17595
rect 19484 17564 19625 17592
rect 19484 17552 19490 17564
rect 19613 17561 19625 17564
rect 19659 17561 19671 17595
rect 19613 17555 19671 17561
rect 20254 17524 20260 17536
rect 18432 17496 20260 17524
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 20806 17484 20812 17536
rect 20864 17524 20870 17536
rect 20916 17524 20944 17691
rect 28074 17688 28080 17700
rect 28132 17728 28138 17740
rect 28902 17728 28908 17740
rect 28132 17700 28908 17728
rect 28132 17688 28138 17700
rect 28902 17688 28908 17700
rect 28960 17688 28966 17740
rect 21177 17527 21235 17533
rect 21177 17524 21189 17527
rect 20864 17496 21189 17524
rect 20864 17484 20870 17496
rect 21177 17493 21189 17496
rect 21223 17493 21235 17527
rect 21177 17487 21235 17493
rect 27338 17484 27344 17536
rect 27396 17524 27402 17536
rect 28077 17527 28135 17533
rect 28077 17524 28089 17527
rect 27396 17496 28089 17524
rect 27396 17484 27402 17496
rect 28077 17493 28089 17496
rect 28123 17493 28135 17527
rect 28077 17487 28135 17493
rect 1104 17434 29256 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 29256 17434
rect 86678 17416 86684 17468
rect 86736 17456 86742 17468
rect 87414 17456 87420 17468
rect 86736 17428 87420 17456
rect 86736 17416 86742 17428
rect 87414 17416 87420 17428
rect 87472 17416 87478 17468
rect 1104 17360 29256 17382
rect 59354 17348 59360 17400
rect 59412 17388 59418 17400
rect 59630 17388 59636 17400
rect 59412 17360 59636 17388
rect 59412 17348 59418 17360
rect 59630 17348 59636 17360
rect 59688 17348 59694 17400
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 9766 17320 9772 17332
rect 4479 17292 9772 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 2590 17184 2596 17196
rect 2551 17156 2596 17184
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17184 2927 17187
rect 4448 17184 4476 17283
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10778 17320 10784 17332
rect 9916 17292 10784 17320
rect 9916 17280 9922 17292
rect 10778 17280 10784 17292
rect 10836 17320 10842 17332
rect 13173 17323 13231 17329
rect 13173 17320 13185 17323
rect 10836 17292 13185 17320
rect 10836 17280 10842 17292
rect 13173 17289 13185 17292
rect 13219 17289 13231 17323
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 13173 17283 13231 17289
rect 14292 17292 15301 17320
rect 13538 17252 13544 17264
rect 2915 17156 4476 17184
rect 6840 17224 13544 17252
rect 2915 17153 2927 17156
rect 2869 17147 2927 17153
rect 6840 17125 6868 17224
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 14292 17252 14320 17292
rect 15289 17289 15301 17292
rect 15335 17320 15347 17323
rect 17310 17320 17316 17332
rect 15335 17292 17316 17320
rect 15335 17289 15347 17292
rect 15289 17283 15347 17289
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 13740 17224 14320 17252
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17184 13507 17187
rect 13630 17184 13636 17196
rect 13495 17156 13636 17184
rect 13495 17153 13507 17156
rect 13449 17147 13507 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 7006 17116 7012 17128
rect 6967 17088 7012 17116
rect 6825 17079 6883 17085
rect 3878 17008 3884 17060
rect 3936 17048 3942 17060
rect 6549 17051 6607 17057
rect 6549 17048 6561 17051
rect 3936 17020 6561 17048
rect 3936 17008 3942 17020
rect 6549 17017 6561 17020
rect 6595 17048 6607 17051
rect 6840 17048 6868 17079
rect 7006 17076 7012 17088
rect 7064 17076 7070 17128
rect 7561 17119 7619 17125
rect 7561 17085 7573 17119
rect 7607 17085 7619 17119
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7561 17079 7619 17085
rect 6595 17020 6868 17048
rect 7024 17048 7052 17076
rect 7576 17048 7604 17079
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 13354 17116 13360 17128
rect 13315 17088 13360 17116
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13740 17125 13768 17224
rect 19426 17184 19432 17196
rect 13832 17156 14228 17184
rect 19387 17156 19432 17184
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 7024 17020 7604 17048
rect 6595 17017 6607 17020
rect 6549 17011 6607 17017
rect 8570 17008 8576 17060
rect 8628 17048 8634 17060
rect 13081 17051 13139 17057
rect 13081 17048 13093 17051
rect 8628 17020 13093 17048
rect 8628 17008 8634 17020
rect 13081 17017 13093 17020
rect 13127 17048 13139 17051
rect 13832 17048 13860 17156
rect 14200 17128 14228 17156
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17184 26387 17187
rect 26421 17187 26479 17193
rect 26421 17184 26433 17187
rect 26375 17156 26433 17184
rect 26375 17153 26387 17156
rect 26329 17147 26387 17153
rect 26421 17153 26433 17156
rect 26467 17184 26479 17187
rect 26510 17184 26516 17196
rect 26467 17156 26516 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 26510 17144 26516 17156
rect 26568 17144 26574 17196
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14182 17116 14188 17128
rect 14143 17088 14188 17116
rect 14001 17079 14059 17085
rect 13127 17020 13860 17048
rect 13127 17017 13139 17020
rect 13081 17011 13139 17017
rect 4154 16980 4160 16992
rect 4115 16952 4160 16980
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 4614 16980 4620 16992
rect 4575 16952 4620 16980
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7340 16952 8033 16980
rect 7340 16940 7346 16952
rect 8021 16949 8033 16952
rect 8067 16949 8079 16983
rect 14016 16980 14044 17079
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 14366 17116 14372 17128
rect 14327 17088 14372 17116
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15194 17116 15200 17128
rect 15151 17088 15200 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15120 17048 15148 17079
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17116 19211 17119
rect 26605 17119 26663 17125
rect 19199 17088 21036 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 20806 17048 20812 17060
rect 14384 17020 15148 17048
rect 20767 17020 20812 17048
rect 14384 16980 14412 17020
rect 20806 17008 20812 17020
rect 20864 17008 20870 17060
rect 14826 16980 14832 16992
rect 14016 16952 14412 16980
rect 14787 16952 14832 16980
rect 8021 16943 8079 16949
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 21008 16989 21036 17088
rect 26605 17085 26617 17119
rect 26651 17085 26663 17119
rect 26605 17079 26663 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17085 27215 17119
rect 27338 17116 27344 17128
rect 27299 17088 27344 17116
rect 27157 17079 27215 17085
rect 26620 17048 26648 17079
rect 27172 17048 27200 17079
rect 27338 17076 27344 17088
rect 27396 17076 27402 17128
rect 27246 17048 27252 17060
rect 26620 17020 27252 17048
rect 27246 17008 27252 17020
rect 27304 17008 27310 17060
rect 20993 16983 21051 16989
rect 20993 16949 21005 16983
rect 21039 16980 21051 16983
rect 21634 16980 21640 16992
rect 21039 16952 21640 16980
rect 21039 16949 21051 16952
rect 20993 16943 21051 16949
rect 21634 16940 21640 16952
rect 21692 16940 21698 16992
rect 26786 16940 26792 16992
rect 26844 16980 26850 16992
rect 27617 16983 27675 16989
rect 27617 16980 27629 16983
rect 26844 16952 27629 16980
rect 26844 16940 26850 16952
rect 27617 16949 27629 16952
rect 27663 16949 27675 16983
rect 27617 16943 27675 16949
rect 1104 16890 29256 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 29256 16890
rect 1104 16816 29256 16838
rect 8570 16776 8576 16788
rect 8531 16748 8576 16776
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 20162 16776 20168 16788
rect 20123 16748 20168 16776
rect 20162 16736 20168 16748
rect 20220 16776 20226 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 20220 16748 20269 16776
rect 20220 16736 20226 16748
rect 20257 16745 20269 16748
rect 20303 16745 20315 16779
rect 20257 16739 20315 16745
rect 21634 16736 21640 16788
rect 21692 16776 21698 16788
rect 23661 16779 23719 16785
rect 23661 16776 23673 16779
rect 21692 16748 23673 16776
rect 21692 16736 21698 16748
rect 23661 16745 23673 16748
rect 23707 16776 23719 16779
rect 24854 16776 24860 16788
rect 23707 16748 24860 16776
rect 23707 16745 23719 16748
rect 23661 16739 23719 16745
rect 24854 16736 24860 16748
rect 24912 16776 24918 16788
rect 26237 16779 26295 16785
rect 26237 16776 26249 16779
rect 24912 16748 26249 16776
rect 24912 16736 24918 16748
rect 26237 16745 26249 16748
rect 26283 16745 26295 16779
rect 28074 16776 28080 16788
rect 28035 16748 28080 16776
rect 26237 16739 26295 16745
rect 12342 16708 12348 16720
rect 12255 16680 12348 16708
rect 12342 16668 12348 16680
rect 12400 16708 12406 16720
rect 20180 16708 20208 16736
rect 12400 16680 13492 16708
rect 12400 16668 12406 16680
rect 13464 16652 13492 16680
rect 18800 16680 20208 16708
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 4672 16612 7021 16640
rect 4672 16600 4678 16612
rect 7009 16609 7021 16612
rect 7055 16640 7067 16643
rect 7098 16640 7104 16652
rect 7055 16612 7104 16640
rect 7055 16609 7067 16612
rect 7009 16603 7067 16609
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 7282 16640 7288 16652
rect 7243 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 13078 16640 13084 16652
rect 12492 16612 12537 16640
rect 13039 16612 13084 16640
rect 12492 16600 12498 16612
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16640 13231 16643
rect 13262 16640 13268 16652
rect 13219 16612 13268 16640
rect 13219 16609 13231 16612
rect 13173 16603 13231 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13446 16640 13452 16652
rect 13407 16612 13452 16640
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 14366 16640 14372 16652
rect 13679 16612 14372 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 18322 16600 18328 16652
rect 18380 16640 18386 16652
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 18380 16612 18429 16640
rect 18380 16600 18386 16612
rect 18417 16609 18429 16612
rect 18463 16640 18475 16643
rect 18506 16640 18512 16652
rect 18463 16612 18512 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 18506 16600 18512 16612
rect 18564 16640 18570 16652
rect 18800 16649 18828 16680
rect 19352 16649 19380 16680
rect 18601 16643 18659 16649
rect 18601 16640 18613 16643
rect 18564 16612 18613 16640
rect 18564 16600 18570 16612
rect 18601 16609 18613 16612
rect 18647 16609 18659 16643
rect 18601 16603 18659 16609
rect 18785 16643 18843 16649
rect 18785 16609 18797 16643
rect 18831 16609 18843 16643
rect 18785 16603 18843 16609
rect 19337 16643 19395 16649
rect 19337 16609 19349 16643
rect 19383 16640 19395 16643
rect 19521 16643 19579 16649
rect 19383 16612 19417 16640
rect 19383 16609 19395 16612
rect 19337 16603 19395 16609
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 20990 16640 20996 16652
rect 19567 16612 20996 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 22830 16600 22836 16652
rect 22888 16640 22894 16652
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 22888 16612 23857 16640
rect 22888 16600 22894 16612
rect 23845 16609 23857 16612
rect 23891 16609 23903 16643
rect 26252 16640 26280 16739
rect 28074 16736 28080 16748
rect 28132 16736 28138 16788
rect 26513 16643 26571 16649
rect 26513 16640 26525 16643
rect 26252 16612 26525 16640
rect 23845 16603 23903 16609
rect 26513 16609 26525 16612
rect 26559 16609 26571 16643
rect 26786 16640 26792 16652
rect 26747 16612 26792 16640
rect 26513 16603 26571 16609
rect 26786 16600 26792 16612
rect 26844 16600 26850 16652
rect 7116 16572 7144 16600
rect 8757 16575 8815 16581
rect 8757 16572 8769 16575
rect 7116 16544 8769 16572
rect 8757 16541 8769 16544
rect 8803 16572 8815 16575
rect 8938 16572 8944 16584
rect 8803 16544 8944 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 8938 16532 8944 16544
rect 8996 16572 9002 16584
rect 9582 16572 9588 16584
rect 8996 16544 9588 16572
rect 8996 16532 9002 16544
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 19797 16439 19855 16445
rect 19797 16405 19809 16439
rect 19843 16436 19855 16439
rect 19886 16436 19892 16448
rect 19843 16408 19892 16436
rect 19843 16405 19855 16408
rect 19797 16399 19855 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 1104 16346 29256 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 29256 16346
rect 1104 16272 29256 16294
rect 4433 16235 4491 16241
rect 4433 16201 4445 16235
rect 4479 16232 4491 16235
rect 8662 16232 8668 16244
rect 4479 16204 8668 16232
rect 4479 16201 4491 16204
rect 4433 16195 4491 16201
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16096 2927 16099
rect 4448 16096 4476 16195
rect 8662 16192 8668 16204
rect 8720 16192 8726 16244
rect 8938 16232 8944 16244
rect 8899 16204 8944 16232
rect 8938 16192 8944 16204
rect 8996 16192 9002 16244
rect 9585 16235 9643 16241
rect 9585 16201 9597 16235
rect 9631 16232 9643 16235
rect 12342 16232 12348 16244
rect 9631 16204 12348 16232
rect 9631 16201 9643 16204
rect 9585 16195 9643 16201
rect 2915 16068 4476 16096
rect 2915 16065 2927 16068
rect 2869 16059 2927 16065
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 7156 16068 7205 16096
rect 7156 16056 7162 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 9692 16096 9720 16204
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 21542 16232 21548 16244
rect 14875 16204 21548 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 8895 16068 9720 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 2590 16028 2596 16040
rect 2503 16000 2596 16028
rect 2590 15988 2596 16000
rect 2648 16028 2654 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 2648 16000 4537 16028
rect 2648 15988 2654 16000
rect 4525 15997 4537 16000
rect 4571 16028 4583 16031
rect 4614 16028 4620 16040
rect 4571 16000 4620 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 7466 16028 7472 16040
rect 7427 16000 7472 16028
rect 7466 15988 7472 16000
rect 7524 15988 7530 16040
rect 9692 16037 9720 16068
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 14844 16096 14872 16195
rect 21542 16192 21548 16204
rect 21600 16192 21606 16244
rect 23658 16232 23664 16244
rect 23619 16204 23664 16232
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 24854 16232 24860 16244
rect 24815 16204 24860 16232
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 26510 16232 26516 16244
rect 26423 16204 26516 16232
rect 26510 16192 26516 16204
rect 26568 16232 26574 16244
rect 28902 16232 28908 16244
rect 26568 16204 28908 16232
rect 26568 16192 26574 16204
rect 28902 16192 28908 16204
rect 28960 16192 28966 16244
rect 19886 16096 19892 16108
rect 13311 16068 14872 16096
rect 19847 16068 19892 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 24872 16096 24900 16192
rect 24949 16099 25007 16105
rect 24949 16096 24961 16099
rect 24872 16068 24961 16096
rect 24949 16065 24961 16068
rect 24995 16065 25007 16099
rect 24949 16059 25007 16065
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 9677 15991 9735 15997
rect 12820 16000 13001 16028
rect 4154 15892 4160 15904
rect 4115 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 9766 15892 9772 15904
rect 9727 15864 9772 15892
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 12820 15901 12848 16000
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 19613 16031 19671 16037
rect 19613 15997 19625 16031
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12676 15864 12817 15892
rect 12676 15852 12682 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 13964 15864 14381 15892
rect 13964 15852 13970 15864
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 19628 15892 19656 15991
rect 23658 15988 23664 16040
rect 23716 16028 23722 16040
rect 23845 16031 23903 16037
rect 23845 16028 23857 16031
rect 23716 16000 23857 16028
rect 23716 15988 23722 16000
rect 23845 15997 23857 16000
rect 23891 15997 23903 16031
rect 25222 16028 25228 16040
rect 25183 16000 25228 16028
rect 23845 15991 23903 15997
rect 25222 15988 25228 16000
rect 25280 15988 25286 16040
rect 21266 15960 21272 15972
rect 21227 15932 21272 15960
rect 21266 15920 21272 15932
rect 21324 15920 21330 15972
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 19628 15864 21465 15892
rect 14369 15855 14427 15861
rect 21453 15861 21465 15864
rect 21499 15892 21511 15895
rect 21634 15892 21640 15904
rect 21499 15864 21640 15892
rect 21499 15861 21511 15864
rect 21453 15855 21511 15861
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 24029 15895 24087 15901
rect 24029 15861 24041 15895
rect 24075 15892 24087 15895
rect 24394 15892 24400 15904
rect 24075 15864 24400 15892
rect 24075 15861 24087 15864
rect 24029 15855 24087 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 1104 15802 29256 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 29256 15802
rect 1104 15728 29256 15750
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 7653 15691 7711 15697
rect 7653 15688 7665 15691
rect 7524 15660 7665 15688
rect 7524 15648 7530 15660
rect 7653 15657 7665 15660
rect 7699 15657 7711 15691
rect 20990 15688 20996 15700
rect 20951 15660 20996 15688
rect 7653 15651 7711 15657
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 21266 15688 21272 15700
rect 21227 15660 21272 15688
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 25222 15648 25228 15700
rect 25280 15688 25286 15700
rect 25409 15691 25467 15697
rect 25409 15688 25421 15691
rect 25280 15660 25421 15688
rect 25280 15648 25286 15660
rect 25409 15657 25421 15660
rect 25455 15657 25467 15691
rect 25409 15651 25467 15657
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 7006 15552 7012 15564
rect 6687 15524 7012 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 7006 15512 7012 15524
rect 7064 15552 7070 15564
rect 7193 15555 7251 15561
rect 7193 15552 7205 15555
rect 7064 15524 7205 15552
rect 7064 15512 7070 15524
rect 7193 15521 7205 15524
rect 7239 15521 7251 15555
rect 7193 15515 7251 15521
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15552 7435 15555
rect 9766 15552 9772 15564
rect 7423 15524 9772 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15552 20959 15555
rect 21284 15552 21312 15648
rect 26605 15623 26663 15629
rect 26605 15620 26617 15623
rect 25148 15592 26617 15620
rect 24394 15552 24400 15564
rect 20947 15524 21312 15552
rect 24355 15524 24400 15552
rect 20947 15521 20959 15524
rect 20901 15515 20959 15521
rect 24394 15512 24400 15524
rect 24452 15552 24458 15564
rect 24946 15552 24952 15564
rect 24452 15524 24952 15552
rect 24452 15512 24458 15524
rect 24946 15512 24952 15524
rect 25004 15512 25010 15564
rect 25148 15561 25176 15592
rect 26605 15589 26617 15592
rect 26651 15589 26663 15623
rect 26605 15583 26663 15589
rect 25133 15555 25191 15561
rect 25133 15521 25145 15555
rect 25179 15521 25191 15555
rect 26510 15552 26516 15564
rect 26471 15524 26516 15552
rect 25133 15515 25191 15521
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 6362 15416 6368 15428
rect 6275 15388 6368 15416
rect 6362 15376 6368 15388
rect 6420 15416 6426 15428
rect 6564 15416 6592 15447
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 24029 15487 24087 15493
rect 24029 15484 24041 15487
rect 18656 15456 24041 15484
rect 18656 15444 18662 15456
rect 24029 15453 24041 15456
rect 24075 15484 24087 15487
rect 24213 15487 24271 15493
rect 24213 15484 24225 15487
rect 24075 15456 24225 15484
rect 24075 15453 24087 15456
rect 24029 15447 24087 15453
rect 24213 15453 24225 15456
rect 24259 15453 24271 15487
rect 24213 15447 24271 15453
rect 18322 15416 18328 15428
rect 6420 15388 18328 15416
rect 6420 15376 6426 15388
rect 18322 15376 18328 15388
rect 18380 15416 18386 15428
rect 25406 15416 25412 15428
rect 18380 15388 25412 15416
rect 18380 15376 18386 15388
rect 25406 15376 25412 15388
rect 25464 15376 25470 15428
rect 1104 15258 29256 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 29256 15258
rect 1104 15184 29256 15206
rect 4525 15147 4583 15153
rect 4525 15113 4537 15147
rect 4571 15144 4583 15147
rect 10410 15144 10416 15156
rect 4571 15116 10416 15144
rect 4571 15113 4583 15116
rect 4525 15107 4583 15113
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 4540 15008 4568 15107
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 3007 14980 4568 15008
rect 13817 15011 13875 15017
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 13817 14977 13829 15011
rect 13863 15008 13875 15011
rect 13906 15008 13912 15020
rect 13863 14980 13912 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 2648 14912 2697 14940
rect 2648 14900 2654 14912
rect 2685 14909 2697 14912
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 6362 14940 6368 14952
rect 4028 14912 6368 14940
rect 4028 14900 4034 14912
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13372 14912 13553 14940
rect 4062 14804 4068 14816
rect 4023 14776 4068 14804
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13372 14813 13400 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 12676 14776 13369 14804
rect 12676 14764 12682 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 13357 14767 13415 14773
rect 15010 14764 15016 14816
rect 15068 14804 15074 14816
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 15068 14776 15117 14804
rect 15068 14764 15074 14776
rect 15105 14773 15117 14776
rect 15151 14773 15163 14807
rect 15105 14767 15163 14773
rect 1104 14714 29256 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 29256 14714
rect 1104 14640 29256 14662
rect 21542 14560 21548 14612
rect 21600 14600 21606 14612
rect 21729 14603 21787 14609
rect 21729 14600 21741 14603
rect 21600 14572 21741 14600
rect 21600 14560 21606 14572
rect 21729 14569 21741 14572
rect 21775 14569 21787 14603
rect 21729 14563 21787 14569
rect 14369 14535 14427 14541
rect 14369 14501 14381 14535
rect 14415 14532 14427 14535
rect 14734 14532 14740 14544
rect 14415 14504 14740 14532
rect 14415 14501 14427 14504
rect 14369 14495 14427 14501
rect 14734 14492 14740 14504
rect 14792 14492 14798 14544
rect 18046 14532 18052 14544
rect 18007 14504 18052 14532
rect 18046 14492 18052 14504
rect 18104 14492 18110 14544
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14464 8355 14467
rect 12434 14464 12440 14476
rect 8343 14436 12440 14464
rect 8343 14433 8355 14436
rect 8297 14427 8355 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 16393 14467 16451 14473
rect 16393 14433 16405 14467
rect 16439 14464 16451 14467
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 16439 14436 18153 14464
rect 16439 14433 16451 14436
rect 16393 14427 16451 14433
rect 18141 14433 18153 14436
rect 18187 14464 18199 14467
rect 20622 14464 20628 14476
rect 18187 14436 20628 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21560 14464 21588 14560
rect 20947 14436 21588 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 12713 14399 12771 14405
rect 12713 14396 12725 14399
rect 12636 14368 12725 14396
rect 8386 14288 8392 14340
rect 8444 14328 8450 14340
rect 9030 14328 9036 14340
rect 8444 14300 9036 14328
rect 8444 14288 8450 14300
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 12636 14272 12664 14368
rect 12713 14365 12725 14368
rect 12759 14365 12771 14399
rect 12986 14396 12992 14408
rect 12947 14368 12992 14396
rect 12713 14359 12771 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 16666 14396 16672 14408
rect 16627 14368 16672 14396
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 8481 14263 8539 14269
rect 8481 14260 8493 14263
rect 4948 14232 8493 14260
rect 4948 14220 4954 14232
rect 8481 14229 8493 14232
rect 8527 14229 8539 14263
rect 12618 14260 12624 14272
rect 12579 14232 12624 14260
rect 8481 14223 8539 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 20990 14220 20996 14272
rect 21048 14260 21054 14272
rect 21545 14263 21603 14269
rect 21545 14260 21557 14263
rect 21048 14232 21557 14260
rect 21048 14220 21054 14232
rect 21545 14229 21557 14232
rect 21591 14229 21603 14263
rect 21545 14223 21603 14229
rect 1104 14170 29256 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 29256 14170
rect 1104 14096 29256 14118
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 6178 14016 6184 14068
rect 6236 14056 6242 14068
rect 6822 14056 6828 14068
rect 6236 14028 6828 14056
rect 6236 14016 6242 14028
rect 6822 14016 6828 14028
rect 6880 14056 6886 14068
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6880 14028 7205 14056
rect 6880 14016 6886 14028
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 8941 14059 8999 14065
rect 8941 14025 8953 14059
rect 8987 14025 8999 14059
rect 8941 14019 8999 14025
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 12618 14056 12624 14068
rect 10643 14028 12624 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 8956 13988 8984 14019
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20717 14059 20775 14065
rect 20717 14056 20729 14059
rect 20680 14028 20729 14056
rect 20680 14016 20686 14028
rect 20717 14025 20729 14028
rect 20763 14025 20775 14059
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 20717 14019 20775 14025
rect 15194 13988 15200 14000
rect 3752 13960 8984 13988
rect 12728 13960 15200 13988
rect 3752 13948 3758 13960
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13920 2927 13923
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 2915 13892 4445 13920
rect 2915 13889 2927 13892
rect 2869 13883 2927 13889
rect 4433 13889 4445 13892
rect 4479 13920 4491 13923
rect 8386 13920 8392 13932
rect 4479 13892 8392 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 10594 13920 10600 13932
rect 8588 13892 10600 13920
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 6880 13824 7389 13852
rect 6880 13812 6886 13824
rect 7377 13821 7389 13824
rect 7423 13852 7435 13855
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 7423 13824 8309 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 8297 13821 8309 13824
rect 8343 13852 8355 13855
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8343 13824 8493 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 8588 13784 8616 13892
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 12728 13929 12756 13960
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 12713 13923 12771 13929
rect 12713 13920 12725 13923
rect 12452 13892 12725 13920
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13852 8818 13864
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 8812 13824 9321 13852
rect 8812 13812 8818 13824
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 10778 13852 10784 13864
rect 10739 13824 10784 13852
rect 9309 13815 9367 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 12452 13861 12480 13892
rect 12713 13889 12725 13892
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13044 13892 14013 13920
rect 13044 13880 13050 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13920 14611 13923
rect 20732 13920 20760 14019
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 14599 13892 15424 13920
rect 20732 13892 20913 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 14645 13855 14703 13861
rect 12584 13824 12629 13852
rect 12584 13812 12590 13824
rect 14645 13821 14657 13855
rect 14691 13852 14703 13855
rect 14734 13852 14740 13864
rect 14691 13824 14740 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15010 13852 15016 13864
rect 14971 13824 15016 13852
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15194 13852 15200 13864
rect 15155 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 8665 13787 8723 13793
rect 8665 13784 8677 13787
rect 8588 13756 8677 13784
rect 8665 13753 8677 13756
rect 8711 13753 8723 13787
rect 8665 13747 8723 13753
rect 3970 13716 3976 13728
rect 3931 13688 3976 13716
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 7561 13719 7619 13725
rect 7561 13685 7573 13719
rect 7607 13716 7619 13719
rect 8202 13716 8208 13728
rect 7607 13688 8208 13716
rect 7607 13685 7619 13688
rect 7561 13679 7619 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 15396 13725 15424 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 25424 13920 25452 14016
rect 25593 13923 25651 13929
rect 25593 13920 25605 13923
rect 25424 13892 25605 13920
rect 20901 13883 20959 13889
rect 25593 13889 25605 13892
rect 25639 13889 25651 13923
rect 27893 13923 27951 13929
rect 27893 13920 27905 13923
rect 25593 13883 25651 13889
rect 27080 13892 27905 13920
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 21048 13824 21189 13852
rect 21048 13812 21054 13824
rect 21177 13821 21189 13824
rect 21223 13821 21235 13855
rect 21177 13815 21235 13821
rect 24946 13812 24952 13864
rect 25004 13852 25010 13864
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25004 13824 25789 13852
rect 25004 13812 25010 13824
rect 25777 13821 25789 13824
rect 25823 13852 25835 13855
rect 26329 13855 26387 13861
rect 26329 13852 26341 13855
rect 25823 13824 26341 13852
rect 25823 13821 25835 13824
rect 25777 13815 25835 13821
rect 26329 13821 26341 13824
rect 26375 13821 26387 13855
rect 26329 13815 26387 13821
rect 26513 13855 26571 13861
rect 26513 13821 26525 13855
rect 26559 13852 26571 13855
rect 27080 13852 27108 13892
rect 27893 13889 27905 13892
rect 27939 13889 27951 13923
rect 27893 13883 27951 13889
rect 27798 13852 27804 13864
rect 26559 13824 27108 13852
rect 27759 13824 27804 13852
rect 26559 13821 26571 13824
rect 26513 13815 26571 13821
rect 27798 13812 27804 13824
rect 27856 13812 27862 13864
rect 15381 13719 15439 13725
rect 15381 13685 15393 13719
rect 15427 13716 15439 13719
rect 15746 13716 15752 13728
rect 15427 13688 15752 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 22278 13716 22284 13728
rect 22239 13688 22284 13716
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 26786 13716 26792 13728
rect 26747 13688 26792 13716
rect 26786 13676 26792 13688
rect 26844 13676 26850 13728
rect 1104 13626 29256 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 29256 13626
rect 1104 13552 29256 13574
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6236 13484 6469 13512
rect 6236 13472 6242 13484
rect 6457 13481 6469 13484
rect 6503 13481 6515 13515
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 6457 13475 6515 13481
rect 6472 13376 6500 13475
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 10502 13512 10508 13524
rect 10463 13484 10508 13512
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 18046 13472 18052 13524
rect 18104 13472 18110 13524
rect 21634 13472 21640 13524
rect 21692 13512 21698 13524
rect 23477 13515 23535 13521
rect 23477 13512 23489 13515
rect 21692 13484 23489 13512
rect 21692 13472 21698 13484
rect 23477 13481 23489 13484
rect 23523 13512 23535 13515
rect 24302 13512 24308 13524
rect 23523 13484 24308 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 24302 13472 24308 13484
rect 24360 13512 24366 13524
rect 26237 13515 26295 13521
rect 26237 13512 26249 13515
rect 24360 13484 26249 13512
rect 24360 13472 24366 13484
rect 26237 13481 26249 13484
rect 26283 13481 26295 13515
rect 26237 13475 26295 13481
rect 6825 13447 6883 13453
rect 6825 13413 6837 13447
rect 6871 13444 6883 13447
rect 7282 13444 7288 13456
rect 6871 13416 7288 13444
rect 6871 13413 6883 13416
rect 6825 13407 6883 13413
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 6641 13379 6699 13385
rect 6641 13376 6653 13379
rect 6472 13348 6653 13376
rect 6641 13345 6653 13348
rect 6687 13345 6699 13379
rect 6641 13339 6699 13345
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7576 13376 7604 13472
rect 6963 13348 7604 13376
rect 8297 13379 8355 13385
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 8478 13376 8484 13388
rect 8343 13348 8484 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 8478 13336 8484 13348
rect 8536 13376 8542 13388
rect 8849 13379 8907 13385
rect 8849 13376 8861 13379
rect 8536 13348 8861 13376
rect 8536 13336 8542 13348
rect 8849 13345 8861 13348
rect 8895 13345 8907 13379
rect 8849 13339 8907 13345
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 10520 13376 10548 13472
rect 16666 13404 16672 13456
rect 16724 13444 16730 13456
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 16724 13416 17049 13444
rect 16724 13404 16730 13416
rect 17037 13413 17049 13416
rect 17083 13413 17095 13447
rect 18064 13444 18092 13472
rect 17037 13407 17095 13413
rect 17696 13416 18092 13444
rect 17696 13385 17724 13416
rect 9907 13348 10548 13376
rect 17681 13379 17739 13385
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 17681 13345 17693 13379
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 21913 13379 21971 13385
rect 18095 13348 21772 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 8202 13308 8208 13320
rect 8163 13280 8208 13308
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17954 13308 17960 13320
rect 17915 13280 17960 13308
rect 17773 13271 17831 13277
rect 7098 13172 7104 13184
rect 7059 13144 7104 13172
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10045 13175 10103 13181
rect 10045 13172 10057 13175
rect 10008 13144 10057 13172
rect 10008 13132 10014 13144
rect 10045 13141 10057 13144
rect 10091 13141 10103 13175
rect 10045 13135 10103 13141
rect 15746 13132 15752 13184
rect 15804 13172 15810 13184
rect 17788 13172 17816 13271
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 21634 13308 21640 13320
rect 21595 13280 21640 13308
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 21744 13308 21772 13348
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 22278 13376 22284 13388
rect 21959 13348 22284 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22278 13336 22284 13348
rect 22336 13336 22342 13388
rect 26252 13376 26280 13475
rect 26513 13379 26571 13385
rect 26513 13376 26525 13379
rect 26252 13348 26525 13376
rect 26513 13345 26525 13348
rect 26559 13345 26571 13379
rect 26786 13376 26792 13388
rect 26747 13348 26792 13376
rect 26513 13339 26571 13345
rect 26786 13336 26792 13348
rect 26844 13336 26850 13388
rect 23017 13311 23075 13317
rect 23017 13308 23029 13311
rect 21744 13280 23029 13308
rect 23017 13277 23029 13280
rect 23063 13277 23075 13311
rect 23017 13271 23075 13277
rect 23308 13212 26372 13240
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 15804 13144 18429 13172
rect 15804 13132 15810 13144
rect 18417 13141 18429 13144
rect 18463 13172 18475 13175
rect 23308 13172 23336 13212
rect 18463 13144 23336 13172
rect 26344 13172 26372 13212
rect 27614 13172 27620 13184
rect 26344 13144 27620 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 27798 13132 27804 13184
rect 27856 13172 27862 13184
rect 28077 13175 28135 13181
rect 28077 13172 28089 13175
rect 27856 13144 28089 13172
rect 27856 13132 27862 13144
rect 28077 13141 28089 13144
rect 28123 13172 28135 13175
rect 31754 13172 31760 13184
rect 28123 13144 31760 13172
rect 28123 13141 28135 13144
rect 28077 13135 28135 13141
rect 31754 13132 31760 13144
rect 31812 13132 31818 13184
rect 1104 13082 29256 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 29256 13082
rect 1104 13008 29256 13030
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4614 12968 4620 12980
rect 4479 12940 4620 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 7892 12940 8677 12968
rect 7892 12928 7898 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 8665 12931 8723 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 9824 12940 10425 12968
rect 9824 12928 9830 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 15473 12971 15531 12977
rect 15473 12968 15485 12971
rect 15252 12940 15485 12968
rect 15252 12928 15258 12940
rect 15473 12937 15485 12940
rect 15519 12937 15531 12971
rect 15746 12968 15752 12980
rect 15707 12940 15752 12968
rect 15473 12931 15531 12937
rect 8202 12900 8208 12912
rect 8115 12872 8208 12900
rect 8202 12860 8208 12872
rect 8260 12900 8266 12912
rect 9784 12900 9812 12928
rect 8260 12872 9812 12900
rect 15488 12900 15516 12931
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 24302 12968 24308 12980
rect 24263 12940 24308 12968
rect 24302 12928 24308 12940
rect 24360 12928 24366 12980
rect 17954 12900 17960 12912
rect 15488 12872 17960 12900
rect 8260 12860 8266 12872
rect 17954 12860 17960 12872
rect 18012 12860 18018 12912
rect 2590 12832 2596 12844
rect 2551 12804 2596 12832
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 4890 12832 4896 12844
rect 2915 12804 4896 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 24320 12832 24348 12928
rect 24489 12835 24547 12841
rect 24489 12832 24501 12835
rect 24320 12804 24501 12832
rect 24489 12801 24501 12804
rect 24535 12832 24547 12835
rect 24535 12804 25084 12832
rect 24535 12801 24547 12804
rect 24489 12795 24547 12801
rect 25056 12776 25084 12804
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 9122 12764 9128 12776
rect 8527 12736 9128 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 9122 12724 9128 12736
rect 9180 12724 9186 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 14826 12764 14832 12776
rect 10735 12736 14832 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 15378 12764 15384 12776
rect 15291 12736 15384 12764
rect 15378 12724 15384 12736
rect 15436 12764 15442 12776
rect 15746 12764 15752 12776
rect 15436 12736 15752 12764
rect 15436 12724 15442 12736
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 24854 12764 24860 12776
rect 24811 12736 24860 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25038 12724 25044 12776
rect 25096 12724 25102 12776
rect 8386 12696 8392 12708
rect 8347 12668 8392 12696
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 10597 12699 10655 12705
rect 10597 12665 10609 12699
rect 10643 12665 10655 12699
rect 11146 12696 11152 12708
rect 11107 12668 11152 12696
rect 10597 12659 10655 12665
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 10612 12628 10640 12659
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 11054 12628 11060 12640
rect 10612 12600 11060 12628
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 25866 12628 25872 12640
rect 25827 12600 25872 12628
rect 25866 12588 25872 12600
rect 25924 12588 25930 12640
rect 1104 12538 29256 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 29256 12538
rect 1104 12464 29256 12486
rect 7282 12424 7288 12436
rect 7243 12396 7288 12424
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 10594 12424 10600 12436
rect 10555 12396 10600 12424
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11977 12427 12035 12433
rect 11977 12424 11989 12427
rect 11112 12396 11989 12424
rect 11112 12384 11118 12396
rect 11977 12393 11989 12396
rect 12023 12393 12035 12427
rect 11977 12387 12035 12393
rect 20254 12384 20260 12436
rect 20312 12424 20318 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 20312 12396 22661 12424
rect 20312 12384 20318 12396
rect 22649 12393 22661 12396
rect 22695 12393 22707 12427
rect 22830 12424 22836 12436
rect 22791 12396 22836 12424
rect 22649 12387 22707 12393
rect 10321 12359 10379 12365
rect 10321 12356 10333 12359
rect 7024 12328 10333 12356
rect 7024 12300 7052 12328
rect 10321 12325 10333 12328
rect 10367 12356 10379 12359
rect 11701 12359 11759 12365
rect 11701 12356 11713 12359
rect 10367 12328 11713 12356
rect 10367 12325 10379 12328
rect 10321 12319 10379 12325
rect 11701 12325 11713 12328
rect 11747 12356 11759 12359
rect 12526 12356 12532 12368
rect 11747 12328 12532 12356
rect 11747 12325 11759 12328
rect 11701 12319 11759 12325
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 4982 12288 4988 12300
rect 3384 12260 4988 12288
rect 3384 12248 3390 12260
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 7006 12288 7012 12300
rect 6967 12260 7012 12288
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12288 7251 12291
rect 7466 12288 7472 12300
rect 7239 12260 7472 12288
rect 7239 12257 7251 12260
rect 7193 12251 7251 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 11422 12288 11428 12300
rect 10551 12260 11428 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 11885 12291 11943 12297
rect 11885 12257 11897 12291
rect 11931 12288 11943 12291
rect 13814 12288 13820 12300
rect 11931 12260 13820 12288
rect 11931 12257 11943 12260
rect 11885 12251 11943 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 17236 12260 18981 12288
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 17236 12229 17264 12260
rect 18969 12257 18981 12260
rect 19015 12288 19027 12291
rect 20622 12288 20628 12300
rect 19015 12260 20628 12288
rect 19015 12257 19027 12260
rect 18969 12251 19027 12257
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 22664 12288 22692 12387
rect 22830 12384 22836 12396
rect 22888 12384 22894 12436
rect 23017 12291 23075 12297
rect 23017 12288 23029 12291
rect 22664 12260 23029 12288
rect 23017 12257 23029 12260
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 17221 12223 17279 12229
rect 17221 12220 17233 12223
rect 13780 12192 17233 12220
rect 13780 12180 13786 12192
rect 17221 12189 17233 12192
rect 17267 12189 17279 12223
rect 17494 12220 17500 12232
rect 17455 12192 17500 12220
rect 17221 12183 17279 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12220 18935 12223
rect 20070 12220 20076 12232
rect 18923 12192 20076 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 1104 11994 29256 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 29256 11994
rect 1104 11920 29256 11942
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8481 11883 8539 11889
rect 8481 11880 8493 11883
rect 8444 11852 8493 11880
rect 8444 11840 8450 11852
rect 8481 11849 8493 11852
rect 8527 11849 8539 11883
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 8481 11843 8539 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 20070 11880 20076 11892
rect 19475 11852 20076 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 17954 11812 17960 11824
rect 16868 11784 17960 11812
rect 2590 11744 2596 11756
rect 2551 11716 2596 11744
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 11146 11744 11152 11756
rect 2915 11716 11152 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 13722 11744 13728 11756
rect 12483 11716 13728 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 13722 11704 13728 11716
rect 13780 11744 13786 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13780 11716 14197 11744
rect 13780 11704 13786 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7064 11648 8217 11676
rect 7064 11636 7070 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8386 11676 8392 11688
rect 8347 11648 8392 11676
rect 8205 11639 8263 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 12710 11676 12716 11688
rect 12671 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 16868 11685 16896 11784
rect 17954 11772 17960 11784
rect 18012 11812 18018 11824
rect 19150 11812 19156 11824
rect 18012 11784 19156 11812
rect 18012 11772 18018 11784
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17552 11716 18061 11744
rect 17552 11704 17558 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 19444 11744 19472 11843
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 25038 11880 25044 11892
rect 24999 11852 25044 11880
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 20990 11744 20996 11756
rect 18049 11707 18107 11713
rect 18708 11716 19472 11744
rect 20951 11716 20996 11744
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11645 16911 11679
rect 18506 11676 18512 11688
rect 18467 11648 18512 11676
rect 16853 11639 16911 11645
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18708 11685 18736 11716
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 25056 11744 25084 11840
rect 25225 11747 25283 11753
rect 25225 11744 25237 11747
rect 25056 11716 25237 11744
rect 25225 11713 25237 11716
rect 25271 11713 25283 11747
rect 25225 11707 25283 11713
rect 25501 11747 25559 11753
rect 25501 11713 25513 11747
rect 25547 11744 25559 11747
rect 25866 11744 25872 11756
rect 25547 11716 25872 11744
rect 25547 11713 25559 11716
rect 25501 11707 25559 11713
rect 25866 11704 25872 11716
rect 25924 11704 25930 11756
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 19015 11679 19073 11685
rect 19015 11676 19027 11679
rect 18693 11639 18751 11645
rect 18892 11648 19027 11676
rect 18892 11608 18920 11648
rect 19015 11645 19027 11648
rect 19061 11645 19073 11679
rect 19150 11676 19156 11688
rect 19111 11648 19156 11676
rect 19015 11639 19073 11645
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 20622 11608 20628 11620
rect 18892 11580 20628 11608
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4433 11543 4491 11549
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 4614 11540 4620 11552
rect 4479 11512 4620 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 17034 11540 17040 11552
rect 16995 11512 17040 11540
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 21634 11540 21640 11552
rect 21595 11512 21640 11540
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 26418 11500 26424 11552
rect 26476 11540 26482 11552
rect 26605 11543 26663 11549
rect 26605 11540 26617 11543
rect 26476 11512 26617 11540
rect 26476 11500 26482 11512
rect 26605 11509 26617 11512
rect 26651 11509 26663 11543
rect 26605 11503 26663 11509
rect 1104 11450 29256 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 29256 11450
rect 1104 11376 29256 11398
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 13872 11308 14320 11336
rect 13872 11296 13878 11308
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12768 11240 13185 11268
rect 12768 11228 12774 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 14292 11209 14320 11308
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 4672 11172 5641 11200
rect 4672 11160 4678 11172
rect 5629 11169 5641 11172
rect 5675 11200 5687 11203
rect 13817 11203 13875 11209
rect 5675 11172 7052 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 6914 11132 6920 11144
rect 5951 11104 6920 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7024 11064 7052 11172
rect 13817 11169 13829 11203
rect 13863 11169 13875 11203
rect 13817 11163 13875 11169
rect 14185 11203 14243 11209
rect 14185 11169 14197 11203
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11200 14611 11203
rect 15378 11200 15384 11212
rect 14599 11172 15384 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7466 11132 7472 11144
rect 7331 11104 7472 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 7374 11064 7380 11076
rect 7024 11036 7380 11064
rect 7374 11024 7380 11036
rect 7432 11064 7438 11076
rect 8846 11064 8852 11076
rect 7432 11036 8852 11064
rect 7432 11024 7438 11036
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 13832 10996 13860 11163
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11101 13967 11135
rect 14200 11132 14228 11163
rect 14568 11132 14596 11163
rect 15378 11160 15384 11172
rect 15436 11200 15442 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15436 11172 15945 11200
rect 15436 11160 15442 11172
rect 15933 11169 15945 11172
rect 15979 11200 15991 11203
rect 16301 11203 16359 11209
rect 16301 11200 16313 11203
rect 15979 11172 16313 11200
rect 15979 11169 15991 11172
rect 15933 11163 15991 11169
rect 16301 11169 16313 11172
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 14200 11104 14596 11132
rect 13909 11095 13967 11101
rect 13924 11064 13952 11095
rect 14734 11092 14740 11144
rect 14792 11132 14798 11144
rect 17034 11132 17040 11144
rect 14792 11104 17040 11132
rect 14792 11092 14798 11104
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 15194 11064 15200 11076
rect 13924 11036 15200 11064
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 16114 11064 16120 11076
rect 16027 11036 16120 11064
rect 16114 11024 16120 11036
rect 16172 11064 16178 11076
rect 18506 11064 18512 11076
rect 16172 11036 18512 11064
rect 16172 11024 16178 11036
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 14734 10996 14740 11008
rect 8536 10968 14740 10996
rect 8536 10956 8542 10968
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 1104 10906 29256 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 29256 10906
rect 1104 10832 29256 10854
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4028 10764 8340 10792
rect 4028 10752 4034 10764
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 4614 10724 4620 10736
rect 4479 10696 4620 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 8312 10724 8340 10764
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 8444 10764 8769 10792
rect 8444 10752 8450 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 8904 10764 9229 10792
rect 8904 10752 8910 10764
rect 9217 10761 9229 10764
rect 9263 10792 9275 10795
rect 12618 10792 12624 10804
rect 9263 10764 12624 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 20680 10764 22017 10792
rect 20680 10752 20686 10764
rect 22005 10761 22017 10764
rect 22051 10761 22063 10795
rect 22005 10755 22063 10761
rect 11238 10724 11244 10736
rect 8312 10696 11244 10724
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 2590 10656 2596 10668
rect 2551 10628 2596 10656
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 7834 10656 7840 10668
rect 2915 10628 7840 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 14277 10659 14335 10665
rect 11480 10628 14228 10656
rect 11480 10616 11486 10628
rect 2608 10588 2636 10616
rect 4614 10588 4620 10600
rect 2608 10560 4620 10588
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 7374 10588 7380 10600
rect 7335 10560 7380 10588
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7650 10588 7656 10600
rect 7611 10560 7656 10588
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 8110 10548 8116 10600
rect 8168 10588 8174 10600
rect 8168 10560 13860 10588
rect 8168 10548 8174 10560
rect 12986 10480 12992 10532
rect 13044 10520 13050 10532
rect 13541 10523 13599 10529
rect 13541 10520 13553 10523
rect 13044 10492 13553 10520
rect 13044 10480 13050 10492
rect 13541 10489 13553 10492
rect 13587 10489 13599 10523
rect 13832 10520 13860 10560
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14200 10597 14228 10628
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 16114 10656 16120 10668
rect 14323 10628 16120 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 14148 10560 14197 10588
rect 14148 10548 14154 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14292 10520 14320 10619
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10656 26111 10659
rect 26418 10656 26424 10668
rect 26099 10628 26424 10656
rect 26099 10625 26111 10628
rect 26053 10619 26111 10625
rect 26418 10616 26424 10628
rect 26476 10616 26482 10668
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 14734 10588 14740 10600
rect 14695 10560 14740 10588
rect 14553 10551 14611 10557
rect 13832 10492 14320 10520
rect 14568 10520 14596 10551
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 20625 10591 20683 10597
rect 20625 10588 20637 10591
rect 20456 10560 20637 10588
rect 15286 10520 15292 10532
rect 14568 10492 15292 10520
rect 13541 10483 13599 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 20456 10464 20484 10560
rect 20625 10557 20637 10560
rect 20671 10557 20683 10591
rect 20898 10588 20904 10600
rect 20859 10560 20904 10588
rect 20625 10551 20683 10557
rect 20898 10548 20904 10560
rect 20956 10548 20962 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25608 10560 25789 10588
rect 25608 10464 25636 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 4154 10452 4160 10464
rect 4115 10424 4160 10452
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 26786 10412 26792 10464
rect 26844 10452 26850 10464
rect 27157 10455 27215 10461
rect 27157 10452 27169 10455
rect 26844 10424 27169 10452
rect 26844 10412 26850 10424
rect 27157 10421 27169 10424
rect 27203 10421 27215 10455
rect 27157 10415 27215 10421
rect 1104 10362 29256 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 29256 10362
rect 1104 10288 29256 10310
rect 7650 10248 7656 10260
rect 7611 10220 7656 10248
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 14090 10248 14096 10260
rect 14051 10220 14096 10248
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 20956 10220 22293 10248
rect 20956 10208 20962 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 27614 10208 27620 10260
rect 27672 10248 27678 10260
rect 27893 10251 27951 10257
rect 27893 10248 27905 10251
rect 27672 10220 27905 10248
rect 27672 10208 27678 10220
rect 27893 10217 27905 10220
rect 27939 10217 27951 10251
rect 27893 10211 27951 10217
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8386 10112 8392 10124
rect 8251 10084 8392 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9858 10112 9864 10124
rect 8619 10084 9864 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 12636 10112 12664 10208
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 12636 10084 12725 10112
rect 12713 10081 12725 10084
rect 12759 10081 12771 10115
rect 12986 10112 12992 10124
rect 12947 10084 12992 10112
rect 12713 10075 12771 10081
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 21177 10115 21235 10121
rect 19935 10084 21036 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8478 10044 8484 10056
rect 8439 10016 8484 10044
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20640 10016 20913 10044
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19705 9911 19763 9917
rect 19705 9908 19717 9911
rect 19392 9880 19717 9908
rect 19392 9868 19398 9880
rect 19705 9877 19717 9880
rect 19751 9908 19763 9911
rect 20438 9908 20444 9920
rect 19751 9880 20444 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20438 9868 20444 9880
rect 20496 9908 20502 9920
rect 20640 9917 20668 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 21008 10044 21036 10084
rect 21177 10081 21189 10115
rect 21223 10112 21235 10115
rect 21266 10112 21272 10124
rect 21223 10084 21272 10112
rect 21223 10081 21235 10084
rect 21177 10075 21235 10081
rect 21266 10072 21272 10084
rect 21324 10112 21330 10124
rect 21634 10112 21640 10124
rect 21324 10084 21640 10112
rect 21324 10072 21330 10084
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 26786 10112 26792 10124
rect 26747 10084 26792 10112
rect 26786 10072 26792 10084
rect 26844 10072 26850 10124
rect 22830 10044 22836 10056
rect 21008 10016 22836 10044
rect 20901 10007 20959 10013
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10044 26387 10047
rect 26513 10047 26571 10053
rect 26513 10044 26525 10047
rect 26375 10016 26525 10044
rect 26375 10013 26387 10016
rect 26329 10007 26387 10013
rect 26513 10013 26525 10016
rect 26559 10013 26571 10047
rect 26513 10007 26571 10013
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 20496 9880 20637 9908
rect 20496 9868 20502 9880
rect 20625 9877 20637 9880
rect 20671 9877 20683 9911
rect 20625 9871 20683 9877
rect 25590 9868 25596 9920
rect 25648 9908 25654 9920
rect 26344 9908 26372 10007
rect 25648 9880 26372 9908
rect 25648 9868 25654 9880
rect 1104 9818 29256 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 29256 9818
rect 1104 9744 29256 9766
rect 15286 9704 15292 9716
rect 15247 9676 15292 9704
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 19426 9636 19432 9648
rect 19339 9608 19432 9636
rect 19426 9596 19432 9608
rect 19484 9636 19490 9648
rect 19886 9636 19892 9648
rect 19484 9608 19892 9636
rect 19484 9596 19490 9608
rect 19886 9596 19892 9608
rect 19944 9596 19950 9648
rect 6914 9568 6920 9580
rect 6875 9540 6920 9568
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 8110 9568 8116 9580
rect 7607 9540 8116 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 13722 9568 13728 9580
rect 13683 9540 13728 9568
rect 13722 9528 13728 9540
rect 13780 9568 13786 9580
rect 15473 9571 15531 9577
rect 15473 9568 15485 9571
rect 13780 9540 15485 9568
rect 13780 9528 13786 9540
rect 15473 9537 15485 9540
rect 15519 9568 15531 9571
rect 17770 9568 17776 9580
rect 15519 9540 17776 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18506 9568 18512 9580
rect 18467 9540 18512 9568
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 19444 9568 19472 9596
rect 21266 9568 21272 9580
rect 18708 9540 19472 9568
rect 21227 9540 21272 9568
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7834 9500 7840 9512
rect 7795 9472 7840 9500
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8478 9500 8484 9512
rect 8067 9472 8484 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 13998 9500 14004 9512
rect 13959 9472 14004 9500
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 18708 9509 18736 9540
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 18693 9503 18751 9509
rect 17092 9472 18184 9500
rect 17092 9460 17098 9472
rect 18046 9432 18052 9444
rect 18007 9404 18052 9432
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 18156 9432 18184 9472
rect 18693 9469 18705 9503
rect 18739 9469 18751 9503
rect 19058 9500 19064 9512
rect 19019 9472 19064 9500
rect 18693 9463 18751 9469
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 19153 9503 19211 9509
rect 19153 9469 19165 9503
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 19168 9432 19196 9463
rect 18156 9404 19196 9432
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 7742 9364 7748 9376
rect 3568 9336 7748 9364
rect 3568 9324 3574 9336
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 21913 9367 21971 9373
rect 21913 9333 21925 9367
rect 21959 9364 21971 9367
rect 22186 9364 22192 9376
rect 21959 9336 22192 9364
rect 21959 9333 21971 9336
rect 21913 9327 21971 9333
rect 22186 9324 22192 9336
rect 22244 9324 22250 9376
rect 1104 9274 29256 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 29256 9274
rect 1104 9200 29256 9222
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 7834 9160 7840 9172
rect 6595 9132 7840 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 6825 9095 6883 9101
rect 6825 9061 6837 9095
rect 6871 9092 6883 9095
rect 7374 9092 7380 9104
rect 6871 9064 7380 9092
rect 6871 9061 6883 9064
rect 6825 9055 6883 9061
rect 4982 9024 4988 9036
rect 4895 8996 4988 9024
rect 4982 8984 4988 8996
rect 5040 9024 5046 9036
rect 6840 9024 6868 9055
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 19426 9092 19432 9104
rect 19387 9064 19432 9092
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 17770 9024 17776 9036
rect 5040 8996 6868 9024
rect 17731 8996 17776 9024
rect 5040 8984 5046 8996
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 18046 9024 18052 9036
rect 18007 8996 18052 9024
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5626 8956 5632 8968
rect 5307 8928 5632 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 17788 8956 17816 8984
rect 19334 8956 19340 8968
rect 17788 8928 19340 8956
rect 19334 8916 19340 8928
rect 19392 8956 19398 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19392 8928 19533 8956
rect 19392 8916 19398 8928
rect 19521 8925 19533 8928
rect 19567 8956 19579 8959
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 19567 8928 21741 8956
rect 19567 8925 19579 8928
rect 19521 8919 19579 8925
rect 21729 8925 21741 8928
rect 21775 8956 21787 8959
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21775 8928 21925 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 21913 8925 21925 8928
rect 21959 8925 21971 8959
rect 22186 8956 22192 8968
rect 22147 8928 22192 8956
rect 21913 8919 21971 8925
rect 21928 8820 21956 8919
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22278 8820 22284 8832
rect 21928 8792 22284 8820
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 23477 8823 23535 8829
rect 23477 8789 23489 8823
rect 23523 8820 23535 8823
rect 23934 8820 23940 8832
rect 23523 8792 23940 8820
rect 23523 8789 23535 8792
rect 23477 8783 23535 8789
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 1104 8730 29256 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 29256 8730
rect 1104 8656 29256 8678
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 4982 8616 4988 8628
rect 4479 8588 4988 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 14056 8588 14197 8616
rect 14056 8576 14062 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 25041 8619 25099 8625
rect 25041 8616 25053 8619
rect 19116 8588 25053 8616
rect 19116 8576 19122 8588
rect 25041 8585 25053 8588
rect 25087 8585 25099 8619
rect 25041 8579 25099 8585
rect 2590 8480 2596 8492
rect 2551 8452 2596 8480
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 7098 8480 7104 8492
rect 2915 8452 7104 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 7432 8452 8493 8480
rect 7432 8440 7438 8452
rect 8481 8449 8493 8452
rect 8527 8480 8539 8483
rect 9766 8480 9772 8492
rect 8527 8452 9772 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 9766 8440 9772 8452
rect 9824 8480 9830 8492
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 9824 8452 10241 8480
rect 9824 8440 9830 8452
rect 10229 8449 10241 8452
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 11112 8452 13093 8480
rect 11112 8440 11118 8452
rect 13081 8449 13093 8452
rect 13127 8480 13139 8483
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 13127 8452 21465 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 23934 8480 23940 8492
rect 23895 8452 23940 8480
rect 21453 8443 21511 8449
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 8754 8412 8760 8424
rect 8715 8384 8760 8412
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12676 8384 12817 8412
rect 12676 8372 12682 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 20809 8415 20867 8421
rect 20809 8381 20821 8415
rect 20855 8412 20867 8415
rect 22186 8412 22192 8424
rect 20855 8384 22192 8412
rect 20855 8381 20867 8384
rect 20809 8375 20867 8381
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 22278 8372 22284 8424
rect 22336 8412 22342 8424
rect 23477 8415 23535 8421
rect 23477 8412 23489 8415
rect 22336 8384 23489 8412
rect 22336 8372 22342 8384
rect 23477 8381 23489 8384
rect 23523 8412 23535 8415
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23523 8384 23673 8412
rect 23523 8381 23535 8384
rect 23477 8375 23535 8381
rect 23661 8381 23673 8384
rect 23707 8412 23719 8415
rect 25590 8412 25596 8424
rect 23707 8384 25596 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 25590 8372 25596 8384
rect 25648 8372 25654 8424
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 1104 8186 29256 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 29256 8186
rect 1104 8112 29256 8134
rect 5626 8072 5632 8084
rect 5587 8044 5632 8072
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 5905 8075 5963 8081
rect 5905 8041 5917 8075
rect 5951 8072 5963 8075
rect 7374 8072 7380 8084
rect 5951 8044 7380 8072
rect 5951 8041 5963 8044
rect 5905 8035 5963 8041
rect 4062 7936 4068 7948
rect 3975 7908 4068 7936
rect 4062 7896 4068 7908
rect 4120 7936 4126 7948
rect 5920 7936 5948 8035
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 4120 7908 5948 7936
rect 8021 7939 8079 7945
rect 4120 7896 4126 7908
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 11054 7936 11060 7948
rect 8067 7908 11060 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 8110 7868 8116 7880
rect 4387 7840 8116 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 8110 7828 8116 7840
rect 8168 7868 8174 7880
rect 8665 7871 8723 7877
rect 8665 7868 8677 7871
rect 8168 7840 8677 7868
rect 8168 7828 8174 7840
rect 8665 7837 8677 7840
rect 8711 7837 8723 7871
rect 8665 7831 8723 7837
rect 1104 7642 29256 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 29256 7642
rect 1104 7568 29256 7590
rect 4062 7528 4068 7540
rect 2608 7500 4068 7528
rect 2608 7401 2636 7500
rect 4062 7488 4068 7500
rect 4120 7528 4126 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4120 7500 4353 7528
rect 4120 7488 4126 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 8754 7488 8760 7540
rect 8812 7528 8818 7540
rect 9217 7531 9275 7537
rect 9217 7528 9229 7531
rect 8812 7500 9229 7528
rect 8812 7488 8818 7500
rect 9217 7497 9229 7500
rect 9263 7497 9275 7531
rect 9217 7491 9275 7497
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 9766 7528 9772 7540
rect 9723 7500 9772 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 15194 7528 15200 7540
rect 15155 7500 15200 7528
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3694 7392 3700 7404
rect 2915 7364 3700 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7432 7364 7849 7392
rect 7432 7352 7438 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8754 7324 8760 7336
rect 8159 7296 8760 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8754 7284 8760 7296
rect 8812 7324 8818 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 8812 7296 10793 7324
rect 8812 7284 8818 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7293 13691 7327
rect 13906 7324 13912 7336
rect 13867 7296 13912 7324
rect 13633 7287 13691 7293
rect 9766 7216 9772 7268
rect 9824 7256 9830 7268
rect 12066 7256 12072 7268
rect 9824 7228 12072 7256
rect 9824 7216 9830 7228
rect 12066 7216 12072 7228
rect 12124 7256 12130 7268
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 12124 7228 13461 7256
rect 12124 7216 12130 7228
rect 13449 7225 13461 7228
rect 13495 7256 13507 7259
rect 13648 7256 13676 7287
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 13495 7228 13676 7256
rect 13495 7225 13507 7228
rect 13449 7219 13507 7225
rect 4154 7188 4160 7200
rect 4115 7160 4160 7188
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 11425 7191 11483 7197
rect 11425 7157 11437 7191
rect 11471 7188 11483 7191
rect 12526 7188 12532 7200
rect 11471 7160 12532 7188
rect 11471 7157 11483 7160
rect 11425 7151 11483 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 1104 7098 29256 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 29256 7098
rect 1104 7024 29256 7046
rect 13906 6916 13912 6928
rect 13867 6888 13912 6916
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8110 6848 8116 6860
rect 8067 6820 8116 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 8754 6848 8760 6860
rect 8711 6820 8760 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 12066 6848 12072 6860
rect 12027 6820 12072 6848
rect 12066 6808 12072 6820
rect 12124 6848 12130 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12124 6820 12265 6848
rect 12124 6808 12130 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 12526 6848 12532 6860
rect 12487 6820 12532 6848
rect 12253 6811 12311 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 6546 6780 6552 6792
rect 4028 6752 6552 6780
rect 4028 6740 4034 6752
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 1104 6554 29256 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 29256 6554
rect 1104 6480 29256 6502
rect 3878 6440 3884 6452
rect 3160 6412 3884 6440
rect 3160 6313 3188 6412
rect 3878 6400 3884 6412
rect 3936 6440 3942 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 3936 6412 4905 6440
rect 3936 6400 3942 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 4893 6403 4951 6409
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 8570 6304 8576 6316
rect 3467 6276 8576 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4212 6072 4537 6100
rect 4212 6060 4218 6072
rect 4525 6069 4537 6072
rect 4571 6069 4583 6103
rect 4525 6063 4583 6069
rect 1104 6010 29256 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 29256 6010
rect 1104 5936 29256 5958
rect 1104 5466 29256 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 29256 5466
rect 1104 5392 29256 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 4798 5352 4804 5364
rect 3016 5324 4804 5352
rect 3016 5312 3022 5324
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 26326 5352 26332 5364
rect 26287 5324 26332 5352
rect 26326 5312 26332 5324
rect 26384 5312 26390 5364
rect 25590 5244 25596 5296
rect 25648 5284 25654 5296
rect 26053 5287 26111 5293
rect 26053 5284 26065 5287
rect 25648 5256 26065 5284
rect 25648 5244 25654 5256
rect 26053 5253 26065 5256
rect 26099 5253 26111 5287
rect 26053 5247 26111 5253
rect 26068 5148 26096 5247
rect 26344 5216 26372 5312
rect 26697 5219 26755 5225
rect 26697 5216 26709 5219
rect 26344 5188 26709 5216
rect 26697 5185 26709 5188
rect 26743 5185 26755 5219
rect 26697 5179 26755 5185
rect 26421 5151 26479 5157
rect 26421 5148 26433 5151
rect 26068 5120 26433 5148
rect 26421 5117 26433 5120
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 28077 5083 28135 5089
rect 28077 5049 28089 5083
rect 28123 5080 28135 5083
rect 29914 5080 29920 5092
rect 28123 5052 29920 5080
rect 28123 5049 28135 5052
rect 28077 5043 28135 5049
rect 29914 5040 29920 5052
rect 29972 5040 29978 5092
rect 1104 4922 29256 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 29256 4922
rect 1104 4848 29256 4870
rect 11517 4811 11575 4817
rect 11517 4808 11529 4811
rect 9692 4780 11529 4808
rect 9692 4681 9720 4780
rect 11517 4777 11529 4780
rect 11563 4808 11575 4811
rect 12066 4808 12072 4820
rect 11563 4780 12072 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9677 4635 9735 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 1104 4378 29256 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 29256 4378
rect 1104 4304 29256 4326
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 3927 4100 5457 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 5445 4097 5457 4100
rect 5491 4128 5503 4131
rect 5902 4128 5908 4140
rect 5491 4100 5908 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 3970 4060 3976 4072
rect 3651 4032 3976 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 3970 4020 3976 4032
rect 4028 4060 4034 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 4028 4032 5549 4060
rect 4028 4020 4034 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 1104 3834 29256 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 29256 3834
rect 1104 3760 29256 3782
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 11054 3720 11060 3732
rect 4120 3692 11060 3720
rect 4120 3680 4126 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 7926 3652 7932 3664
rect 3384 3624 7932 3652
rect 3384 3612 3390 3624
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 1104 3290 29256 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 29256 3290
rect 1104 3216 29256 3238
rect 4706 3176 4712 3188
rect 4667 3148 4712 3176
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 4724 3040 4752 3136
rect 3283 3012 4752 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3970 2972 3976 2984
rect 3007 2944 3976 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3970 2932 3976 2944
rect 4028 2972 4034 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4028 2944 4905 2972
rect 4028 2932 4034 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 4341 2839 4399 2845
rect 4341 2836 4353 2839
rect 2832 2808 4353 2836
rect 2832 2796 2838 2808
rect 4341 2805 4353 2808
rect 4387 2805 4399 2839
rect 4341 2799 4399 2805
rect 1104 2746 29256 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 29256 2746
rect 1104 2672 29256 2694
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 4982 2292 4988 2304
rect 2924 2264 4988 2292
rect 2924 2252 2930 2264
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 1104 2202 29256 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 29256 2202
rect 1104 2128 29256 2150
rect 3234 1708 3240 1760
rect 3292 1748 3298 1760
rect 8018 1748 8024 1760
rect 3292 1720 8024 1748
rect 3292 1708 3298 1720
rect 8018 1708 8024 1720
rect 8076 1708 8082 1760
rect 3418 688 3424 740
rect 3476 728 3482 740
rect 8202 728 8208 740
rect 3476 700 8208 728
rect 3476 688 3482 700
rect 8202 688 8208 700
rect 8260 688 8266 740
<< via1 >>
rect 4068 48356 4120 48408
rect 14924 48356 14976 48408
rect 3976 48288 4028 48340
rect 73068 48288 73120 48340
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 65686 47846 65738 47898
rect 65750 47846 65802 47898
rect 65814 47846 65866 47898
rect 65878 47846 65930 47898
rect 96406 47846 96458 47898
rect 96470 47846 96522 47898
rect 96534 47846 96586 47898
rect 96598 47846 96650 47898
rect 8392 47651 8444 47660
rect 8392 47617 8401 47651
rect 8401 47617 8435 47651
rect 8435 47617 8444 47651
rect 8392 47608 8444 47617
rect 7932 47583 7984 47592
rect 7932 47549 7941 47583
rect 7941 47549 7975 47583
rect 7975 47549 7984 47583
rect 7932 47540 7984 47549
rect 13728 47540 13780 47592
rect 12072 47404 12124 47456
rect 22468 47404 22520 47456
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 50326 47302 50378 47354
rect 50390 47302 50442 47354
rect 50454 47302 50506 47354
rect 50518 47302 50570 47354
rect 81046 47302 81098 47354
rect 81110 47302 81162 47354
rect 81174 47302 81226 47354
rect 81238 47302 81290 47354
rect 3424 47064 3476 47116
rect 7932 47107 7984 47116
rect 7932 47073 7941 47107
rect 7941 47073 7975 47107
rect 7975 47073 7984 47107
rect 7932 47064 7984 47073
rect 22284 47200 22336 47252
rect 22468 47243 22520 47252
rect 22468 47209 22477 47243
rect 22477 47209 22511 47243
rect 22511 47209 22520 47243
rect 22468 47200 22520 47209
rect 12072 46971 12124 46980
rect 4712 46860 4764 46912
rect 12072 46937 12081 46971
rect 12081 46937 12115 46971
rect 12115 46937 12124 46971
rect 13360 46971 13412 46980
rect 12072 46928 12124 46937
rect 13360 46937 13369 46971
rect 13369 46937 13403 46971
rect 13403 46937 13412 46971
rect 13360 46928 13412 46937
rect 23296 47132 23348 47184
rect 23388 47107 23440 47116
rect 23388 47073 23397 47107
rect 23397 47073 23431 47107
rect 23431 47073 23440 47107
rect 23388 47064 23440 47073
rect 25412 47107 25464 47116
rect 14004 46928 14056 46980
rect 14188 46971 14240 46980
rect 14188 46937 14197 46971
rect 14197 46937 14231 46971
rect 14231 46937 14240 46971
rect 14188 46928 14240 46937
rect 7196 46860 7248 46912
rect 15476 46860 15528 46912
rect 18052 46996 18104 47048
rect 23388 46928 23440 46980
rect 23940 46928 23992 46980
rect 25412 47073 25421 47107
rect 25421 47073 25455 47107
rect 25455 47073 25464 47107
rect 25412 47064 25464 47073
rect 44364 47064 44416 47116
rect 32588 47039 32640 47048
rect 32588 47005 32597 47039
rect 32597 47005 32631 47039
rect 32631 47005 32640 47039
rect 32588 46996 32640 47005
rect 32864 47039 32916 47048
rect 32864 47005 32873 47039
rect 32873 47005 32907 47039
rect 32907 47005 32916 47039
rect 32864 46996 32916 47005
rect 38752 46971 38804 46980
rect 19064 46860 19116 46912
rect 24032 46860 24084 46912
rect 38752 46937 38761 46971
rect 38761 46937 38795 46971
rect 38795 46937 38804 46971
rect 40592 46996 40644 47048
rect 40684 46996 40736 47048
rect 38752 46928 38804 46937
rect 31024 46860 31076 46912
rect 33784 46860 33836 46912
rect 40040 46860 40092 46912
rect 43444 46903 43496 46912
rect 43444 46869 43453 46903
rect 43453 46869 43487 46903
rect 43487 46869 43496 46903
rect 43444 46860 43496 46869
rect 46664 47064 46716 47116
rect 50160 47064 50212 47116
rect 50528 47064 50580 47116
rect 50896 47107 50948 47116
rect 50896 47073 50905 47107
rect 50905 47073 50939 47107
rect 50939 47073 50948 47107
rect 50896 47064 50948 47073
rect 51908 47064 51960 47116
rect 56692 47107 56744 47116
rect 56692 47073 56701 47107
rect 56701 47073 56735 47107
rect 56735 47073 56744 47107
rect 56692 47064 56744 47073
rect 56784 47107 56836 47116
rect 56784 47073 56793 47107
rect 56793 47073 56827 47107
rect 56827 47073 56836 47107
rect 56784 47064 56836 47073
rect 62948 47064 63000 47116
rect 47308 46996 47360 47048
rect 47492 47039 47544 47048
rect 47492 47005 47501 47039
rect 47501 47005 47535 47039
rect 47535 47005 47544 47039
rect 47492 46996 47544 47005
rect 51356 47039 51408 47048
rect 51356 47005 51365 47039
rect 51365 47005 51399 47039
rect 51399 47005 51408 47039
rect 51356 46996 51408 47005
rect 57244 47039 57296 47048
rect 57244 47005 57253 47039
rect 57253 47005 57287 47039
rect 57287 47005 57296 47039
rect 57244 46996 57296 47005
rect 61476 47039 61528 47048
rect 61476 47005 61485 47039
rect 61485 47005 61519 47039
rect 61519 47005 61528 47039
rect 61476 46996 61528 47005
rect 47400 46928 47452 46980
rect 59544 46928 59596 46980
rect 46480 46903 46532 46912
rect 46480 46869 46489 46903
rect 46489 46869 46523 46903
rect 46523 46869 46532 46903
rect 46480 46860 46532 46869
rect 47308 46860 47360 46912
rect 48688 46860 48740 46912
rect 51724 46860 51776 46912
rect 52368 46903 52420 46912
rect 52368 46869 52377 46903
rect 52377 46869 52411 46903
rect 52411 46869 52420 46903
rect 52368 46860 52420 46869
rect 62120 46860 62172 46912
rect 62948 46903 63000 46912
rect 62948 46869 62957 46903
rect 62957 46869 62991 46903
rect 62991 46869 63000 46903
rect 62948 46860 63000 46869
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 65686 46758 65738 46810
rect 65750 46758 65802 46810
rect 65814 46758 65866 46810
rect 65878 46758 65930 46810
rect 96406 46758 96458 46810
rect 96470 46758 96522 46810
rect 96534 46758 96586 46810
rect 96598 46758 96650 46810
rect 2780 46656 2832 46708
rect 22284 46656 22336 46708
rect 24952 46656 25004 46708
rect 25412 46656 25464 46708
rect 14004 46588 14056 46640
rect 2780 46520 2832 46572
rect 8392 46520 8444 46572
rect 2596 46495 2648 46504
rect 2596 46461 2605 46495
rect 2605 46461 2639 46495
rect 2639 46461 2648 46495
rect 2596 46452 2648 46461
rect 7196 46452 7248 46504
rect 13360 46520 13412 46572
rect 13728 46520 13780 46572
rect 40592 46699 40644 46708
rect 30840 46520 30892 46572
rect 40592 46665 40601 46699
rect 40601 46665 40635 46699
rect 40635 46665 40644 46699
rect 40592 46656 40644 46665
rect 47400 46656 47452 46708
rect 50896 46656 50948 46708
rect 45008 46588 45060 46640
rect 62120 46699 62172 46708
rect 13452 46452 13504 46504
rect 18144 46452 18196 46504
rect 19064 46495 19116 46504
rect 19064 46461 19073 46495
rect 19073 46461 19107 46495
rect 19107 46461 19116 46495
rect 19064 46452 19116 46461
rect 20720 46495 20772 46504
rect 20720 46461 20729 46495
rect 20729 46461 20763 46495
rect 20763 46461 20772 46495
rect 20720 46452 20772 46461
rect 23296 46452 23348 46504
rect 21916 46384 21968 46436
rect 4160 46359 4212 46368
rect 4160 46325 4169 46359
rect 4169 46325 4203 46359
rect 4203 46325 4212 46359
rect 4160 46316 4212 46325
rect 4712 46316 4764 46368
rect 7932 46316 7984 46368
rect 13912 46316 13964 46368
rect 18144 46359 18196 46368
rect 18144 46325 18153 46359
rect 18153 46325 18187 46359
rect 18187 46325 18196 46359
rect 18144 46316 18196 46325
rect 19156 46359 19208 46368
rect 19156 46325 19165 46359
rect 19165 46325 19199 46359
rect 19199 46325 19208 46359
rect 19156 46316 19208 46325
rect 21824 46316 21876 46368
rect 24032 46452 24084 46504
rect 26700 46495 26752 46504
rect 26700 46461 26709 46495
rect 26709 46461 26743 46495
rect 26743 46461 26752 46495
rect 26700 46452 26752 46461
rect 29184 46452 29236 46504
rect 31944 46452 31996 46504
rect 32036 46495 32088 46504
rect 32036 46461 32045 46495
rect 32045 46461 32079 46495
rect 32079 46461 32088 46495
rect 33784 46495 33836 46504
rect 32036 46452 32088 46461
rect 33784 46461 33793 46495
rect 33793 46461 33827 46495
rect 33827 46461 33836 46495
rect 33784 46452 33836 46461
rect 34428 46452 34480 46504
rect 43444 46520 43496 46572
rect 45376 46520 45428 46572
rect 38752 46452 38804 46504
rect 38936 46427 38988 46436
rect 27068 46316 27120 46368
rect 30840 46316 30892 46368
rect 31024 46316 31076 46368
rect 32128 46316 32180 46368
rect 32312 46359 32364 46368
rect 32312 46325 32321 46359
rect 32321 46325 32355 46359
rect 32355 46325 32364 46359
rect 32312 46316 32364 46325
rect 33876 46359 33928 46368
rect 33876 46325 33885 46359
rect 33885 46325 33919 46359
rect 33919 46325 33928 46359
rect 33876 46316 33928 46325
rect 34980 46359 35032 46368
rect 34980 46325 34989 46359
rect 34989 46325 35023 46359
rect 35023 46325 35032 46359
rect 34980 46316 35032 46325
rect 38936 46393 38945 46427
rect 38945 46393 38979 46427
rect 38979 46393 38988 46427
rect 38936 46384 38988 46393
rect 40684 46452 40736 46504
rect 50528 46563 50580 46572
rect 38476 46316 38528 46368
rect 39212 46359 39264 46368
rect 39212 46325 39221 46359
rect 39221 46325 39255 46359
rect 39255 46325 39264 46359
rect 39212 46316 39264 46325
rect 44456 46384 44508 46436
rect 46112 46427 46164 46436
rect 46112 46393 46121 46427
rect 46121 46393 46155 46427
rect 46155 46393 46164 46427
rect 46112 46384 46164 46393
rect 47492 46495 47544 46504
rect 47492 46461 47501 46495
rect 47501 46461 47535 46495
rect 47535 46461 47544 46495
rect 47492 46452 47544 46461
rect 48688 46495 48740 46504
rect 48688 46461 48697 46495
rect 48697 46461 48731 46495
rect 48731 46461 48740 46495
rect 48688 46452 48740 46461
rect 46940 46384 46992 46436
rect 47400 46384 47452 46436
rect 50528 46529 50537 46563
rect 50537 46529 50571 46563
rect 50571 46529 50580 46563
rect 50528 46520 50580 46529
rect 51356 46520 51408 46572
rect 50160 46495 50212 46504
rect 50160 46461 50169 46495
rect 50169 46461 50203 46495
rect 50203 46461 50212 46495
rect 50160 46452 50212 46461
rect 51172 46452 51224 46504
rect 51448 46452 51500 46504
rect 54852 46495 54904 46504
rect 54852 46461 54861 46495
rect 54861 46461 54895 46495
rect 54895 46461 54904 46495
rect 54852 46452 54904 46461
rect 62120 46665 62129 46699
rect 62129 46665 62163 46699
rect 62163 46665 62172 46699
rect 62120 46656 62172 46665
rect 56692 46520 56744 46572
rect 57244 46520 57296 46572
rect 57336 46495 57388 46504
rect 57336 46461 57345 46495
rect 57345 46461 57379 46495
rect 57379 46461 57388 46495
rect 57336 46452 57388 46461
rect 57428 46452 57480 46504
rect 62120 46452 62172 46504
rect 51356 46316 51408 46368
rect 52000 46316 52052 46368
rect 56600 46359 56652 46368
rect 56600 46325 56609 46359
rect 56609 46325 56643 46359
rect 56643 46325 56652 46359
rect 56600 46316 56652 46325
rect 59176 46359 59228 46368
rect 59176 46325 59185 46359
rect 59185 46325 59219 46359
rect 59219 46325 59228 46359
rect 59176 46316 59228 46325
rect 62028 46316 62080 46368
rect 83832 46316 83884 46368
rect 90824 46316 90876 46368
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 50326 46214 50378 46266
rect 50390 46214 50442 46266
rect 50454 46214 50506 46266
rect 50518 46214 50570 46266
rect 81046 46214 81098 46266
rect 81110 46214 81162 46266
rect 81174 46214 81226 46266
rect 81238 46214 81290 46266
rect 4620 46112 4672 46164
rect 14004 46155 14056 46164
rect 14004 46121 14013 46155
rect 14013 46121 14047 46155
rect 14047 46121 14056 46155
rect 14004 46112 14056 46121
rect 7104 45976 7156 46028
rect 8024 46019 8076 46028
rect 8024 45985 8033 46019
rect 8033 45985 8067 46019
rect 8067 45985 8076 46019
rect 8024 45976 8076 45985
rect 13912 46019 13964 46028
rect 13912 45985 13921 46019
rect 13921 45985 13955 46019
rect 13955 45985 13964 46019
rect 13912 45976 13964 45985
rect 14188 45976 14240 46028
rect 23388 46112 23440 46164
rect 26700 46112 26752 46164
rect 19156 45976 19208 46028
rect 18052 45951 18104 45960
rect 16764 45883 16816 45892
rect 16764 45849 16773 45883
rect 16773 45849 16807 45883
rect 16807 45849 16816 45883
rect 18052 45917 18061 45951
rect 18061 45917 18095 45951
rect 18095 45917 18104 45951
rect 18052 45908 18104 45917
rect 20720 45976 20772 46028
rect 22652 46044 22704 46096
rect 32128 46112 32180 46164
rect 34428 46155 34480 46164
rect 21916 46019 21968 46028
rect 21916 45985 21925 46019
rect 21925 45985 21959 46019
rect 21959 45985 21968 46019
rect 21916 45976 21968 45985
rect 22192 45976 22244 46028
rect 23940 46019 23992 46028
rect 23940 45985 23949 46019
rect 23949 45985 23983 46019
rect 23983 45985 23992 46019
rect 24492 46019 24544 46028
rect 23940 45976 23992 45985
rect 24492 45985 24501 46019
rect 24501 45985 24535 46019
rect 24535 45985 24544 46019
rect 24492 45976 24544 45985
rect 24676 46019 24728 46028
rect 24676 45985 24685 46019
rect 24685 45985 24719 46019
rect 24719 45985 24728 46019
rect 24676 45976 24728 45985
rect 27068 46019 27120 46028
rect 27068 45985 27077 46019
rect 27077 45985 27111 46019
rect 27111 45985 27120 46019
rect 27068 45976 27120 45985
rect 27804 45976 27856 46028
rect 29092 46019 29144 46028
rect 29092 45985 29101 46019
rect 29101 45985 29135 46019
rect 29135 45985 29144 46019
rect 29092 45976 29144 45985
rect 32036 46044 32088 46096
rect 34428 46121 34437 46155
rect 34437 46121 34471 46155
rect 34471 46121 34480 46155
rect 34428 46112 34480 46121
rect 39212 46155 39264 46164
rect 32312 45976 32364 46028
rect 38476 46019 38528 46028
rect 38476 45985 38485 46019
rect 38485 45985 38519 46019
rect 38519 45985 38528 46019
rect 38476 45976 38528 45985
rect 39212 46121 39221 46155
rect 39221 46121 39255 46155
rect 39255 46121 39264 46155
rect 39212 46112 39264 46121
rect 46112 46112 46164 46164
rect 46940 46112 46992 46164
rect 57428 46112 57480 46164
rect 40776 46044 40828 46096
rect 44364 46087 44416 46096
rect 44364 46053 44373 46087
rect 44373 46053 44407 46087
rect 44407 46053 44416 46087
rect 44364 46044 44416 46053
rect 45008 46019 45060 46028
rect 45008 45985 45017 46019
rect 45017 45985 45051 46019
rect 45051 45985 45060 46019
rect 45008 45976 45060 45985
rect 45376 46019 45428 46028
rect 45376 45985 45385 46019
rect 45385 45985 45419 46019
rect 45419 45985 45428 46019
rect 45376 45976 45428 45985
rect 47308 46044 47360 46096
rect 46664 46019 46716 46028
rect 46664 45985 46673 46019
rect 46673 45985 46707 46019
rect 46707 45985 46716 46019
rect 46664 45976 46716 45985
rect 16764 45840 16816 45849
rect 24952 45908 25004 45960
rect 24492 45840 24544 45892
rect 29184 45840 29236 45892
rect 22192 45772 22244 45824
rect 24676 45772 24728 45824
rect 27160 45815 27212 45824
rect 27160 45781 27169 45815
rect 27169 45781 27203 45815
rect 27203 45781 27212 45815
rect 27160 45772 27212 45781
rect 32588 45908 32640 45960
rect 35440 45908 35492 45960
rect 34980 45840 35032 45892
rect 30380 45772 30432 45824
rect 40132 45840 40184 45892
rect 45928 45908 45980 45960
rect 48688 45908 48740 45960
rect 51172 46019 51224 46028
rect 51172 45985 51181 46019
rect 51181 45985 51215 46019
rect 51215 45985 51224 46019
rect 51172 45976 51224 45985
rect 51632 45976 51684 46028
rect 51724 46019 51776 46028
rect 51724 45985 51733 46019
rect 51733 45985 51767 46019
rect 51767 45985 51776 46019
rect 54852 46044 54904 46096
rect 56784 46044 56836 46096
rect 61476 46044 61528 46096
rect 51724 45976 51776 45985
rect 55956 45976 56008 46028
rect 63224 45976 63276 46028
rect 62304 45951 62356 45960
rect 62304 45917 62313 45951
rect 62313 45917 62347 45951
rect 62347 45917 62356 45951
rect 62304 45908 62356 45917
rect 62028 45840 62080 45892
rect 45928 45815 45980 45824
rect 45928 45781 45937 45815
rect 45937 45781 45971 45815
rect 45971 45781 45980 45815
rect 45928 45772 45980 45781
rect 46480 45772 46532 45824
rect 47308 45815 47360 45824
rect 47308 45781 47317 45815
rect 47317 45781 47351 45815
rect 47351 45781 47360 45815
rect 47308 45772 47360 45781
rect 52644 45772 52696 45824
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 65686 45670 65738 45722
rect 65750 45670 65802 45722
rect 65814 45670 65866 45722
rect 65878 45670 65930 45722
rect 96406 45670 96458 45722
rect 96470 45670 96522 45722
rect 96534 45670 96586 45722
rect 96598 45670 96650 45722
rect 27160 45568 27212 45620
rect 38568 45568 38620 45620
rect 46664 45568 46716 45620
rect 54484 45568 54536 45620
rect 55128 45568 55180 45620
rect 15660 45500 15712 45552
rect 44548 45500 44600 45552
rect 47676 45500 47728 45552
rect 65064 45500 65116 45552
rect 4620 45432 4672 45484
rect 13452 45475 13504 45484
rect 13452 45441 13461 45475
rect 13461 45441 13495 45475
rect 13495 45441 13504 45475
rect 13452 45432 13504 45441
rect 15476 45432 15528 45484
rect 30840 45432 30892 45484
rect 32864 45432 32916 45484
rect 2596 45407 2648 45416
rect 2596 45373 2605 45407
rect 2605 45373 2639 45407
rect 2639 45373 2648 45407
rect 2596 45364 2648 45373
rect 13820 45364 13872 45416
rect 23388 45364 23440 45416
rect 31852 45364 31904 45416
rect 44456 45407 44508 45416
rect 30380 45296 30432 45348
rect 2964 45228 3016 45280
rect 4436 45271 4488 45280
rect 4436 45237 4445 45271
rect 4445 45237 4479 45271
rect 4479 45237 4488 45271
rect 4436 45228 4488 45237
rect 30840 45271 30892 45280
rect 30840 45237 30849 45271
rect 30849 45237 30883 45271
rect 30883 45237 30892 45271
rect 30840 45228 30892 45237
rect 44456 45373 44465 45407
rect 44465 45373 44499 45407
rect 44499 45373 44508 45407
rect 44456 45364 44508 45373
rect 46112 45407 46164 45416
rect 46112 45373 46121 45407
rect 46121 45373 46155 45407
rect 46155 45373 46164 45407
rect 46112 45364 46164 45373
rect 51908 45407 51960 45416
rect 51908 45373 51917 45407
rect 51917 45373 51951 45407
rect 51951 45373 51960 45407
rect 51908 45364 51960 45373
rect 33876 45228 33928 45280
rect 52460 45407 52512 45416
rect 52460 45373 52469 45407
rect 52469 45373 52503 45407
rect 52503 45373 52512 45407
rect 52460 45364 52512 45373
rect 56600 45364 56652 45416
rect 58532 45364 58584 45416
rect 54944 45296 54996 45348
rect 55864 45296 55916 45348
rect 65248 45296 65300 45348
rect 43812 45228 43864 45280
rect 45376 45228 45428 45280
rect 51908 45228 51960 45280
rect 55956 45228 56008 45280
rect 56600 45228 56652 45280
rect 57520 45228 57572 45280
rect 57704 45228 57756 45280
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 50326 45126 50378 45178
rect 50390 45126 50442 45178
rect 50454 45126 50506 45178
rect 50518 45126 50570 45178
rect 81046 45126 81098 45178
rect 81110 45126 81162 45178
rect 81174 45126 81226 45178
rect 81238 45126 81290 45178
rect 4436 45024 4488 45076
rect 4712 45024 4764 45076
rect 7196 45067 7248 45076
rect 7196 45033 7205 45067
rect 7205 45033 7239 45067
rect 7239 45033 7248 45067
rect 7196 45024 7248 45033
rect 15292 45024 15344 45076
rect 6920 44820 6972 44872
rect 23388 45024 23440 45076
rect 29184 45067 29236 45076
rect 29184 45033 29193 45067
rect 29193 45033 29227 45067
rect 29227 45033 29236 45067
rect 29184 45024 29236 45033
rect 44548 45067 44600 45076
rect 44548 45033 44557 45067
rect 44557 45033 44591 45067
rect 44591 45033 44600 45067
rect 44548 45024 44600 45033
rect 44732 45067 44784 45076
rect 44732 45033 44741 45067
rect 44741 45033 44775 45067
rect 44775 45033 44784 45067
rect 44732 45024 44784 45033
rect 45468 45024 45520 45076
rect 47308 45024 47360 45076
rect 60924 45024 60976 45076
rect 62304 45024 62356 45076
rect 44456 44956 44508 45008
rect 23848 44888 23900 44940
rect 29184 44888 29236 44940
rect 44364 44888 44416 44940
rect 44548 44888 44600 44940
rect 45468 44931 45520 44940
rect 38752 44820 38804 44872
rect 39212 44863 39264 44872
rect 39212 44829 39221 44863
rect 39221 44829 39255 44863
rect 39255 44829 39264 44863
rect 39212 44820 39264 44829
rect 45468 44897 45477 44931
rect 45477 44897 45511 44931
rect 45511 44897 45520 44931
rect 45468 44888 45520 44897
rect 61568 44956 61620 45008
rect 46848 44888 46900 44940
rect 46572 44820 46624 44872
rect 55864 44888 55916 44940
rect 57704 44931 57756 44940
rect 57704 44897 57713 44931
rect 57713 44897 57747 44931
rect 57747 44897 57756 44931
rect 57704 44888 57756 44897
rect 60372 44931 60424 44940
rect 60372 44897 60381 44931
rect 60381 44897 60415 44931
rect 60415 44897 60424 44931
rect 60372 44888 60424 44897
rect 61752 44931 61804 44940
rect 61752 44897 61761 44931
rect 61761 44897 61795 44931
rect 61795 44897 61804 44931
rect 61752 44888 61804 44897
rect 65524 44956 65576 45008
rect 52644 44863 52696 44872
rect 46480 44752 46532 44804
rect 47124 44752 47176 44804
rect 51724 44752 51776 44804
rect 52644 44829 52653 44863
rect 52653 44829 52687 44863
rect 52687 44829 52696 44863
rect 52644 44820 52696 44829
rect 57336 44820 57388 44872
rect 59176 44820 59228 44872
rect 57244 44752 57296 44804
rect 60740 44820 60792 44872
rect 62028 44820 62080 44872
rect 63224 44863 63276 44872
rect 63224 44829 63233 44863
rect 63233 44829 63267 44863
rect 63267 44829 63276 44863
rect 63224 44820 63276 44829
rect 64328 44820 64380 44872
rect 66904 44820 66956 44872
rect 62948 44752 63000 44804
rect 7012 44684 7064 44736
rect 23848 44684 23900 44736
rect 38752 44727 38804 44736
rect 38752 44693 38761 44727
rect 38761 44693 38795 44727
rect 38795 44693 38804 44727
rect 38752 44684 38804 44693
rect 40500 44727 40552 44736
rect 40500 44693 40509 44727
rect 40509 44693 40543 44727
rect 40543 44693 40552 44727
rect 40500 44684 40552 44693
rect 52460 44727 52512 44736
rect 52460 44693 52484 44727
rect 52484 44693 52512 44727
rect 52460 44684 52512 44693
rect 52552 44727 52604 44736
rect 52552 44693 52561 44727
rect 52561 44693 52595 44727
rect 52595 44693 52604 44727
rect 52552 44684 52604 44693
rect 54576 44684 54628 44736
rect 59084 44684 59136 44736
rect 60464 44727 60516 44736
rect 60464 44693 60473 44727
rect 60473 44693 60507 44727
rect 60507 44693 60516 44727
rect 60464 44684 60516 44693
rect 68560 44684 68612 44736
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 65686 44582 65738 44634
rect 65750 44582 65802 44634
rect 65814 44582 65866 44634
rect 65878 44582 65930 44634
rect 96406 44582 96458 44634
rect 96470 44582 96522 44634
rect 96534 44582 96586 44634
rect 96598 44582 96650 44634
rect 4712 44480 4764 44532
rect 7840 44480 7892 44532
rect 39212 44480 39264 44532
rect 15292 44455 15344 44464
rect 15292 44421 15301 44455
rect 15301 44421 15335 44455
rect 15335 44421 15344 44455
rect 15292 44412 15344 44421
rect 15476 44455 15528 44464
rect 15476 44421 15485 44455
rect 15485 44421 15519 44455
rect 15519 44421 15528 44455
rect 15476 44412 15528 44421
rect 2596 44319 2648 44328
rect 2596 44285 2605 44319
rect 2605 44285 2639 44319
rect 2639 44285 2648 44319
rect 2596 44276 2648 44285
rect 6736 44276 6788 44328
rect 2872 44140 2924 44192
rect 4620 44140 4672 44192
rect 8944 44276 8996 44328
rect 9036 44276 9088 44328
rect 24768 44344 24820 44396
rect 13452 44276 13504 44328
rect 14004 44319 14056 44328
rect 14004 44285 14013 44319
rect 14013 44285 14047 44319
rect 14047 44285 14056 44319
rect 14004 44276 14056 44285
rect 18972 44319 19024 44328
rect 9680 44208 9732 44260
rect 18972 44285 18981 44319
rect 18981 44285 19015 44319
rect 19015 44285 19024 44319
rect 18972 44276 19024 44285
rect 22652 44276 22704 44328
rect 27804 44319 27856 44328
rect 27804 44285 27813 44319
rect 27813 44285 27847 44319
rect 27847 44285 27856 44319
rect 27804 44276 27856 44285
rect 20904 44208 20956 44260
rect 21088 44208 21140 44260
rect 21916 44208 21968 44260
rect 28264 44208 28316 44260
rect 29000 44208 29052 44260
rect 31944 44344 31996 44396
rect 56784 44480 56836 44532
rect 58532 44523 58584 44532
rect 58532 44489 58541 44523
rect 58541 44489 58575 44523
rect 58575 44489 58584 44523
rect 58532 44480 58584 44489
rect 60464 44480 60516 44532
rect 60740 44523 60792 44532
rect 60740 44489 60749 44523
rect 60749 44489 60783 44523
rect 60783 44489 60792 44523
rect 60924 44523 60976 44532
rect 60740 44480 60792 44489
rect 60924 44489 60933 44523
rect 60933 44489 60967 44523
rect 60967 44489 60976 44523
rect 60924 44480 60976 44489
rect 65248 44523 65300 44532
rect 65248 44489 65257 44523
rect 65257 44489 65291 44523
rect 65291 44489 65300 44523
rect 65984 44523 66036 44532
rect 65248 44480 65300 44489
rect 65984 44489 65993 44523
rect 65993 44489 66027 44523
rect 66027 44489 66036 44523
rect 65984 44480 66036 44489
rect 71320 44480 71372 44532
rect 73620 44480 73672 44532
rect 44364 44412 44416 44464
rect 45468 44412 45520 44464
rect 47676 44455 47728 44464
rect 31852 44276 31904 44328
rect 32864 44276 32916 44328
rect 40500 44276 40552 44328
rect 47676 44421 47685 44455
rect 47685 44421 47719 44455
rect 47719 44421 47728 44455
rect 47676 44412 47728 44421
rect 51724 44387 51776 44396
rect 51724 44353 51733 44387
rect 51733 44353 51767 44387
rect 51767 44353 51776 44387
rect 51724 44344 51776 44353
rect 46848 44319 46900 44328
rect 46848 44285 46857 44319
rect 46857 44285 46891 44319
rect 46891 44285 46900 44319
rect 46848 44276 46900 44285
rect 51264 44276 51316 44328
rect 51908 44319 51960 44328
rect 51908 44285 51917 44319
rect 51917 44285 51951 44319
rect 51951 44285 51960 44319
rect 51908 44276 51960 44285
rect 21824 44140 21876 44192
rect 52828 44412 52880 44464
rect 57244 44344 57296 44396
rect 66076 44412 66128 44464
rect 66168 44412 66220 44464
rect 71412 44412 71464 44464
rect 60740 44344 60792 44396
rect 65984 44344 66036 44396
rect 29092 44140 29144 44192
rect 45560 44183 45612 44192
rect 45560 44149 45569 44183
rect 45569 44149 45603 44183
rect 45603 44149 45612 44183
rect 45560 44140 45612 44149
rect 47124 44140 47176 44192
rect 50712 44140 50764 44192
rect 59176 44276 59228 44328
rect 59452 44319 59504 44328
rect 59452 44285 59461 44319
rect 59461 44285 59495 44319
rect 59495 44285 59504 44319
rect 59452 44276 59504 44285
rect 65064 44319 65116 44328
rect 65064 44285 65073 44319
rect 65073 44285 65107 44319
rect 65107 44285 65116 44319
rect 65064 44276 65116 44285
rect 54668 44208 54720 44260
rect 60188 44208 60240 44260
rect 65524 44276 65576 44328
rect 66996 44319 67048 44328
rect 66996 44285 67005 44319
rect 67005 44285 67039 44319
rect 67039 44285 67048 44319
rect 66996 44276 67048 44285
rect 68560 44319 68612 44328
rect 68560 44285 68569 44319
rect 68569 44285 68603 44319
rect 68603 44285 68612 44319
rect 68560 44276 68612 44285
rect 53288 44183 53340 44192
rect 53288 44149 53297 44183
rect 53297 44149 53331 44183
rect 53331 44149 53340 44183
rect 53288 44140 53340 44149
rect 66168 44140 66220 44192
rect 68744 44140 68796 44192
rect 71320 44140 71372 44192
rect 72884 44276 72936 44328
rect 77392 44208 77444 44260
rect 72976 44183 73028 44192
rect 72976 44149 72985 44183
rect 72985 44149 73019 44183
rect 73019 44149 73028 44183
rect 72976 44140 73028 44149
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 81046 44038 81098 44090
rect 81110 44038 81162 44090
rect 81174 44038 81226 44090
rect 81238 44038 81290 44090
rect 6920 43979 6972 43988
rect 6920 43945 6929 43979
rect 6929 43945 6963 43979
rect 6963 43945 6972 43979
rect 6920 43936 6972 43945
rect 7104 43800 7156 43852
rect 7840 43936 7892 43988
rect 13820 43936 13872 43988
rect 15660 43979 15712 43988
rect 15660 43945 15669 43979
rect 15669 43945 15703 43979
rect 15703 43945 15712 43979
rect 15660 43936 15712 43945
rect 17224 43936 17276 43988
rect 31944 43979 31996 43988
rect 31944 43945 31953 43979
rect 31953 43945 31987 43979
rect 31987 43945 31996 43979
rect 31944 43936 31996 43945
rect 9680 43843 9732 43852
rect 9680 43809 9689 43843
rect 9689 43809 9723 43843
rect 9723 43809 9732 43843
rect 9680 43800 9732 43809
rect 14280 43868 14332 43920
rect 3700 43664 3752 43716
rect 12716 43707 12768 43716
rect 12716 43673 12725 43707
rect 12725 43673 12759 43707
rect 12759 43673 12768 43707
rect 12716 43664 12768 43673
rect 12900 43664 12952 43716
rect 20904 43843 20956 43852
rect 17132 43732 17184 43784
rect 20904 43809 20913 43843
rect 20913 43809 20947 43843
rect 20947 43809 20956 43843
rect 20904 43800 20956 43809
rect 29184 43868 29236 43920
rect 27804 43800 27856 43852
rect 28264 43843 28316 43852
rect 28264 43809 28273 43843
rect 28273 43809 28307 43843
rect 28307 43809 28316 43843
rect 28264 43800 28316 43809
rect 28632 43800 28684 43852
rect 32036 43868 32088 43920
rect 32956 43936 33008 43988
rect 34244 43936 34296 43988
rect 45560 43936 45612 43988
rect 45836 43936 45888 43988
rect 46572 43979 46624 43988
rect 46572 43945 46581 43979
rect 46581 43945 46615 43979
rect 46615 43945 46624 43979
rect 46572 43936 46624 43945
rect 54116 43936 54168 43988
rect 59452 43936 59504 43988
rect 60372 43936 60424 43988
rect 60464 43936 60516 43988
rect 72884 43979 72936 43988
rect 22192 43775 22244 43784
rect 9772 43639 9824 43648
rect 9772 43605 9781 43639
rect 9781 43605 9815 43639
rect 9815 43605 9824 43639
rect 9772 43596 9824 43605
rect 22192 43741 22201 43775
rect 22201 43741 22235 43775
rect 22235 43741 22244 43775
rect 22192 43732 22244 43741
rect 29000 43732 29052 43784
rect 32956 43843 33008 43852
rect 32956 43809 32965 43843
rect 32965 43809 32999 43843
rect 32999 43809 33008 43843
rect 32956 43800 33008 43809
rect 36360 43800 36412 43852
rect 38476 43843 38528 43852
rect 38476 43809 38485 43843
rect 38485 43809 38519 43843
rect 38519 43809 38528 43843
rect 38476 43800 38528 43809
rect 44548 43800 44600 43852
rect 45284 43843 45336 43852
rect 39488 43732 39540 43784
rect 20352 43596 20404 43648
rect 20996 43639 21048 43648
rect 20996 43605 21005 43639
rect 21005 43605 21039 43639
rect 21039 43605 21048 43639
rect 20996 43596 21048 43605
rect 21916 43596 21968 43648
rect 23388 43596 23440 43648
rect 23664 43596 23716 43648
rect 28632 43639 28684 43648
rect 28632 43605 28641 43639
rect 28641 43605 28675 43639
rect 28675 43605 28684 43639
rect 28632 43596 28684 43605
rect 45284 43809 45293 43843
rect 45293 43809 45327 43843
rect 45327 43809 45336 43843
rect 45284 43800 45336 43809
rect 45836 43843 45888 43852
rect 45836 43809 45845 43843
rect 45845 43809 45879 43843
rect 45879 43809 45888 43843
rect 45836 43800 45888 43809
rect 45100 43775 45152 43784
rect 45100 43741 45109 43775
rect 45109 43741 45143 43775
rect 45143 43741 45152 43775
rect 45100 43732 45152 43741
rect 51264 43843 51316 43852
rect 51264 43809 51273 43843
rect 51273 43809 51307 43843
rect 51307 43809 51316 43843
rect 51264 43800 51316 43809
rect 51908 43800 51960 43852
rect 52460 43868 52512 43920
rect 52828 43868 52880 43920
rect 34244 43596 34296 43648
rect 35440 43596 35492 43648
rect 37188 43596 37240 43648
rect 38752 43596 38804 43648
rect 39488 43639 39540 43648
rect 39488 43605 39497 43639
rect 39497 43605 39531 43639
rect 39531 43605 39540 43639
rect 39488 43596 39540 43605
rect 52460 43664 52512 43716
rect 54668 43800 54720 43852
rect 59084 43868 59136 43920
rect 60188 43843 60240 43852
rect 60188 43809 60197 43843
rect 60197 43809 60231 43843
rect 60231 43809 60240 43843
rect 60188 43800 60240 43809
rect 60740 43868 60792 43920
rect 65984 43911 66036 43920
rect 60556 43800 60608 43852
rect 65984 43877 65993 43911
rect 65993 43877 66027 43911
rect 66027 43877 66036 43911
rect 65984 43868 66036 43877
rect 66904 43868 66956 43920
rect 72516 43868 72568 43920
rect 54944 43775 54996 43784
rect 54944 43741 54953 43775
rect 54953 43741 54987 43775
rect 54987 43741 54996 43775
rect 54944 43732 54996 43741
rect 66260 43800 66312 43852
rect 66996 43843 67048 43852
rect 66996 43809 67005 43843
rect 67005 43809 67039 43843
rect 67039 43809 67048 43843
rect 66996 43800 67048 43809
rect 71596 43843 71648 43852
rect 71596 43809 71605 43843
rect 71605 43809 71639 43843
rect 71639 43809 71648 43843
rect 71596 43800 71648 43809
rect 71780 43732 71832 43784
rect 72884 43945 72893 43979
rect 72893 43945 72927 43979
rect 72927 43945 72936 43979
rect 72884 43936 72936 43945
rect 77392 43979 77444 43988
rect 77392 43945 77401 43979
rect 77401 43945 77435 43979
rect 77435 43945 77444 43979
rect 77392 43936 77444 43945
rect 72792 43843 72844 43852
rect 72792 43809 72801 43843
rect 72801 43809 72835 43843
rect 72835 43809 72844 43843
rect 72792 43800 72844 43809
rect 79600 43800 79652 43852
rect 77760 43732 77812 43784
rect 53288 43664 53340 43716
rect 42248 43639 42300 43648
rect 42248 43605 42257 43639
rect 42257 43605 42291 43639
rect 42291 43605 42300 43639
rect 42248 43596 42300 43605
rect 44548 43596 44600 43648
rect 45100 43596 45152 43648
rect 46756 43639 46808 43648
rect 46756 43605 46765 43639
rect 46765 43605 46799 43639
rect 46799 43605 46808 43639
rect 46756 43596 46808 43605
rect 52920 43596 52972 43648
rect 60004 43664 60056 43716
rect 60280 43596 60332 43648
rect 60464 43639 60516 43648
rect 60464 43605 60473 43639
rect 60473 43605 60507 43639
rect 60507 43605 60516 43639
rect 60464 43596 60516 43605
rect 63224 43664 63276 43716
rect 79692 43596 79744 43648
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 65686 43494 65738 43546
rect 65750 43494 65802 43546
rect 65814 43494 65866 43546
rect 65878 43494 65930 43546
rect 96406 43494 96458 43546
rect 96470 43494 96522 43546
rect 96534 43494 96586 43546
rect 96598 43494 96650 43546
rect 3976 43435 4028 43444
rect 3976 43401 3985 43435
rect 3985 43401 4019 43435
rect 4019 43401 4028 43435
rect 3976 43392 4028 43401
rect 11612 43392 11664 43444
rect 12716 43435 12768 43444
rect 12716 43401 12725 43435
rect 12725 43401 12759 43435
rect 12759 43401 12768 43435
rect 14004 43435 14056 43444
rect 12716 43392 12768 43401
rect 4712 43324 4764 43376
rect 2596 43231 2648 43240
rect 2596 43197 2605 43231
rect 2605 43197 2639 43231
rect 2639 43197 2648 43231
rect 2596 43188 2648 43197
rect 8668 43324 8720 43376
rect 8944 43367 8996 43376
rect 8944 43333 8953 43367
rect 8953 43333 8987 43367
rect 8987 43333 8996 43367
rect 8944 43324 8996 43333
rect 14004 43401 14013 43435
rect 14013 43401 14047 43435
rect 14047 43401 14056 43435
rect 14004 43392 14056 43401
rect 15292 43435 15344 43444
rect 15292 43401 15301 43435
rect 15301 43401 15335 43435
rect 15335 43401 15344 43435
rect 15292 43392 15344 43401
rect 16580 43256 16632 43308
rect 4712 43052 4764 43104
rect 7564 43052 7616 43104
rect 8668 43188 8720 43240
rect 8944 43188 8996 43240
rect 12900 43188 12952 43240
rect 9772 43052 9824 43104
rect 10140 43052 10192 43104
rect 13636 43120 13688 43172
rect 15292 43188 15344 43240
rect 16580 43120 16632 43172
rect 18972 43324 19024 43376
rect 22192 43392 22244 43444
rect 22652 43435 22704 43444
rect 22652 43401 22661 43435
rect 22661 43401 22695 43435
rect 22695 43401 22704 43435
rect 22652 43392 22704 43401
rect 23388 43392 23440 43444
rect 19892 43324 19944 43376
rect 20996 43324 21048 43376
rect 24768 43367 24820 43376
rect 20260 43188 20312 43240
rect 20352 43188 20404 43240
rect 24124 43256 24176 43308
rect 22468 43231 22520 43240
rect 22468 43197 22477 43231
rect 22477 43197 22511 43231
rect 22511 43197 22520 43231
rect 22468 43188 22520 43197
rect 23664 43231 23716 43240
rect 23664 43197 23673 43231
rect 23673 43197 23707 43231
rect 23707 43197 23716 43231
rect 23664 43188 23716 43197
rect 20812 43120 20864 43172
rect 24768 43333 24777 43367
rect 24777 43333 24811 43367
rect 24811 43333 24820 43367
rect 24768 43324 24820 43333
rect 28632 43392 28684 43444
rect 33324 43392 33376 43444
rect 38384 43392 38436 43444
rect 52920 43435 52972 43444
rect 52920 43401 52929 43435
rect 52929 43401 52963 43435
rect 52963 43401 52972 43435
rect 52920 43392 52972 43401
rect 53196 43392 53248 43444
rect 59084 43392 59136 43444
rect 59544 43392 59596 43444
rect 37188 43367 37240 43376
rect 37188 43333 37197 43367
rect 37197 43333 37231 43367
rect 37231 43333 37240 43367
rect 37188 43324 37240 43333
rect 32772 43256 32824 43308
rect 35440 43299 35492 43308
rect 35440 43265 35449 43299
rect 35449 43265 35483 43299
rect 35483 43265 35492 43299
rect 35440 43256 35492 43265
rect 26240 43231 26292 43240
rect 26240 43197 26249 43231
rect 26249 43197 26283 43231
rect 26283 43197 26292 43231
rect 26240 43188 26292 43197
rect 32956 43188 33008 43240
rect 33324 43231 33376 43240
rect 33324 43197 33333 43231
rect 33333 43197 33367 43231
rect 33367 43197 33376 43231
rect 33324 43188 33376 43197
rect 35716 43231 35768 43240
rect 35716 43197 35725 43231
rect 35725 43197 35759 43231
rect 35759 43197 35768 43231
rect 35716 43188 35768 43197
rect 42248 43324 42300 43376
rect 56600 43324 56652 43376
rect 60188 43324 60240 43376
rect 37832 43256 37884 43308
rect 44824 43256 44876 43308
rect 53012 43256 53064 43308
rect 58716 43256 58768 43308
rect 17776 43095 17828 43104
rect 17776 43061 17785 43095
rect 17785 43061 17819 43095
rect 17819 43061 17828 43095
rect 17776 43052 17828 43061
rect 17868 43052 17920 43104
rect 22468 43052 22520 43104
rect 23756 43095 23808 43104
rect 23756 43061 23765 43095
rect 23765 43061 23799 43095
rect 23799 43061 23808 43095
rect 23756 43052 23808 43061
rect 25044 43095 25096 43104
rect 25044 43061 25053 43095
rect 25053 43061 25087 43095
rect 25087 43061 25096 43095
rect 25044 43052 25096 43061
rect 27528 43095 27580 43104
rect 27528 43061 27537 43095
rect 27537 43061 27571 43095
rect 27571 43061 27580 43095
rect 27528 43052 27580 43061
rect 32312 43095 32364 43104
rect 32312 43061 32321 43095
rect 32321 43061 32355 43095
rect 32355 43061 32364 43095
rect 32312 43052 32364 43061
rect 51448 43188 51500 43240
rect 52000 43188 52052 43240
rect 33968 43095 34020 43104
rect 33968 43061 33977 43095
rect 33977 43061 34011 43095
rect 34011 43061 34020 43095
rect 33968 43052 34020 43061
rect 44824 43120 44876 43172
rect 53196 43188 53248 43240
rect 60464 43256 60516 43308
rect 71044 43324 71096 43376
rect 72976 43367 73028 43376
rect 59452 43188 59504 43240
rect 60096 43231 60148 43240
rect 39488 43095 39540 43104
rect 39488 43061 39497 43095
rect 39497 43061 39531 43095
rect 39531 43061 39540 43095
rect 39488 43052 39540 43061
rect 51448 43095 51500 43104
rect 51448 43061 51457 43095
rect 51457 43061 51491 43095
rect 51491 43061 51500 43095
rect 51448 43052 51500 43061
rect 59176 43052 59228 43104
rect 59636 43052 59688 43104
rect 60096 43197 60105 43231
rect 60105 43197 60139 43231
rect 60139 43197 60148 43231
rect 60096 43188 60148 43197
rect 61568 43231 61620 43240
rect 61568 43197 61577 43231
rect 61577 43197 61611 43231
rect 61611 43197 61620 43231
rect 61568 43188 61620 43197
rect 66904 43231 66956 43240
rect 66904 43197 66913 43231
rect 66913 43197 66947 43231
rect 66947 43197 66956 43231
rect 66904 43188 66956 43197
rect 67088 43188 67140 43240
rect 71044 43188 71096 43240
rect 60004 43163 60056 43172
rect 60004 43129 60013 43163
rect 60013 43129 60047 43163
rect 60047 43129 60056 43163
rect 60004 43120 60056 43129
rect 60188 43120 60240 43172
rect 60556 43120 60608 43172
rect 66720 43163 66772 43172
rect 60648 43095 60700 43104
rect 60648 43061 60657 43095
rect 60657 43061 60691 43095
rect 60691 43061 60700 43095
rect 60648 43052 60700 43061
rect 66720 43129 66729 43163
rect 66729 43129 66763 43163
rect 66763 43129 66772 43163
rect 66720 43120 66772 43129
rect 71228 43231 71280 43240
rect 71228 43197 71237 43231
rect 71237 43197 71271 43231
rect 71271 43197 71280 43231
rect 71228 43188 71280 43197
rect 71872 43188 71924 43240
rect 72976 43333 72985 43367
rect 72985 43333 73019 43367
rect 73019 43333 73028 43367
rect 72976 43324 73028 43333
rect 77760 43256 77812 43308
rect 77852 43188 77904 43240
rect 78404 43231 78456 43240
rect 78404 43197 78413 43231
rect 78413 43197 78447 43231
rect 78447 43197 78456 43231
rect 78404 43188 78456 43197
rect 78588 43231 78640 43240
rect 78588 43197 78597 43231
rect 78597 43197 78631 43231
rect 78631 43197 78640 43231
rect 78588 43188 78640 43197
rect 71964 43163 72016 43172
rect 71964 43129 71973 43163
rect 71973 43129 72007 43163
rect 72007 43129 72016 43163
rect 71964 43120 72016 43129
rect 66352 43052 66404 43104
rect 66996 43095 67048 43104
rect 66996 43061 67005 43095
rect 67005 43061 67039 43095
rect 67039 43061 67048 43095
rect 66996 43052 67048 43061
rect 72424 43052 72476 43104
rect 77484 43095 77536 43104
rect 77484 43061 77493 43095
rect 77493 43061 77527 43095
rect 77527 43061 77536 43095
rect 77484 43052 77536 43061
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 81046 42950 81098 43002
rect 81110 42950 81162 43002
rect 81174 42950 81226 43002
rect 81238 42950 81290 43002
rect 4068 42848 4120 42900
rect 32312 42848 32364 42900
rect 33968 42848 34020 42900
rect 44732 42848 44784 42900
rect 44824 42891 44876 42900
rect 44824 42857 44833 42891
rect 44833 42857 44867 42891
rect 44867 42857 44876 42891
rect 46572 42891 46624 42900
rect 44824 42848 44876 42857
rect 46572 42857 46581 42891
rect 46581 42857 46615 42891
rect 46615 42857 46624 42891
rect 46572 42848 46624 42857
rect 51264 42848 51316 42900
rect 51816 42848 51868 42900
rect 52000 42848 52052 42900
rect 53012 42891 53064 42900
rect 53012 42857 53021 42891
rect 53021 42857 53055 42891
rect 53055 42857 53064 42891
rect 53012 42848 53064 42857
rect 53196 42891 53248 42900
rect 53196 42857 53205 42891
rect 53205 42857 53239 42891
rect 53239 42857 53248 42891
rect 53196 42848 53248 42857
rect 77852 42891 77904 42900
rect 77852 42857 77861 42891
rect 77861 42857 77895 42891
rect 77895 42857 77904 42891
rect 77852 42848 77904 42857
rect 6736 42780 6788 42832
rect 7104 42755 7156 42764
rect 7104 42721 7113 42755
rect 7113 42721 7147 42755
rect 7147 42721 7156 42755
rect 7104 42712 7156 42721
rect 17224 42780 17276 42832
rect 23756 42780 23808 42832
rect 44548 42780 44600 42832
rect 13728 42755 13780 42764
rect 13728 42721 13737 42755
rect 13737 42721 13771 42755
rect 13771 42721 13780 42755
rect 13728 42712 13780 42721
rect 14004 42712 14056 42764
rect 14280 42755 14332 42764
rect 14280 42721 14289 42755
rect 14289 42721 14323 42755
rect 14323 42721 14332 42755
rect 14280 42712 14332 42721
rect 16396 42712 16448 42764
rect 29920 42712 29972 42764
rect 32312 42712 32364 42764
rect 32864 42755 32916 42764
rect 32864 42721 32873 42755
rect 32873 42721 32907 42755
rect 32907 42721 32916 42755
rect 32864 42712 32916 42721
rect 34244 42755 34296 42764
rect 34244 42721 34253 42755
rect 34253 42721 34287 42755
rect 34287 42721 34296 42755
rect 34244 42712 34296 42721
rect 39488 42712 39540 42764
rect 44364 42712 44416 42764
rect 45284 42780 45336 42832
rect 45560 42712 45612 42764
rect 46572 42712 46624 42764
rect 46756 42755 46808 42764
rect 46756 42721 46765 42755
rect 46765 42721 46799 42755
rect 46799 42721 46808 42755
rect 46756 42712 46808 42721
rect 11060 42644 11112 42696
rect 13636 42687 13688 42696
rect 13636 42653 13645 42687
rect 13645 42653 13679 42687
rect 13679 42653 13688 42687
rect 13636 42644 13688 42653
rect 35716 42644 35768 42696
rect 4068 42576 4120 42628
rect 30840 42576 30892 42628
rect 44548 42576 44600 42628
rect 51264 42644 51316 42696
rect 51724 42712 51776 42764
rect 52184 42755 52236 42764
rect 52184 42721 52193 42755
rect 52193 42721 52227 42755
rect 52227 42721 52236 42755
rect 66352 42823 66404 42832
rect 52184 42712 52236 42721
rect 58900 42712 58952 42764
rect 66352 42789 66361 42823
rect 66361 42789 66395 42823
rect 66395 42789 66404 42823
rect 66352 42780 66404 42789
rect 59452 42755 59504 42764
rect 59452 42721 59461 42755
rect 59461 42721 59495 42755
rect 59495 42721 59504 42755
rect 59452 42712 59504 42721
rect 60188 42755 60240 42764
rect 60188 42721 60197 42755
rect 60197 42721 60231 42755
rect 60231 42721 60240 42755
rect 60188 42712 60240 42721
rect 21088 42551 21140 42560
rect 21088 42517 21097 42551
rect 21097 42517 21131 42551
rect 21131 42517 21140 42551
rect 21088 42508 21140 42517
rect 32864 42508 32916 42560
rect 51724 42576 51776 42628
rect 52184 42576 52236 42628
rect 52552 42619 52604 42628
rect 52552 42585 52561 42619
rect 52561 42585 52595 42619
rect 52595 42585 52604 42619
rect 52552 42576 52604 42585
rect 51172 42508 51224 42560
rect 52276 42508 52328 42560
rect 58808 42508 58860 42560
rect 60096 42576 60148 42628
rect 66996 42712 67048 42764
rect 68744 42755 68796 42764
rect 68744 42721 68753 42755
rect 68753 42721 68787 42755
rect 68787 42721 68796 42755
rect 68744 42712 68796 42721
rect 71596 42780 71648 42832
rect 71228 42712 71280 42764
rect 72056 42755 72108 42764
rect 72056 42721 72065 42755
rect 72065 42721 72099 42755
rect 72099 42721 72108 42755
rect 72056 42712 72108 42721
rect 77484 42780 77536 42832
rect 72424 42755 72476 42764
rect 72424 42721 72433 42755
rect 72433 42721 72467 42755
rect 72467 42721 72476 42755
rect 72424 42712 72476 42721
rect 72516 42755 72568 42764
rect 72516 42721 72525 42755
rect 72525 42721 72559 42755
rect 72559 42721 72568 42755
rect 78588 42780 78640 42832
rect 72516 42712 72568 42721
rect 71412 42644 71464 42696
rect 73344 42644 73396 42696
rect 73620 42644 73672 42696
rect 67456 42576 67508 42628
rect 72792 42576 72844 42628
rect 60740 42508 60792 42560
rect 66628 42551 66680 42560
rect 66628 42517 66637 42551
rect 66637 42517 66671 42551
rect 66671 42517 66680 42551
rect 66628 42508 66680 42517
rect 66812 42508 66864 42560
rect 69204 42551 69256 42560
rect 69204 42517 69213 42551
rect 69213 42517 69247 42551
rect 69247 42517 69256 42551
rect 69204 42508 69256 42517
rect 77484 42508 77536 42560
rect 79692 42755 79744 42764
rect 79692 42721 79701 42755
rect 79701 42721 79735 42755
rect 79735 42721 79744 42755
rect 79692 42712 79744 42721
rect 78404 42644 78456 42696
rect 77760 42576 77812 42628
rect 82176 42644 82228 42696
rect 79784 42551 79836 42560
rect 79784 42517 79793 42551
rect 79793 42517 79827 42551
rect 79827 42517 79836 42551
rect 79784 42508 79836 42517
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 65686 42406 65738 42458
rect 65750 42406 65802 42458
rect 65814 42406 65866 42458
rect 65878 42406 65930 42458
rect 96406 42406 96458 42458
rect 96470 42406 96522 42458
rect 96534 42406 96586 42458
rect 96598 42406 96650 42458
rect 3976 42347 4028 42356
rect 3976 42313 3985 42347
rect 3985 42313 4019 42347
rect 4019 42313 4028 42347
rect 3976 42304 4028 42313
rect 4620 42347 4672 42356
rect 4620 42313 4629 42347
rect 4629 42313 4663 42347
rect 4663 42313 4672 42347
rect 4620 42304 4672 42313
rect 7104 42304 7156 42356
rect 16672 42304 16724 42356
rect 17868 42304 17920 42356
rect 2596 42211 2648 42220
rect 2596 42177 2605 42211
rect 2605 42177 2639 42211
rect 2639 42177 2648 42211
rect 13728 42236 13780 42288
rect 2596 42168 2648 42177
rect 4804 42100 4856 42152
rect 7288 42100 7340 42152
rect 16672 42100 16724 42152
rect 19156 42100 19208 42152
rect 17408 42032 17460 42084
rect 16212 41964 16264 42016
rect 20812 42304 20864 42356
rect 26240 42304 26292 42356
rect 19892 42236 19944 42288
rect 20260 42168 20312 42220
rect 19340 41964 19392 42016
rect 23756 41964 23808 42016
rect 25136 42143 25188 42152
rect 25136 42109 25145 42143
rect 25145 42109 25179 42143
rect 25179 42109 25188 42143
rect 25136 42100 25188 42109
rect 27528 42304 27580 42356
rect 53012 42304 53064 42356
rect 53472 42304 53524 42356
rect 58900 42304 58952 42356
rect 64328 42347 64380 42356
rect 64328 42313 64337 42347
rect 64337 42313 64371 42347
rect 64371 42313 64380 42347
rect 64328 42304 64380 42313
rect 66996 42347 67048 42356
rect 66996 42313 67005 42347
rect 67005 42313 67039 42347
rect 67039 42313 67048 42347
rect 66996 42304 67048 42313
rect 70492 42304 70544 42356
rect 72056 42304 72108 42356
rect 77852 42304 77904 42356
rect 29184 42236 29236 42288
rect 31208 42236 31260 42288
rect 32036 42236 32088 42288
rect 32128 42236 32180 42288
rect 58164 42236 58216 42288
rect 59268 42236 59320 42288
rect 61108 42236 61160 42288
rect 27344 42168 27396 42220
rect 29000 42168 29052 42220
rect 40132 42168 40184 42220
rect 53012 42168 53064 42220
rect 58808 42168 58860 42220
rect 66628 42168 66680 42220
rect 66720 42168 66772 42220
rect 29644 42032 29696 42084
rect 26516 41964 26568 42016
rect 29276 41964 29328 42016
rect 31208 42100 31260 42152
rect 36268 42100 36320 42152
rect 46296 42143 46348 42152
rect 46296 42109 46305 42143
rect 46305 42109 46339 42143
rect 46339 42109 46348 42143
rect 46296 42100 46348 42109
rect 40040 41964 40092 42016
rect 41236 41964 41288 42016
rect 46756 41964 46808 42016
rect 52276 42100 52328 42152
rect 49516 42032 49568 42084
rect 51448 42032 51500 42084
rect 59268 42100 59320 42152
rect 72516 42168 72568 42220
rect 77576 42211 77628 42220
rect 77576 42177 77585 42211
rect 77585 42177 77619 42211
rect 77619 42177 77628 42211
rect 77576 42168 77628 42177
rect 67456 42143 67508 42152
rect 53012 42075 53064 42084
rect 53012 42041 53021 42075
rect 53021 42041 53055 42075
rect 53055 42041 53064 42075
rect 53012 42032 53064 42041
rect 47676 42007 47728 42016
rect 47676 41973 47685 42007
rect 47685 41973 47719 42007
rect 47719 41973 47728 42007
rect 47676 41964 47728 41973
rect 51172 42007 51224 42016
rect 51172 41973 51181 42007
rect 51181 41973 51215 42007
rect 51215 41973 51224 42007
rect 51172 41964 51224 41973
rect 51264 41964 51316 42016
rect 59636 42032 59688 42084
rect 58440 41964 58492 42016
rect 59728 42007 59780 42016
rect 59728 41973 59737 42007
rect 59737 41973 59771 42007
rect 59771 41973 59780 42007
rect 67456 42109 67465 42143
rect 67465 42109 67499 42143
rect 67499 42109 67508 42143
rect 67456 42100 67508 42109
rect 66076 42032 66128 42084
rect 69204 42100 69256 42152
rect 65984 42007 66036 42016
rect 59728 41964 59780 41973
rect 65984 41973 65993 42007
rect 65993 41973 66027 42007
rect 66027 41973 66036 42007
rect 65984 41964 66036 41973
rect 66444 41964 66496 42016
rect 66904 41964 66956 42016
rect 67456 41964 67508 42016
rect 71964 42100 72016 42152
rect 77668 42100 77720 42152
rect 71872 42075 71924 42084
rect 71872 42041 71881 42075
rect 71881 42041 71915 42075
rect 71915 42041 71924 42075
rect 71872 42032 71924 42041
rect 72700 42032 72752 42084
rect 77760 42075 77812 42084
rect 77760 42041 77769 42075
rect 77769 42041 77803 42075
rect 77803 42041 77812 42075
rect 77760 42032 77812 42041
rect 71780 41964 71832 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 81046 41862 81098 41914
rect 81110 41862 81162 41914
rect 81174 41862 81226 41914
rect 81238 41862 81290 41914
rect 4620 41760 4672 41812
rect 11152 41692 11204 41744
rect 7288 41624 7340 41676
rect 13452 41760 13504 41812
rect 14004 41760 14056 41812
rect 16212 41760 16264 41812
rect 16396 41803 16448 41812
rect 16396 41769 16405 41803
rect 16405 41769 16439 41803
rect 16439 41769 16448 41803
rect 16396 41760 16448 41769
rect 19432 41760 19484 41812
rect 25136 41760 25188 41812
rect 16120 41624 16172 41676
rect 16396 41624 16448 41676
rect 26516 41667 26568 41676
rect 26516 41633 26525 41667
rect 26525 41633 26559 41667
rect 26559 41633 26568 41667
rect 26516 41624 26568 41633
rect 27344 41760 27396 41812
rect 29644 41803 29696 41812
rect 29644 41769 29653 41803
rect 29653 41769 29687 41803
rect 29687 41769 29696 41803
rect 29644 41760 29696 41769
rect 29920 41803 29972 41812
rect 29920 41769 29929 41803
rect 29929 41769 29963 41803
rect 29963 41769 29972 41803
rect 29920 41760 29972 41769
rect 51264 41760 51316 41812
rect 53472 41803 53524 41812
rect 53472 41769 53481 41803
rect 53481 41769 53515 41803
rect 53515 41769 53524 41803
rect 53472 41760 53524 41769
rect 60740 41760 60792 41812
rect 6828 41556 6880 41608
rect 11336 41599 11388 41608
rect 11336 41565 11345 41599
rect 11345 41565 11379 41599
rect 11379 41565 11388 41599
rect 11336 41556 11388 41565
rect 29368 41624 29420 41676
rect 31760 41624 31812 41676
rect 35440 41692 35492 41744
rect 38568 41692 38620 41744
rect 39396 41624 39448 41676
rect 40040 41667 40092 41676
rect 40040 41633 40049 41667
rect 40049 41633 40083 41667
rect 40083 41633 40092 41667
rect 40040 41624 40092 41633
rect 35072 41556 35124 41608
rect 39304 41599 39356 41608
rect 27712 41488 27764 41540
rect 30748 41488 30800 41540
rect 39304 41565 39313 41599
rect 39313 41565 39347 41599
rect 39347 41565 39356 41599
rect 39304 41556 39356 41565
rect 41236 41556 41288 41608
rect 46112 41624 46164 41676
rect 47676 41692 47728 41744
rect 46756 41667 46808 41676
rect 46756 41633 46765 41667
rect 46765 41633 46799 41667
rect 46799 41633 46808 41667
rect 47400 41667 47452 41676
rect 46756 41624 46808 41633
rect 47400 41633 47409 41667
rect 47409 41633 47443 41667
rect 47443 41633 47452 41667
rect 47400 41624 47452 41633
rect 48780 41624 48832 41676
rect 49608 41556 49660 41608
rect 38568 41488 38620 41540
rect 38752 41488 38804 41540
rect 52276 41624 52328 41676
rect 52552 41624 52604 41676
rect 53380 41624 53432 41676
rect 58164 41624 58216 41676
rect 60832 41624 60884 41676
rect 53472 41556 53524 41608
rect 70492 41692 70544 41744
rect 66812 41667 66864 41676
rect 66812 41633 66821 41667
rect 66821 41633 66855 41667
rect 66855 41633 66864 41667
rect 66812 41624 66864 41633
rect 71872 41624 71924 41676
rect 72148 41624 72200 41676
rect 72424 41624 72476 41676
rect 74264 41624 74316 41676
rect 72792 41556 72844 41608
rect 79784 41760 79836 41812
rect 77392 41735 77444 41744
rect 77392 41701 77401 41735
rect 77401 41701 77435 41735
rect 77435 41701 77444 41735
rect 77392 41692 77444 41701
rect 77116 41624 77168 41676
rect 77852 41667 77904 41676
rect 77852 41633 77861 41667
rect 77861 41633 77895 41667
rect 77895 41633 77904 41667
rect 77852 41624 77904 41633
rect 83372 41599 83424 41608
rect 83372 41565 83381 41599
rect 83381 41565 83415 41599
rect 83415 41565 83424 41599
rect 83372 41556 83424 41565
rect 83648 41599 83700 41608
rect 83648 41565 83657 41599
rect 83657 41565 83691 41599
rect 83691 41565 83700 41599
rect 83648 41556 83700 41565
rect 77484 41488 77536 41540
rect 12532 41420 12584 41472
rect 26608 41420 26660 41472
rect 27988 41463 28040 41472
rect 27988 41429 27997 41463
rect 27997 41429 28031 41463
rect 28031 41429 28040 41463
rect 27988 41420 28040 41429
rect 40500 41463 40552 41472
rect 40500 41429 40509 41463
rect 40509 41429 40543 41463
rect 40543 41429 40552 41463
rect 40500 41420 40552 41429
rect 41604 41420 41656 41472
rect 45468 41463 45520 41472
rect 45468 41429 45477 41463
rect 45477 41429 45511 41463
rect 45511 41429 45520 41463
rect 45468 41420 45520 41429
rect 51816 41463 51868 41472
rect 51816 41429 51825 41463
rect 51825 41429 51859 41463
rect 51859 41429 51868 41463
rect 51816 41420 51868 41429
rect 52552 41420 52604 41472
rect 66628 41420 66680 41472
rect 72608 41463 72660 41472
rect 72608 41429 72617 41463
rect 72617 41429 72651 41463
rect 72651 41429 72660 41463
rect 72608 41420 72660 41429
rect 78956 41463 79008 41472
rect 78956 41429 78965 41463
rect 78965 41429 78999 41463
rect 78999 41429 79008 41463
rect 78956 41420 79008 41429
rect 84568 41420 84620 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 65686 41318 65738 41370
rect 65750 41318 65802 41370
rect 65814 41318 65866 41370
rect 65878 41318 65930 41370
rect 96406 41318 96458 41370
rect 96470 41318 96522 41370
rect 96534 41318 96586 41370
rect 96598 41318 96650 41370
rect 4068 41216 4120 41268
rect 7012 41216 7064 41268
rect 4712 41148 4764 41200
rect 3976 41123 4028 41132
rect 3976 41089 3985 41123
rect 3985 41089 4019 41123
rect 4019 41089 4028 41123
rect 3976 41080 4028 41089
rect 2596 41055 2648 41064
rect 2596 41021 2612 41055
rect 2612 41021 2646 41055
rect 2646 41021 2648 41055
rect 2596 41012 2648 41021
rect 4620 41012 4672 41064
rect 5540 41012 5592 41064
rect 6828 41055 6880 41064
rect 3608 40944 3660 40996
rect 6828 41021 6837 41055
rect 6837 41021 6871 41055
rect 6871 41021 6880 41055
rect 6828 41012 6880 41021
rect 11060 41216 11112 41268
rect 11336 41259 11388 41268
rect 11336 41225 11345 41259
rect 11345 41225 11379 41259
rect 11379 41225 11388 41259
rect 11336 41216 11388 41225
rect 11428 41216 11480 41268
rect 16764 41216 16816 41268
rect 18420 41216 18472 41268
rect 27712 41259 27764 41268
rect 16580 41148 16632 41200
rect 27712 41225 27721 41259
rect 27721 41225 27755 41259
rect 27755 41225 27764 41259
rect 27712 41216 27764 41225
rect 30564 41216 30616 41268
rect 38844 41216 38896 41268
rect 40224 41259 40276 41268
rect 40224 41225 40233 41259
rect 40233 41225 40267 41259
rect 40267 41225 40276 41259
rect 40224 41216 40276 41225
rect 42064 41259 42116 41268
rect 42064 41225 42073 41259
rect 42073 41225 42107 41259
rect 42107 41225 42116 41259
rect 42064 41216 42116 41225
rect 45468 41148 45520 41200
rect 46756 41148 46808 41200
rect 49608 41216 49660 41268
rect 55864 41216 55916 41268
rect 72792 41259 72844 41268
rect 12716 41055 12768 41064
rect 12716 41021 12725 41055
rect 12725 41021 12759 41055
rect 12759 41021 12768 41055
rect 12716 41012 12768 41021
rect 17408 41080 17460 41132
rect 18696 41123 18748 41132
rect 18696 41089 18705 41123
rect 18705 41089 18739 41123
rect 18739 41089 18748 41123
rect 18696 41080 18748 41089
rect 19432 41123 19484 41132
rect 19432 41089 19441 41123
rect 19441 41089 19475 41123
rect 19475 41089 19484 41123
rect 19432 41080 19484 41089
rect 23756 41080 23808 41132
rect 26516 41080 26568 41132
rect 13452 41055 13504 41064
rect 13452 41021 13461 41055
rect 13461 41021 13495 41055
rect 13495 41021 13504 41055
rect 13452 41012 13504 41021
rect 13728 41012 13780 41064
rect 14004 41055 14056 41064
rect 14004 41021 14013 41055
rect 14013 41021 14047 41055
rect 14047 41021 14056 41055
rect 14004 41012 14056 41021
rect 7012 40876 7064 40928
rect 7564 40876 7616 40928
rect 19248 41012 19300 41064
rect 11060 40876 11112 40928
rect 13084 40919 13136 40928
rect 13084 40885 13093 40919
rect 13093 40885 13127 40919
rect 13127 40885 13136 40919
rect 13084 40876 13136 40885
rect 19432 40944 19484 40996
rect 24124 41055 24176 41064
rect 24124 41021 24133 41055
rect 24133 41021 24167 41055
rect 24167 41021 24176 41055
rect 24676 41055 24728 41064
rect 24124 41012 24176 41021
rect 24676 41021 24685 41055
rect 24685 41021 24719 41055
rect 24719 41021 24728 41055
rect 24676 41012 24728 41021
rect 26148 41055 26200 41064
rect 26148 41021 26157 41055
rect 26157 41021 26191 41055
rect 26191 41021 26200 41055
rect 26148 41012 26200 41021
rect 27988 41012 28040 41064
rect 21824 40876 21876 40928
rect 23756 40919 23808 40928
rect 23756 40885 23765 40919
rect 23765 40885 23799 40919
rect 23799 40885 23808 40919
rect 23756 40876 23808 40885
rect 26148 40876 26200 40928
rect 27896 40919 27948 40928
rect 27896 40885 27905 40919
rect 27905 40885 27939 40919
rect 27939 40885 27948 40919
rect 27896 40876 27948 40885
rect 29184 40876 29236 40928
rect 40408 41080 40460 41132
rect 40592 41080 40644 41132
rect 41696 41123 41748 41132
rect 29644 41012 29696 41064
rect 30564 41055 30616 41064
rect 30564 41021 30573 41055
rect 30573 41021 30607 41055
rect 30607 41021 30616 41055
rect 30564 41012 30616 41021
rect 33416 40944 33468 40996
rect 38016 41012 38068 41064
rect 38752 41012 38804 41064
rect 38660 40944 38712 40996
rect 39396 41012 39448 41064
rect 39120 40944 39172 40996
rect 41696 41089 41705 41123
rect 41705 41089 41739 41123
rect 41739 41089 41748 41123
rect 41696 41080 41748 41089
rect 59176 41148 59228 41200
rect 60832 41191 60884 41200
rect 60832 41157 60841 41191
rect 60841 41157 60875 41191
rect 60875 41157 60884 41191
rect 60832 41148 60884 41157
rect 61108 41191 61160 41200
rect 61108 41157 61117 41191
rect 61117 41157 61151 41191
rect 61151 41157 61160 41191
rect 61108 41148 61160 41157
rect 64328 41148 64380 41200
rect 66444 41148 66496 41200
rect 72792 41225 72801 41259
rect 72801 41225 72835 41259
rect 72835 41225 72844 41259
rect 72792 41216 72844 41225
rect 40592 40944 40644 40996
rect 41236 41055 41288 41064
rect 41236 41021 41245 41055
rect 41245 41021 41279 41055
rect 41279 41021 41288 41055
rect 41236 41012 41288 41021
rect 41420 41012 41472 41064
rect 47400 41055 47452 41064
rect 42064 40944 42116 40996
rect 47400 41021 47409 41055
rect 47409 41021 47443 41055
rect 47443 41021 47452 41055
rect 47400 41012 47452 41021
rect 53196 41080 53248 41132
rect 53472 41123 53524 41132
rect 53472 41089 53481 41123
rect 53481 41089 53515 41123
rect 53515 41089 53524 41123
rect 53472 41080 53524 41089
rect 59268 41123 59320 41132
rect 59268 41089 59277 41123
rect 59277 41089 59311 41123
rect 59311 41089 59320 41123
rect 59268 41080 59320 41089
rect 59544 41123 59596 41132
rect 59544 41089 59553 41123
rect 59553 41089 59587 41123
rect 59587 41089 59596 41123
rect 59544 41080 59596 41089
rect 66904 41080 66956 41132
rect 71872 41080 71924 41132
rect 58900 41012 58952 41064
rect 65340 41055 65392 41064
rect 65340 41021 65349 41055
rect 65349 41021 65383 41055
rect 65383 41021 65392 41055
rect 65340 41012 65392 41021
rect 65984 41012 66036 41064
rect 66628 41055 66680 41064
rect 66628 41021 66637 41055
rect 66637 41021 66671 41055
rect 66671 41021 66680 41055
rect 66628 41012 66680 41021
rect 38016 40919 38068 40928
rect 38016 40885 38025 40919
rect 38025 40885 38059 40919
rect 38059 40885 38068 40919
rect 38016 40876 38068 40885
rect 39304 40876 39356 40928
rect 39580 40876 39632 40928
rect 40224 40876 40276 40928
rect 41052 40876 41104 40928
rect 48228 40944 48280 40996
rect 48136 40876 48188 40928
rect 48780 40876 48832 40928
rect 54484 40876 54536 40928
rect 58716 40876 58768 40928
rect 66720 40944 66772 40996
rect 67088 40987 67140 40996
rect 67088 40953 67097 40987
rect 67097 40953 67131 40987
rect 67131 40953 67140 40987
rect 67088 40944 67140 40953
rect 67364 41012 67416 41064
rect 71596 41012 71648 41064
rect 83740 41148 83792 41200
rect 71688 40944 71740 40996
rect 72424 41080 72476 41132
rect 72700 41123 72752 41132
rect 72700 41089 72709 41123
rect 72709 41089 72743 41123
rect 72743 41089 72752 41123
rect 72700 41080 72752 41089
rect 72332 41055 72384 41064
rect 72332 41021 72346 41055
rect 72346 41021 72384 41055
rect 72332 41012 72384 41021
rect 76196 41055 76248 41064
rect 76196 41021 76205 41055
rect 76205 41021 76239 41055
rect 76239 41021 76248 41055
rect 76196 41012 76248 41021
rect 77208 41055 77260 41064
rect 77208 41021 77217 41055
rect 77217 41021 77251 41055
rect 77251 41021 77260 41055
rect 77208 41012 77260 41021
rect 77668 41080 77720 41132
rect 77484 41012 77536 41064
rect 72516 40944 72568 40996
rect 84108 40944 84160 40996
rect 66904 40876 66956 40928
rect 67640 40876 67692 40928
rect 71780 40919 71832 40928
rect 71780 40885 71789 40919
rect 71789 40885 71823 40919
rect 71823 40885 71832 40919
rect 71780 40876 71832 40885
rect 76196 40876 76248 40928
rect 78956 40876 79008 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 81046 40774 81098 40826
rect 81110 40774 81162 40826
rect 81174 40774 81226 40826
rect 81238 40774 81290 40826
rect 7748 40672 7800 40724
rect 10140 40672 10192 40724
rect 11060 40672 11112 40724
rect 12716 40672 12768 40724
rect 13452 40672 13504 40724
rect 5540 40604 5592 40656
rect 3056 40468 3108 40520
rect 6828 40536 6880 40588
rect 13084 40604 13136 40656
rect 13544 40604 13596 40656
rect 10232 40579 10284 40588
rect 10232 40545 10241 40579
rect 10241 40545 10275 40579
rect 10275 40545 10284 40579
rect 10232 40536 10284 40545
rect 12532 40579 12584 40588
rect 12532 40545 12541 40579
rect 12541 40545 12575 40579
rect 12575 40545 12584 40579
rect 12532 40536 12584 40545
rect 19248 40604 19300 40656
rect 20352 40647 20404 40656
rect 7840 40468 7892 40520
rect 11428 40468 11480 40520
rect 19524 40536 19576 40588
rect 16028 40511 16080 40520
rect 16028 40477 16037 40511
rect 16037 40477 16071 40511
rect 16071 40477 16080 40511
rect 16028 40468 16080 40477
rect 18420 40468 18472 40520
rect 20352 40613 20361 40647
rect 20361 40613 20395 40647
rect 20395 40613 20404 40647
rect 20352 40604 20404 40613
rect 26976 40604 27028 40656
rect 27344 40672 27396 40724
rect 27436 40672 27488 40724
rect 41512 40672 41564 40724
rect 41604 40672 41656 40724
rect 55864 40672 55916 40724
rect 58440 40715 58492 40724
rect 58440 40681 58449 40715
rect 58449 40681 58483 40715
rect 58483 40681 58492 40715
rect 58440 40672 58492 40681
rect 58900 40672 58952 40724
rect 65432 40672 65484 40724
rect 71688 40672 71740 40724
rect 76196 40672 76248 40724
rect 77760 40672 77812 40724
rect 84108 40672 84160 40724
rect 21916 40468 21968 40520
rect 22376 40511 22428 40520
rect 22376 40477 22385 40511
rect 22385 40477 22419 40511
rect 22419 40477 22428 40511
rect 22376 40468 22428 40477
rect 27252 40536 27304 40588
rect 29000 40604 29052 40656
rect 27988 40468 28040 40520
rect 29460 40536 29512 40588
rect 34152 40604 34204 40656
rect 40224 40647 40276 40656
rect 29092 40468 29144 40520
rect 29184 40468 29236 40520
rect 38844 40579 38896 40588
rect 38844 40545 38853 40579
rect 38853 40545 38887 40579
rect 38887 40545 38896 40579
rect 38844 40536 38896 40545
rect 39396 40579 39448 40588
rect 39396 40545 39405 40579
rect 39405 40545 39439 40579
rect 39439 40545 39448 40579
rect 39396 40536 39448 40545
rect 39580 40579 39632 40588
rect 39580 40545 39589 40579
rect 39589 40545 39623 40579
rect 39623 40545 39632 40579
rect 39580 40536 39632 40545
rect 40224 40613 40233 40647
rect 40233 40613 40267 40647
rect 40267 40613 40276 40647
rect 40224 40604 40276 40613
rect 40684 40604 40736 40656
rect 40776 40604 40828 40656
rect 40960 40604 41012 40656
rect 52736 40604 52788 40656
rect 52828 40604 52880 40656
rect 58808 40604 58860 40656
rect 61568 40604 61620 40656
rect 83648 40604 83700 40656
rect 44456 40536 44508 40588
rect 31760 40468 31812 40520
rect 32956 40468 33008 40520
rect 33416 40511 33468 40520
rect 33416 40477 33425 40511
rect 33425 40477 33459 40511
rect 33459 40477 33468 40511
rect 33416 40468 33468 40477
rect 38568 40511 38620 40520
rect 38568 40477 38577 40511
rect 38577 40477 38611 40511
rect 38611 40477 38620 40511
rect 38568 40468 38620 40477
rect 44824 40536 44876 40588
rect 46572 40536 46624 40588
rect 9864 40332 9916 40384
rect 12532 40332 12584 40384
rect 21088 40332 21140 40384
rect 21916 40375 21968 40384
rect 21916 40341 21925 40375
rect 21925 40341 21959 40375
rect 21959 40341 21968 40375
rect 21916 40332 21968 40341
rect 23664 40375 23716 40384
rect 23664 40341 23673 40375
rect 23673 40341 23707 40375
rect 23707 40341 23716 40375
rect 23664 40332 23716 40341
rect 24676 40332 24728 40384
rect 29000 40332 29052 40384
rect 29184 40375 29236 40384
rect 29184 40341 29193 40375
rect 29193 40341 29227 40375
rect 29227 40341 29236 40375
rect 29184 40332 29236 40341
rect 32956 40375 33008 40384
rect 32956 40341 32965 40375
rect 32965 40341 32999 40375
rect 32999 40341 33008 40375
rect 32956 40332 33008 40341
rect 40592 40400 40644 40452
rect 44364 40400 44416 40452
rect 34704 40375 34756 40384
rect 34704 40341 34713 40375
rect 34713 40341 34747 40375
rect 34747 40341 34756 40375
rect 34704 40332 34756 40341
rect 40500 40332 40552 40384
rect 41512 40375 41564 40384
rect 41512 40341 41521 40375
rect 41521 40341 41555 40375
rect 41555 40341 41564 40375
rect 41512 40332 41564 40341
rect 41604 40332 41656 40384
rect 44180 40332 44232 40384
rect 44916 40468 44968 40520
rect 45744 40468 45796 40520
rect 48872 40468 48924 40520
rect 44640 40400 44692 40452
rect 52460 40536 52512 40588
rect 52920 40536 52972 40588
rect 58072 40536 58124 40588
rect 58440 40536 58492 40588
rect 59176 40536 59228 40588
rect 59728 40536 59780 40588
rect 67088 40536 67140 40588
rect 52828 40468 52880 40520
rect 53012 40511 53064 40520
rect 53012 40477 53021 40511
rect 53021 40477 53055 40511
rect 53055 40477 53064 40511
rect 53012 40468 53064 40477
rect 53104 40468 53156 40520
rect 65340 40468 65392 40520
rect 45560 40332 45612 40384
rect 45744 40375 45796 40384
rect 45744 40341 45753 40375
rect 45753 40341 45787 40375
rect 45787 40341 45796 40375
rect 45744 40332 45796 40341
rect 46020 40375 46072 40384
rect 46020 40341 46029 40375
rect 46029 40341 46063 40375
rect 46063 40341 46072 40375
rect 46020 40332 46072 40341
rect 46572 40332 46624 40384
rect 49516 40332 49568 40384
rect 54300 40400 54352 40452
rect 63132 40400 63184 40452
rect 66812 40468 66864 40520
rect 67456 40468 67508 40520
rect 72424 40511 72476 40520
rect 72424 40477 72433 40511
rect 72433 40477 72467 40511
rect 72467 40477 72476 40511
rect 72424 40468 72476 40477
rect 72608 40468 72660 40520
rect 77208 40468 77260 40520
rect 77484 40536 77536 40588
rect 83556 40579 83608 40588
rect 83556 40545 83565 40579
rect 83565 40545 83599 40579
rect 83599 40545 83608 40579
rect 83556 40536 83608 40545
rect 83740 40579 83792 40588
rect 83740 40545 83749 40579
rect 83749 40545 83783 40579
rect 83783 40545 83792 40579
rect 83740 40536 83792 40545
rect 84568 40579 84620 40588
rect 84568 40545 84577 40579
rect 84577 40545 84611 40579
rect 84611 40545 84620 40579
rect 84568 40536 84620 40545
rect 83280 40511 83332 40520
rect 83280 40477 83289 40511
rect 83289 40477 83323 40511
rect 83323 40477 83332 40511
rect 83280 40468 83332 40477
rect 53932 40332 53984 40384
rect 58716 40332 58768 40384
rect 61016 40332 61068 40384
rect 61752 40332 61804 40384
rect 73528 40375 73580 40384
rect 73528 40341 73537 40375
rect 73537 40341 73571 40375
rect 73571 40341 73580 40375
rect 73528 40332 73580 40341
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 65686 40230 65738 40282
rect 65750 40230 65802 40282
rect 65814 40230 65866 40282
rect 65878 40230 65930 40282
rect 96406 40230 96458 40282
rect 96470 40230 96522 40282
rect 96534 40230 96586 40282
rect 96598 40230 96650 40282
rect 3884 40128 3936 40180
rect 4804 40060 4856 40112
rect 4988 40060 5040 40112
rect 10232 40128 10284 40180
rect 27344 40128 27396 40180
rect 27528 40128 27580 40180
rect 27712 40128 27764 40180
rect 29460 40171 29512 40180
rect 29460 40137 29469 40171
rect 29469 40137 29503 40171
rect 29503 40137 29512 40171
rect 29460 40128 29512 40137
rect 34704 40128 34756 40180
rect 57796 40171 57848 40180
rect 57796 40137 57805 40171
rect 57805 40137 57839 40171
rect 57839 40137 57848 40171
rect 57796 40128 57848 40137
rect 58808 40171 58860 40180
rect 58808 40137 58817 40171
rect 58817 40137 58851 40171
rect 58851 40137 58860 40171
rect 58808 40128 58860 40137
rect 72424 40128 72476 40180
rect 74264 40171 74316 40180
rect 74264 40137 74273 40171
rect 74273 40137 74307 40171
rect 74307 40137 74316 40171
rect 74264 40128 74316 40137
rect 83740 40171 83792 40180
rect 83740 40137 83749 40171
rect 83749 40137 83783 40171
rect 83783 40137 83792 40171
rect 83740 40128 83792 40137
rect 12532 40060 12584 40112
rect 38568 40060 38620 40112
rect 40500 40060 40552 40112
rect 45744 40060 45796 40112
rect 4804 39924 4856 39976
rect 9404 39924 9456 39976
rect 17132 39992 17184 40044
rect 18420 40035 18472 40044
rect 17316 39924 17368 39976
rect 18420 40001 18429 40035
rect 18429 40001 18463 40035
rect 18463 40001 18472 40035
rect 18420 39992 18472 40001
rect 40684 40035 40736 40044
rect 40684 40001 40690 40035
rect 40690 40001 40736 40035
rect 40684 39992 40736 40001
rect 23664 39967 23716 39976
rect 23664 39933 23673 39967
rect 23673 39933 23707 39967
rect 23707 39933 23716 39967
rect 23664 39924 23716 39933
rect 28448 39924 28500 39976
rect 29460 39924 29512 39976
rect 15568 39856 15620 39908
rect 22744 39856 22796 39908
rect 40316 39924 40368 39976
rect 40408 39924 40460 39976
rect 38936 39856 38988 39908
rect 40960 39992 41012 40044
rect 41696 39992 41748 40044
rect 44456 39992 44508 40044
rect 44916 39992 44968 40044
rect 46020 39992 46072 40044
rect 46848 39924 46900 39976
rect 48136 40060 48188 40112
rect 48780 40060 48832 40112
rect 53104 40060 53156 40112
rect 54116 40103 54168 40112
rect 54116 40069 54140 40103
rect 54140 40069 54168 40103
rect 54116 40060 54168 40069
rect 54392 40060 54444 40112
rect 52460 39992 52512 40044
rect 54668 39992 54720 40044
rect 54852 40103 54904 40112
rect 54852 40069 54861 40103
rect 54861 40069 54895 40103
rect 54895 40069 54904 40103
rect 54852 40060 54904 40069
rect 59544 40060 59596 40112
rect 83280 40060 83332 40112
rect 44272 39856 44324 39908
rect 51080 39924 51132 39976
rect 53380 39924 53432 39976
rect 53932 39967 53984 39976
rect 53932 39933 53941 39967
rect 53941 39933 53975 39967
rect 53975 39933 53984 39967
rect 53932 39924 53984 39933
rect 54208 39924 54260 39976
rect 57796 39924 57848 39976
rect 58072 39967 58124 39976
rect 58072 39933 58081 39967
rect 58081 39933 58115 39967
rect 58115 39933 58124 39967
rect 58072 39924 58124 39933
rect 58808 39924 58860 39976
rect 59176 39967 59228 39976
rect 59176 39933 59185 39967
rect 59185 39933 59219 39967
rect 59219 39933 59228 39967
rect 59176 39924 59228 39933
rect 48228 39856 48280 39908
rect 49056 39856 49108 39908
rect 54392 39856 54444 39908
rect 10600 39831 10652 39840
rect 10600 39797 10609 39831
rect 10609 39797 10643 39831
rect 10643 39797 10652 39831
rect 10600 39788 10652 39797
rect 15108 39788 15160 39840
rect 16580 39788 16632 39840
rect 17316 39831 17368 39840
rect 17316 39797 17325 39831
rect 17325 39797 17359 39831
rect 17359 39797 17368 39831
rect 17316 39788 17368 39797
rect 19340 39788 19392 39840
rect 24124 39788 24176 39840
rect 29460 39788 29512 39840
rect 32404 39788 32456 39840
rect 40868 39788 40920 39840
rect 46848 39831 46900 39840
rect 46848 39797 46857 39831
rect 46857 39797 46891 39831
rect 46891 39797 46900 39831
rect 46848 39788 46900 39797
rect 46940 39788 46992 39840
rect 59544 39856 59596 39908
rect 56508 39788 56560 39840
rect 57796 39788 57848 39840
rect 59452 39788 59504 39840
rect 60556 39924 60608 39976
rect 71136 39924 71188 39976
rect 72148 39924 72200 39976
rect 72516 39967 72568 39976
rect 60832 39856 60884 39908
rect 65156 39856 65208 39908
rect 66076 39856 66128 39908
rect 67640 39856 67692 39908
rect 72516 39933 72525 39967
rect 72525 39933 72559 39967
rect 72559 39933 72568 39967
rect 72516 39924 72568 39933
rect 60004 39788 60056 39840
rect 67364 39788 67416 39840
rect 71688 39788 71740 39840
rect 72608 39856 72660 39908
rect 79692 39992 79744 40044
rect 83556 39992 83608 40044
rect 73528 39924 73580 39976
rect 77208 39924 77260 39976
rect 82176 39924 82228 39976
rect 82268 39856 82320 39908
rect 83740 39924 83792 39976
rect 77576 39831 77628 39840
rect 77576 39797 77585 39831
rect 77585 39797 77619 39831
rect 77619 39797 77628 39831
rect 77576 39788 77628 39797
rect 77760 39788 77812 39840
rect 82360 39831 82412 39840
rect 82360 39797 82369 39831
rect 82369 39797 82403 39831
rect 82403 39797 82412 39831
rect 82360 39788 82412 39797
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 81046 39686 81098 39738
rect 81110 39686 81162 39738
rect 81174 39686 81226 39738
rect 81238 39686 81290 39738
rect 3792 39584 3844 39636
rect 12072 39584 12124 39636
rect 22376 39627 22428 39636
rect 22376 39593 22385 39627
rect 22385 39593 22419 39627
rect 22419 39593 22428 39627
rect 22376 39584 22428 39593
rect 22744 39627 22796 39636
rect 22744 39593 22753 39627
rect 22753 39593 22787 39627
rect 22787 39593 22796 39627
rect 22744 39584 22796 39593
rect 24124 39584 24176 39636
rect 38016 39584 38068 39636
rect 44272 39584 44324 39636
rect 44364 39584 44416 39636
rect 46020 39584 46072 39636
rect 46940 39584 46992 39636
rect 4620 39448 4672 39500
rect 9128 39448 9180 39500
rect 4712 39244 4764 39296
rect 9128 39244 9180 39296
rect 21088 39448 21140 39500
rect 21364 39491 21416 39500
rect 21364 39457 21373 39491
rect 21373 39457 21407 39491
rect 21407 39457 21416 39491
rect 21364 39448 21416 39457
rect 16396 39423 16448 39432
rect 16396 39389 16405 39423
rect 16405 39389 16439 39423
rect 16439 39389 16448 39423
rect 16396 39380 16448 39389
rect 17868 39380 17920 39432
rect 19248 39244 19300 39296
rect 20720 39244 20772 39296
rect 21364 39312 21416 39364
rect 27896 39448 27948 39500
rect 32956 39516 33008 39568
rect 44824 39516 44876 39568
rect 39028 39491 39080 39500
rect 39028 39457 39037 39491
rect 39037 39457 39071 39491
rect 39071 39457 39080 39491
rect 39028 39448 39080 39457
rect 39488 39491 39540 39500
rect 39488 39457 39497 39491
rect 39497 39457 39531 39491
rect 39531 39457 39540 39491
rect 39488 39448 39540 39457
rect 39948 39448 40000 39500
rect 43812 39448 43864 39500
rect 44180 39491 44232 39500
rect 44180 39457 44189 39491
rect 44189 39457 44223 39491
rect 44223 39457 44232 39491
rect 44180 39448 44232 39457
rect 28264 39423 28316 39432
rect 28264 39389 28273 39423
rect 28273 39389 28307 39423
rect 28307 39389 28316 39423
rect 28264 39380 28316 39389
rect 33324 39423 33376 39432
rect 33324 39389 33333 39423
rect 33333 39389 33367 39423
rect 33367 39389 33376 39423
rect 33324 39380 33376 39389
rect 38936 39423 38988 39432
rect 38936 39389 38945 39423
rect 38945 39389 38979 39423
rect 38979 39389 38988 39423
rect 38936 39380 38988 39389
rect 44456 39491 44508 39500
rect 44456 39457 44465 39491
rect 44465 39457 44499 39491
rect 44499 39457 44508 39491
rect 44916 39491 44968 39500
rect 44456 39448 44508 39457
rect 44916 39457 44925 39491
rect 44925 39457 44959 39491
rect 44959 39457 44968 39491
rect 44916 39448 44968 39457
rect 26700 39312 26752 39364
rect 29552 39287 29604 39296
rect 29552 39253 29561 39287
rect 29561 39253 29595 39287
rect 29595 39253 29604 39287
rect 29552 39244 29604 39253
rect 34612 39287 34664 39296
rect 34612 39253 34621 39287
rect 34621 39253 34655 39287
rect 34655 39253 34664 39287
rect 34612 39244 34664 39253
rect 39580 39244 39632 39296
rect 40040 39287 40092 39296
rect 40040 39253 40049 39287
rect 40049 39253 40083 39287
rect 40083 39253 40092 39287
rect 40040 39244 40092 39253
rect 40684 39244 40736 39296
rect 42616 39244 42668 39296
rect 46572 39380 46624 39432
rect 47032 39448 47084 39500
rect 48044 39584 48096 39636
rect 48136 39516 48188 39568
rect 48780 39516 48832 39568
rect 48872 39516 48924 39568
rect 54392 39516 54444 39568
rect 54484 39516 54536 39568
rect 47400 39491 47452 39500
rect 47400 39457 47409 39491
rect 47409 39457 47443 39491
rect 47443 39457 47452 39491
rect 47400 39448 47452 39457
rect 47584 39448 47636 39500
rect 51816 39448 51868 39500
rect 52276 39491 52328 39500
rect 52276 39457 52285 39491
rect 52285 39457 52319 39491
rect 52319 39457 52328 39491
rect 52276 39448 52328 39457
rect 48136 39380 48188 39432
rect 51724 39380 51776 39432
rect 52828 39491 52880 39500
rect 52828 39457 52837 39491
rect 52837 39457 52871 39491
rect 52871 39457 52880 39491
rect 52828 39448 52880 39457
rect 53656 39423 53708 39432
rect 53656 39389 53665 39423
rect 53665 39389 53699 39423
rect 53699 39389 53708 39423
rect 53656 39380 53708 39389
rect 55220 39516 55272 39568
rect 58440 39584 58492 39636
rect 60372 39584 60424 39636
rect 60832 39584 60884 39636
rect 60740 39516 60792 39568
rect 54852 39448 54904 39500
rect 60832 39491 60884 39500
rect 54944 39423 54996 39432
rect 54944 39389 54950 39423
rect 54950 39389 54984 39423
rect 54984 39389 54996 39423
rect 54944 39380 54996 39389
rect 55220 39380 55272 39432
rect 60556 39380 60608 39432
rect 54208 39312 54260 39364
rect 54576 39312 54628 39364
rect 47308 39244 47360 39296
rect 47400 39244 47452 39296
rect 47860 39244 47912 39296
rect 51724 39287 51776 39296
rect 51724 39253 51733 39287
rect 51733 39253 51767 39287
rect 51767 39253 51776 39287
rect 51724 39244 51776 39253
rect 52276 39244 52328 39296
rect 52828 39244 52880 39296
rect 53288 39287 53340 39296
rect 53288 39253 53297 39287
rect 53297 39253 53331 39287
rect 53331 39253 53340 39287
rect 53288 39244 53340 39253
rect 60096 39312 60148 39364
rect 60832 39457 60841 39491
rect 60841 39457 60875 39491
rect 60875 39457 60884 39491
rect 60832 39448 60884 39457
rect 67364 39584 67416 39636
rect 69756 39584 69808 39636
rect 71688 39584 71740 39636
rect 66076 39516 66128 39568
rect 71596 39559 71648 39568
rect 71596 39525 71605 39559
rect 71605 39525 71639 39559
rect 71639 39525 71648 39559
rect 71964 39584 72016 39636
rect 72516 39584 72568 39636
rect 77760 39627 77812 39636
rect 77760 39593 77769 39627
rect 77769 39593 77803 39627
rect 77803 39593 77812 39627
rect 77760 39584 77812 39593
rect 83372 39584 83424 39636
rect 71596 39516 71648 39525
rect 61200 39491 61252 39500
rect 61200 39457 61209 39491
rect 61209 39457 61243 39491
rect 61243 39457 61252 39491
rect 61200 39448 61252 39457
rect 61568 39448 61620 39500
rect 61936 39448 61988 39500
rect 65524 39448 65576 39500
rect 66812 39448 66864 39500
rect 67456 39448 67508 39500
rect 71412 39448 71464 39500
rect 71780 39491 71832 39500
rect 71780 39457 71789 39491
rect 71789 39457 71823 39491
rect 71823 39457 71832 39491
rect 71780 39448 71832 39457
rect 72148 39491 72200 39500
rect 72148 39457 72157 39491
rect 72157 39457 72191 39491
rect 72191 39457 72200 39491
rect 72148 39448 72200 39457
rect 68836 39380 68888 39432
rect 71596 39380 71648 39432
rect 71964 39380 72016 39432
rect 66076 39312 66128 39364
rect 71136 39312 71188 39364
rect 72424 39312 72476 39364
rect 79692 39516 79744 39568
rect 78220 39491 78272 39500
rect 78220 39457 78229 39491
rect 78229 39457 78263 39491
rect 78263 39457 78272 39491
rect 78220 39448 78272 39457
rect 86316 39448 86368 39500
rect 84384 39380 84436 39432
rect 57888 39244 57940 39296
rect 60280 39287 60332 39296
rect 60280 39253 60289 39287
rect 60289 39253 60323 39287
rect 60323 39253 60332 39287
rect 60280 39244 60332 39253
rect 60372 39244 60424 39296
rect 61200 39244 61252 39296
rect 66904 39244 66956 39296
rect 71412 39287 71464 39296
rect 71412 39253 71421 39287
rect 71421 39253 71455 39287
rect 71455 39253 71464 39287
rect 71412 39244 71464 39253
rect 78404 39287 78456 39296
rect 78404 39253 78413 39287
rect 78413 39253 78447 39287
rect 78447 39253 78456 39287
rect 78404 39244 78456 39253
rect 85396 39244 85448 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 65686 39142 65738 39194
rect 65750 39142 65802 39194
rect 65814 39142 65866 39194
rect 65878 39142 65930 39194
rect 96406 39142 96458 39194
rect 96470 39142 96522 39194
rect 96534 39142 96586 39194
rect 96598 39142 96650 39194
rect 4620 39040 4672 39092
rect 4804 39083 4856 39092
rect 4804 39049 4813 39083
rect 4813 39049 4847 39083
rect 4847 39049 4856 39083
rect 4804 39040 4856 39049
rect 9864 39083 9916 39092
rect 4804 38904 4856 38956
rect 4620 38836 4672 38888
rect 3516 38700 3568 38752
rect 9864 39049 9873 39083
rect 9873 39049 9907 39083
rect 9907 39049 9916 39083
rect 9864 39040 9916 39049
rect 13544 39040 13596 39092
rect 13820 39083 13872 39092
rect 13820 39049 13829 39083
rect 13829 39049 13863 39083
rect 13863 39049 13872 39083
rect 13820 39040 13872 39049
rect 17132 39040 17184 39092
rect 22192 39040 22244 39092
rect 28448 39083 28500 39092
rect 9404 39015 9456 39024
rect 9404 38981 9413 39015
rect 9413 38981 9447 39015
rect 9447 38981 9456 39015
rect 9404 38972 9456 38981
rect 10232 38972 10284 39024
rect 15108 38972 15160 39024
rect 16028 39015 16080 39024
rect 16028 38981 16037 39015
rect 16037 38981 16071 39015
rect 16071 38981 16080 39015
rect 16028 38972 16080 38981
rect 26700 38972 26752 39024
rect 28448 39049 28457 39083
rect 28457 39049 28491 39083
rect 28491 39049 28500 39083
rect 28448 39040 28500 39049
rect 29552 39040 29604 39092
rect 53104 39040 53156 39092
rect 53288 39040 53340 39092
rect 54668 39083 54720 39092
rect 54668 39049 54677 39083
rect 54677 39049 54711 39083
rect 54711 39049 54720 39083
rect 54668 39040 54720 39049
rect 42156 38972 42208 39024
rect 44916 38972 44968 39024
rect 46112 39015 46164 39024
rect 46112 38981 46121 39015
rect 46121 38981 46155 39015
rect 46155 38981 46164 39015
rect 46112 38972 46164 38981
rect 39028 38904 39080 38956
rect 40408 38904 40460 38956
rect 40684 38904 40736 38956
rect 46388 38947 46440 38956
rect 46388 38913 46397 38947
rect 46397 38913 46431 38947
rect 46431 38913 46440 38947
rect 48044 38947 48096 38956
rect 46388 38904 46440 38913
rect 48044 38913 48053 38947
rect 48053 38913 48087 38947
rect 48087 38913 48096 38947
rect 48044 38904 48096 38913
rect 48136 38947 48188 38956
rect 48136 38913 48145 38947
rect 48145 38913 48179 38947
rect 48179 38913 48188 38947
rect 53380 38972 53432 39024
rect 54576 38947 54628 38956
rect 48136 38904 48188 38913
rect 10232 38836 10284 38888
rect 15108 38879 15160 38888
rect 15108 38845 15117 38879
rect 15117 38845 15151 38879
rect 15151 38845 15160 38879
rect 15108 38836 15160 38845
rect 15568 38879 15620 38888
rect 15568 38845 15577 38879
rect 15577 38845 15611 38879
rect 15611 38845 15620 38879
rect 15568 38836 15620 38845
rect 21364 38836 21416 38888
rect 23664 38879 23716 38888
rect 23664 38845 23673 38879
rect 23673 38845 23707 38879
rect 23707 38845 23716 38879
rect 23664 38836 23716 38845
rect 28448 38836 28500 38888
rect 44732 38836 44784 38888
rect 46572 38836 46624 38888
rect 47032 38879 47084 38888
rect 47032 38845 47041 38879
rect 47041 38845 47075 38879
rect 47075 38845 47084 38879
rect 47032 38836 47084 38845
rect 47124 38836 47176 38888
rect 17868 38768 17920 38820
rect 15108 38700 15160 38752
rect 36360 38743 36412 38752
rect 36360 38709 36369 38743
rect 36369 38709 36403 38743
rect 36403 38709 36412 38743
rect 36360 38700 36412 38709
rect 49240 38768 49292 38820
rect 51448 38768 51500 38820
rect 52276 38836 52328 38888
rect 53656 38879 53708 38888
rect 53656 38845 53665 38879
rect 53665 38845 53699 38879
rect 53699 38845 53708 38879
rect 53656 38836 53708 38845
rect 54208 38879 54260 38888
rect 54208 38845 54217 38879
rect 54217 38845 54251 38879
rect 54251 38845 54260 38879
rect 54208 38836 54260 38845
rect 54576 38913 54585 38947
rect 54585 38913 54619 38947
rect 54619 38913 54628 38947
rect 54576 38904 54628 38913
rect 58072 38972 58124 39024
rect 59176 38972 59228 39024
rect 59452 38972 59504 39024
rect 61476 38972 61528 39024
rect 68376 38972 68428 39024
rect 68836 39015 68888 39024
rect 68836 38981 68845 39015
rect 68845 38981 68879 39015
rect 68879 38981 68888 39015
rect 68836 38972 68888 38981
rect 69756 38972 69808 39024
rect 73068 39040 73120 39092
rect 77760 39040 77812 39092
rect 84384 39083 84436 39092
rect 84384 39049 84393 39083
rect 84393 39049 84427 39083
rect 84427 39049 84436 39083
rect 84384 39040 84436 39049
rect 86316 39083 86368 39092
rect 86316 39049 86325 39083
rect 86325 39049 86359 39083
rect 86359 39049 86368 39083
rect 86316 39040 86368 39049
rect 53104 38768 53156 38820
rect 59084 38836 59136 38888
rect 46848 38700 46900 38752
rect 47124 38700 47176 38752
rect 52736 38700 52788 38752
rect 54392 38700 54444 38752
rect 59452 38836 59504 38888
rect 65984 38904 66036 38956
rect 66076 38904 66128 38956
rect 69296 38904 69348 38956
rect 71412 38904 71464 38956
rect 59728 38768 59780 38820
rect 61660 38836 61712 38888
rect 61936 38879 61988 38888
rect 61936 38845 61945 38879
rect 61945 38845 61979 38879
rect 61979 38845 61988 38879
rect 61936 38836 61988 38845
rect 64972 38879 65024 38888
rect 64972 38845 64981 38879
rect 64981 38845 65015 38879
rect 65015 38845 65024 38879
rect 64972 38836 65024 38845
rect 65156 38879 65208 38888
rect 65156 38845 65165 38879
rect 65165 38845 65199 38879
rect 65199 38845 65208 38879
rect 65156 38836 65208 38845
rect 65524 38879 65576 38888
rect 65524 38845 65533 38879
rect 65533 38845 65567 38879
rect 65567 38845 65576 38879
rect 65524 38836 65576 38845
rect 66904 38879 66956 38888
rect 64236 38768 64288 38820
rect 66904 38845 66913 38879
rect 66913 38845 66947 38879
rect 66947 38845 66956 38879
rect 66904 38836 66956 38845
rect 71688 38879 71740 38888
rect 71688 38845 71697 38879
rect 71697 38845 71731 38879
rect 71731 38845 71740 38879
rect 71688 38836 71740 38845
rect 71964 38904 72016 38956
rect 77116 38972 77168 39024
rect 72792 38836 72844 38888
rect 73068 38879 73120 38888
rect 73068 38845 73077 38879
rect 73077 38845 73111 38879
rect 73111 38845 73120 38879
rect 73068 38836 73120 38845
rect 77116 38879 77168 38888
rect 77116 38845 77125 38879
rect 77125 38845 77159 38879
rect 77159 38845 77168 38879
rect 77116 38836 77168 38845
rect 78404 38904 78456 38956
rect 79048 38836 79100 38888
rect 79600 38836 79652 38888
rect 82268 38836 82320 38888
rect 84292 38879 84344 38888
rect 84292 38845 84301 38879
rect 84301 38845 84335 38879
rect 84335 38845 84344 38879
rect 84292 38836 84344 38845
rect 85396 38879 85448 38888
rect 85396 38845 85405 38879
rect 85405 38845 85439 38879
rect 85439 38845 85448 38879
rect 85396 38836 85448 38845
rect 86316 38836 86368 38888
rect 86776 38879 86828 38888
rect 86776 38845 86785 38879
rect 86785 38845 86819 38879
rect 86819 38845 86828 38879
rect 86776 38836 86828 38845
rect 84752 38768 84804 38820
rect 60004 38743 60056 38752
rect 60004 38709 60013 38743
rect 60013 38709 60047 38743
rect 60047 38709 60056 38743
rect 60004 38700 60056 38709
rect 60096 38700 60148 38752
rect 61384 38700 61436 38752
rect 64972 38700 65024 38752
rect 68284 38700 68336 38752
rect 71412 38700 71464 38752
rect 72608 38743 72660 38752
rect 72608 38709 72617 38743
rect 72617 38709 72651 38743
rect 72651 38709 72660 38743
rect 72608 38700 72660 38709
rect 73160 38743 73212 38752
rect 73160 38709 73169 38743
rect 73169 38709 73203 38743
rect 73203 38709 73212 38743
rect 73160 38700 73212 38709
rect 79876 38743 79928 38752
rect 79876 38709 79885 38743
rect 79885 38709 79919 38743
rect 79919 38709 79928 38743
rect 79876 38700 79928 38709
rect 83372 38743 83424 38752
rect 83372 38709 83381 38743
rect 83381 38709 83415 38743
rect 83415 38709 83424 38743
rect 83372 38700 83424 38709
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 81046 38598 81098 38650
rect 81110 38598 81162 38650
rect 81174 38598 81226 38650
rect 81238 38598 81290 38650
rect 4068 38496 4120 38548
rect 23756 38496 23808 38548
rect 12256 38428 12308 38480
rect 10600 38360 10652 38412
rect 11060 38335 11112 38344
rect 11060 38301 11069 38335
rect 11069 38301 11103 38335
rect 11103 38301 11112 38335
rect 11060 38292 11112 38301
rect 13820 38360 13872 38412
rect 17868 38471 17920 38480
rect 17868 38437 17877 38471
rect 17877 38437 17911 38471
rect 17911 38437 17920 38471
rect 17868 38428 17920 38437
rect 20812 38428 20864 38480
rect 21088 38428 21140 38480
rect 15844 38360 15896 38412
rect 16028 38403 16080 38412
rect 16028 38369 16037 38403
rect 16037 38369 16071 38403
rect 16071 38369 16080 38403
rect 16028 38360 16080 38369
rect 16212 38403 16264 38412
rect 16212 38369 16221 38403
rect 16221 38369 16255 38403
rect 16255 38369 16264 38403
rect 16212 38360 16264 38369
rect 23664 38428 23716 38480
rect 26240 38428 26292 38480
rect 16396 38267 16448 38276
rect 16396 38233 16405 38267
rect 16405 38233 16439 38267
rect 16439 38233 16448 38267
rect 16396 38224 16448 38233
rect 5080 38156 5132 38208
rect 12256 38156 12308 38208
rect 12440 38156 12492 38208
rect 15108 38199 15160 38208
rect 15108 38165 15117 38199
rect 15117 38165 15151 38199
rect 15151 38165 15160 38199
rect 15108 38156 15160 38165
rect 15844 38156 15896 38208
rect 26700 38360 26752 38412
rect 28264 38428 28316 38480
rect 37096 38496 37148 38548
rect 40224 38496 40276 38548
rect 40408 38539 40460 38548
rect 40408 38505 40417 38539
rect 40417 38505 40451 38539
rect 40451 38505 40460 38539
rect 40408 38496 40460 38505
rect 40960 38496 41012 38548
rect 51816 38496 51868 38548
rect 54944 38496 54996 38548
rect 55036 38496 55088 38548
rect 72424 38539 72476 38548
rect 64972 38428 65024 38480
rect 38476 38360 38528 38412
rect 21732 38335 21784 38344
rect 21732 38301 21741 38335
rect 21741 38301 21775 38335
rect 21775 38301 21784 38335
rect 21732 38292 21784 38301
rect 23848 38224 23900 38276
rect 32772 38224 32824 38276
rect 33416 38335 33468 38344
rect 33416 38301 33425 38335
rect 33425 38301 33459 38335
rect 33459 38301 33468 38335
rect 33416 38292 33468 38301
rect 38752 38335 38804 38344
rect 38752 38301 38761 38335
rect 38761 38301 38795 38335
rect 38795 38301 38804 38335
rect 38752 38292 38804 38301
rect 39028 38360 39080 38412
rect 40224 38360 40276 38412
rect 41236 38360 41288 38412
rect 49240 38360 49292 38412
rect 52644 38403 52696 38412
rect 52644 38369 52650 38403
rect 52650 38369 52696 38403
rect 52644 38360 52696 38369
rect 57888 38360 57940 38412
rect 60280 38360 60332 38412
rect 39948 38292 40000 38344
rect 40040 38292 40092 38344
rect 46020 38292 46072 38344
rect 52368 38292 52420 38344
rect 53104 38292 53156 38344
rect 58716 38292 58768 38344
rect 59728 38292 59780 38344
rect 62212 38360 62264 38412
rect 64236 38403 64288 38412
rect 64236 38369 64245 38403
rect 64245 38369 64279 38403
rect 64279 38369 64288 38403
rect 64236 38360 64288 38369
rect 60740 38292 60792 38344
rect 71688 38428 71740 38480
rect 34796 38224 34848 38276
rect 39120 38224 39172 38276
rect 39856 38267 39908 38276
rect 39856 38233 39865 38267
rect 39865 38233 39899 38267
rect 39899 38233 39908 38267
rect 39856 38224 39908 38233
rect 24676 38156 24728 38208
rect 25504 38156 25556 38208
rect 32956 38199 33008 38208
rect 32956 38165 32965 38199
rect 32965 38165 32999 38199
rect 32999 38165 33008 38199
rect 32956 38156 33008 38165
rect 38292 38156 38344 38208
rect 38844 38156 38896 38208
rect 40868 38224 40920 38276
rect 52736 38267 52788 38276
rect 52736 38233 52745 38267
rect 52745 38233 52779 38267
rect 52779 38233 52788 38267
rect 52736 38224 52788 38233
rect 72424 38505 72433 38539
rect 72433 38505 72467 38539
rect 72467 38505 72476 38539
rect 72424 38496 72476 38505
rect 76656 38539 76708 38548
rect 76656 38505 76665 38539
rect 76665 38505 76699 38539
rect 76699 38505 76708 38539
rect 76656 38496 76708 38505
rect 77116 38496 77168 38548
rect 79048 38496 79100 38548
rect 79968 38496 80020 38548
rect 83372 38496 83424 38548
rect 73528 38428 73580 38480
rect 73160 38360 73212 38412
rect 76012 38360 76064 38412
rect 79140 38428 79192 38480
rect 79692 38471 79744 38480
rect 79692 38437 79701 38471
rect 79701 38437 79735 38471
rect 79735 38437 79744 38471
rect 79692 38428 79744 38437
rect 84292 38428 84344 38480
rect 77484 38292 77536 38344
rect 78220 38292 78272 38344
rect 40040 38156 40092 38208
rect 41236 38199 41288 38208
rect 41236 38165 41245 38199
rect 41245 38165 41279 38199
rect 41279 38165 41288 38199
rect 41236 38156 41288 38165
rect 55312 38156 55364 38208
rect 60832 38199 60884 38208
rect 60832 38165 60841 38199
rect 60841 38165 60875 38199
rect 60875 38165 60884 38199
rect 60832 38156 60884 38165
rect 62212 38156 62264 38208
rect 66260 38224 66312 38276
rect 73344 38224 73396 38276
rect 79784 38360 79836 38412
rect 80336 38360 80388 38412
rect 80888 38360 80940 38412
rect 79048 38292 79100 38344
rect 84200 38335 84252 38344
rect 78956 38224 79008 38276
rect 65432 38199 65484 38208
rect 65432 38165 65441 38199
rect 65441 38165 65475 38199
rect 65475 38165 65484 38199
rect 78772 38199 78824 38208
rect 65432 38156 65484 38165
rect 78772 38165 78781 38199
rect 78781 38165 78815 38199
rect 78815 38165 78824 38199
rect 79416 38224 79468 38276
rect 84200 38301 84209 38335
rect 84209 38301 84243 38335
rect 84243 38301 84252 38335
rect 84200 38292 84252 38301
rect 85396 38224 85448 38276
rect 78772 38156 78824 38165
rect 79968 38156 80020 38208
rect 83372 38156 83424 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 65686 38054 65738 38106
rect 65750 38054 65802 38106
rect 65814 38054 65866 38106
rect 65878 38054 65930 38106
rect 96406 38054 96458 38106
rect 96470 38054 96522 38106
rect 96534 38054 96586 38106
rect 96598 38054 96650 38106
rect 4620 37952 4672 38004
rect 4712 37995 4764 38004
rect 4712 37961 4721 37995
rect 4721 37961 4755 37995
rect 4755 37961 4764 37995
rect 4712 37952 4764 37961
rect 5080 37995 5132 38004
rect 5080 37961 5089 37995
rect 5089 37961 5123 37995
rect 5123 37961 5132 37995
rect 5080 37952 5132 37961
rect 11060 37952 11112 38004
rect 22192 37995 22244 38004
rect 22192 37961 22201 37995
rect 22201 37961 22235 37995
rect 22235 37961 22244 37995
rect 22192 37952 22244 37961
rect 51724 37952 51776 38004
rect 54576 37952 54628 38004
rect 58716 37952 58768 38004
rect 58900 37995 58952 38004
rect 58900 37961 58909 37995
rect 58909 37961 58943 37995
rect 58943 37961 58952 37995
rect 58900 37952 58952 37961
rect 60832 37952 60884 38004
rect 70124 37952 70176 38004
rect 72332 37952 72384 38004
rect 73068 37952 73120 38004
rect 77484 37995 77536 38004
rect 77484 37961 77493 37995
rect 77493 37961 77527 37995
rect 77527 37961 77536 37995
rect 77484 37952 77536 37961
rect 77760 37995 77812 38004
rect 77760 37961 77769 37995
rect 77769 37961 77803 37995
rect 77803 37961 77812 37995
rect 77760 37952 77812 37961
rect 86776 37952 86828 38004
rect 3424 37748 3476 37800
rect 15844 37884 15896 37936
rect 21732 37927 21784 37936
rect 21732 37893 21741 37927
rect 21741 37893 21775 37927
rect 21775 37893 21784 37927
rect 21732 37884 21784 37893
rect 22652 37884 22704 37936
rect 27620 37884 27672 37936
rect 10968 37816 11020 37868
rect 12532 37859 12584 37868
rect 12532 37825 12541 37859
rect 12541 37825 12575 37859
rect 12575 37825 12584 37859
rect 12532 37816 12584 37825
rect 16028 37816 16080 37868
rect 5080 37748 5132 37800
rect 5632 37791 5684 37800
rect 5632 37757 5641 37791
rect 5641 37757 5675 37791
rect 5675 37757 5684 37791
rect 5632 37748 5684 37757
rect 5724 37723 5776 37732
rect 5724 37689 5733 37723
rect 5733 37689 5767 37723
rect 5767 37689 5776 37723
rect 5724 37680 5776 37689
rect 3792 37612 3844 37664
rect 10232 37791 10284 37800
rect 10232 37757 10241 37791
rect 10241 37757 10275 37791
rect 10275 37757 10284 37791
rect 10232 37748 10284 37757
rect 12440 37791 12492 37800
rect 12440 37757 12449 37791
rect 12449 37757 12483 37791
rect 12483 37757 12492 37791
rect 12440 37748 12492 37757
rect 20720 37748 20772 37800
rect 23664 37816 23716 37868
rect 25504 37859 25556 37868
rect 25504 37825 25513 37859
rect 25513 37825 25547 37859
rect 25547 37825 25556 37859
rect 25504 37816 25556 37825
rect 25596 37816 25648 37868
rect 21364 37791 21416 37800
rect 21364 37757 21373 37791
rect 21373 37757 21407 37791
rect 21407 37757 21416 37791
rect 21364 37748 21416 37757
rect 22192 37748 22244 37800
rect 10508 37680 10560 37732
rect 23756 37723 23808 37732
rect 23756 37689 23765 37723
rect 23765 37689 23799 37723
rect 23799 37689 23808 37723
rect 23756 37680 23808 37689
rect 17316 37612 17368 37664
rect 17868 37612 17920 37664
rect 20076 37612 20128 37664
rect 21364 37612 21416 37664
rect 26148 37791 26200 37800
rect 26148 37757 26157 37791
rect 26157 37757 26191 37791
rect 26191 37757 26200 37791
rect 26148 37748 26200 37757
rect 27712 37748 27764 37800
rect 36360 37816 36412 37868
rect 34612 37748 34664 37800
rect 34796 37748 34848 37800
rect 36636 37884 36688 37936
rect 37280 37816 37332 37868
rect 39856 37816 39908 37868
rect 51448 37884 51500 37936
rect 52368 37884 52420 37936
rect 58624 37884 58676 37936
rect 46572 37748 46624 37800
rect 52000 37748 52052 37800
rect 52368 37791 52420 37800
rect 52368 37757 52377 37791
rect 52377 37757 52411 37791
rect 52411 37757 52420 37791
rect 52368 37748 52420 37757
rect 52552 37748 52604 37800
rect 53380 37816 53432 37868
rect 85580 37884 85632 37936
rect 53564 37748 53616 37800
rect 55036 37748 55088 37800
rect 27160 37680 27212 37732
rect 38844 37723 38896 37732
rect 26148 37612 26200 37664
rect 32312 37612 32364 37664
rect 32956 37655 33008 37664
rect 32956 37621 32965 37655
rect 32965 37621 32999 37655
rect 32999 37621 33008 37655
rect 32956 37612 33008 37621
rect 33692 37655 33744 37664
rect 33692 37621 33701 37655
rect 33701 37621 33735 37655
rect 33735 37621 33744 37655
rect 33692 37612 33744 37621
rect 34980 37655 35032 37664
rect 34980 37621 34989 37655
rect 34989 37621 35023 37655
rect 35023 37621 35032 37655
rect 34980 37612 35032 37621
rect 38844 37689 38853 37723
rect 38853 37689 38887 37723
rect 38887 37689 38896 37723
rect 38844 37680 38896 37689
rect 46020 37680 46072 37732
rect 56508 37680 56560 37732
rect 61016 37748 61068 37800
rect 63316 37748 63368 37800
rect 64696 37816 64748 37868
rect 79876 37816 79928 37868
rect 64880 37748 64932 37800
rect 65156 37791 65208 37800
rect 65156 37757 65165 37791
rect 65165 37757 65199 37791
rect 65199 37757 65208 37791
rect 65156 37748 65208 37757
rect 65524 37791 65576 37800
rect 65524 37757 65533 37791
rect 65533 37757 65567 37791
rect 65567 37757 65576 37791
rect 65524 37748 65576 37757
rect 72332 37791 72384 37800
rect 72332 37757 72341 37791
rect 72341 37757 72375 37791
rect 72375 37757 72384 37791
rect 72332 37748 72384 37757
rect 65064 37680 65116 37732
rect 66444 37680 66496 37732
rect 68560 37680 68612 37732
rect 73160 37748 73212 37800
rect 77760 37748 77812 37800
rect 79784 37791 79836 37800
rect 79784 37757 79793 37791
rect 79793 37757 79827 37791
rect 79827 37757 79836 37791
rect 79784 37748 79836 37757
rect 79968 37791 80020 37800
rect 79968 37757 79977 37791
rect 79977 37757 80011 37791
rect 80011 37757 80020 37791
rect 79968 37748 80020 37757
rect 86592 37791 86644 37800
rect 86592 37757 86601 37791
rect 86601 37757 86635 37791
rect 86635 37757 86644 37791
rect 86592 37748 86644 37757
rect 79324 37680 79376 37732
rect 80336 37723 80388 37732
rect 46204 37655 46256 37664
rect 46204 37621 46213 37655
rect 46213 37621 46247 37655
rect 46247 37621 46256 37655
rect 46204 37612 46256 37621
rect 52000 37612 52052 37664
rect 53564 37612 53616 37664
rect 60188 37612 60240 37664
rect 60924 37655 60976 37664
rect 60924 37621 60933 37655
rect 60933 37621 60967 37655
rect 60967 37621 60976 37655
rect 60924 37612 60976 37621
rect 63132 37612 63184 37664
rect 63316 37655 63368 37664
rect 63316 37621 63325 37655
rect 63325 37621 63359 37655
rect 63359 37621 63368 37655
rect 63316 37612 63368 37621
rect 64696 37612 64748 37664
rect 66168 37612 66220 37664
rect 72516 37655 72568 37664
rect 72516 37621 72525 37655
rect 72525 37621 72559 37655
rect 72559 37621 72568 37655
rect 72516 37612 72568 37621
rect 72608 37612 72660 37664
rect 79416 37612 79468 37664
rect 80336 37689 80345 37723
rect 80345 37689 80379 37723
rect 80379 37689 80388 37723
rect 80336 37680 80388 37689
rect 84200 37612 84252 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 81046 37510 81098 37562
rect 81110 37510 81162 37562
rect 81174 37510 81226 37562
rect 81238 37510 81290 37562
rect 4804 37408 4856 37460
rect 5632 37408 5684 37460
rect 10968 37451 11020 37460
rect 10968 37417 10977 37451
rect 10977 37417 11011 37451
rect 11011 37417 11020 37451
rect 10968 37408 11020 37417
rect 11060 37408 11112 37460
rect 6000 37340 6052 37392
rect 5724 37272 5776 37324
rect 10324 37315 10376 37324
rect 4804 37204 4856 37256
rect 9680 37247 9732 37256
rect 9680 37213 9689 37247
rect 9689 37213 9723 37247
rect 9723 37213 9732 37247
rect 9680 37204 9732 37213
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 10876 37315 10928 37324
rect 10508 37204 10560 37256
rect 10876 37281 10885 37315
rect 10885 37281 10919 37315
rect 10919 37281 10928 37315
rect 10876 37272 10928 37281
rect 11060 37204 11112 37256
rect 15568 37272 15620 37324
rect 16120 37272 16172 37324
rect 17132 37272 17184 37324
rect 20812 37272 20864 37324
rect 30380 37408 30432 37460
rect 32864 37408 32916 37460
rect 22192 37340 22244 37392
rect 21456 37272 21508 37324
rect 22744 37340 22796 37392
rect 63316 37408 63368 37460
rect 66076 37408 66128 37460
rect 66260 37451 66312 37460
rect 66260 37417 66269 37451
rect 66269 37417 66303 37451
rect 66303 37417 66312 37451
rect 66260 37408 66312 37417
rect 71688 37408 71740 37460
rect 73620 37408 73672 37460
rect 78956 37451 79008 37460
rect 78956 37417 78965 37451
rect 78965 37417 78999 37451
rect 78999 37417 79008 37451
rect 78956 37408 79008 37417
rect 33416 37383 33468 37392
rect 33416 37349 33425 37383
rect 33425 37349 33459 37383
rect 33459 37349 33468 37383
rect 33416 37340 33468 37349
rect 21824 37204 21876 37256
rect 22376 37315 22428 37324
rect 22376 37281 22385 37315
rect 22385 37281 22419 37315
rect 22419 37281 22428 37315
rect 27160 37315 27212 37324
rect 22376 37272 22428 37281
rect 27160 37281 27169 37315
rect 27169 37281 27203 37315
rect 27203 37281 27212 37315
rect 27160 37272 27212 37281
rect 32956 37272 33008 37324
rect 33048 37315 33100 37324
rect 33048 37281 33057 37315
rect 33057 37281 33091 37315
rect 33091 37281 33100 37315
rect 34980 37340 35032 37392
rect 38292 37383 38344 37392
rect 38292 37349 38301 37383
rect 38301 37349 38335 37383
rect 38335 37349 38344 37383
rect 38292 37340 38344 37349
rect 46572 37383 46624 37392
rect 46572 37349 46581 37383
rect 46581 37349 46615 37383
rect 46615 37349 46624 37383
rect 46572 37340 46624 37349
rect 46664 37340 46716 37392
rect 50988 37340 51040 37392
rect 53104 37383 53156 37392
rect 53104 37349 53113 37383
rect 53113 37349 53147 37383
rect 53147 37349 53156 37383
rect 53104 37340 53156 37349
rect 53380 37383 53432 37392
rect 53380 37349 53389 37383
rect 53389 37349 53423 37383
rect 53423 37349 53432 37383
rect 53380 37340 53432 37349
rect 53564 37383 53616 37392
rect 53564 37349 53573 37383
rect 53573 37349 53607 37383
rect 53607 37349 53616 37383
rect 53564 37340 53616 37349
rect 59728 37340 59780 37392
rect 63132 37340 63184 37392
rect 34336 37315 34388 37324
rect 33048 37272 33100 37281
rect 34336 37281 34345 37315
rect 34345 37281 34379 37315
rect 34379 37281 34388 37315
rect 34336 37272 34388 37281
rect 26792 37204 26844 37256
rect 27896 37204 27948 37256
rect 4068 37068 4120 37120
rect 7932 37068 7984 37120
rect 14280 37068 14332 37120
rect 32956 37136 33008 37188
rect 38476 37247 38528 37256
rect 38476 37213 38485 37247
rect 38485 37213 38519 37247
rect 38519 37213 38528 37247
rect 38476 37204 38528 37213
rect 38752 37247 38804 37256
rect 38752 37213 38761 37247
rect 38761 37213 38795 37247
rect 38795 37213 38804 37247
rect 38752 37204 38804 37213
rect 40960 37315 41012 37324
rect 40960 37281 40969 37315
rect 40969 37281 41003 37315
rect 41003 37281 41012 37315
rect 40960 37272 41012 37281
rect 44548 37315 44600 37324
rect 44548 37281 44557 37315
rect 44557 37281 44591 37315
rect 44591 37281 44600 37315
rect 44548 37272 44600 37281
rect 44824 37315 44876 37324
rect 44824 37281 44841 37315
rect 44841 37281 44875 37315
rect 44875 37281 44876 37315
rect 51816 37315 51868 37324
rect 44824 37272 44876 37281
rect 51816 37281 51825 37315
rect 51825 37281 51859 37315
rect 51859 37281 51868 37315
rect 51816 37272 51868 37281
rect 52000 37315 52052 37324
rect 52000 37281 52009 37315
rect 52009 37281 52043 37315
rect 52043 37281 52052 37315
rect 52000 37272 52052 37281
rect 52552 37315 52604 37324
rect 52552 37281 52561 37315
rect 52561 37281 52595 37315
rect 52595 37281 52604 37315
rect 52552 37272 52604 37281
rect 60188 37315 60240 37324
rect 60188 37281 60197 37315
rect 60197 37281 60231 37315
rect 60231 37281 60240 37315
rect 60188 37272 60240 37281
rect 64604 37272 64656 37324
rect 42156 37204 42208 37256
rect 44916 37247 44968 37256
rect 44916 37213 44925 37247
rect 44925 37213 44959 37247
rect 44959 37213 44968 37247
rect 44916 37204 44968 37213
rect 45192 37247 45244 37256
rect 45192 37213 45201 37247
rect 45201 37213 45235 37247
rect 45235 37213 45244 37247
rect 45192 37204 45244 37213
rect 53104 37204 53156 37256
rect 65340 37272 65392 37324
rect 66996 37340 67048 37392
rect 32220 37068 32272 37120
rect 32772 37068 32824 37120
rect 34336 37068 34388 37120
rect 38384 37068 38436 37120
rect 38936 37068 38988 37120
rect 44732 37068 44784 37120
rect 46756 37111 46808 37120
rect 46756 37077 46765 37111
rect 46765 37077 46799 37111
rect 46799 37077 46808 37111
rect 46756 37068 46808 37077
rect 63224 37068 63276 37120
rect 65248 37204 65300 37256
rect 65984 37272 66036 37324
rect 78772 37340 78824 37392
rect 79324 37383 79376 37392
rect 70124 37315 70176 37324
rect 70124 37281 70133 37315
rect 70133 37281 70167 37315
rect 70167 37281 70176 37315
rect 70124 37272 70176 37281
rect 71136 37272 71188 37324
rect 72516 37272 72568 37324
rect 73160 37272 73212 37324
rect 77208 37272 77260 37324
rect 79324 37349 79333 37383
rect 79333 37349 79367 37383
rect 79367 37349 79376 37383
rect 79324 37340 79376 37349
rect 80888 37383 80940 37392
rect 80888 37349 80897 37383
rect 80897 37349 80931 37383
rect 80931 37349 80940 37383
rect 80888 37340 80940 37349
rect 79876 37272 79928 37324
rect 79692 37247 79744 37256
rect 79692 37213 79701 37247
rect 79701 37213 79735 37247
rect 79735 37213 79744 37247
rect 79692 37204 79744 37213
rect 79784 37204 79836 37256
rect 81348 37272 81400 37324
rect 84200 37408 84252 37460
rect 85580 37383 85632 37392
rect 85580 37349 85589 37383
rect 85589 37349 85623 37383
rect 85623 37349 85632 37383
rect 85580 37340 85632 37349
rect 85856 37272 85908 37324
rect 85948 37315 86000 37324
rect 85948 37281 85957 37315
rect 85957 37281 85991 37315
rect 85991 37281 86000 37315
rect 85948 37272 86000 37281
rect 85764 37247 85816 37256
rect 85764 37213 85773 37247
rect 85773 37213 85807 37247
rect 85807 37213 85816 37247
rect 87328 37272 87380 37324
rect 85764 37204 85816 37213
rect 64880 37136 64932 37188
rect 78956 37136 79008 37188
rect 65248 37111 65300 37120
rect 65248 37077 65257 37111
rect 65257 37077 65291 37111
rect 65291 37077 65300 37111
rect 65248 37068 65300 37077
rect 79968 37111 80020 37120
rect 79968 37077 79977 37111
rect 79977 37077 80011 37111
rect 80011 37077 80020 37111
rect 79968 37068 80020 37077
rect 80428 37068 80480 37120
rect 88432 37068 88484 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 65686 36966 65738 37018
rect 65750 36966 65802 37018
rect 65814 36966 65866 37018
rect 65878 36966 65930 37018
rect 96406 36966 96458 37018
rect 96470 36966 96522 37018
rect 96534 36966 96586 37018
rect 96598 36966 96650 37018
rect 4804 36796 4856 36848
rect 3332 36524 3384 36576
rect 3792 36660 3844 36712
rect 5724 36864 5776 36916
rect 9864 36864 9916 36916
rect 9956 36907 10008 36916
rect 9956 36873 9965 36907
rect 9965 36873 9999 36907
rect 9999 36873 10008 36907
rect 9956 36864 10008 36873
rect 11060 36864 11112 36916
rect 19248 36864 19300 36916
rect 5540 36796 5592 36848
rect 16396 36796 16448 36848
rect 16672 36839 16724 36848
rect 16672 36805 16681 36839
rect 16681 36805 16715 36839
rect 16715 36805 16724 36839
rect 16672 36796 16724 36805
rect 9128 36771 9180 36780
rect 9128 36737 9137 36771
rect 9137 36737 9171 36771
rect 9171 36737 9180 36771
rect 9128 36728 9180 36737
rect 9956 36728 10008 36780
rect 16580 36728 16632 36780
rect 25504 36796 25556 36848
rect 26240 36796 26292 36848
rect 26332 36839 26384 36848
rect 26332 36805 26341 36839
rect 26341 36805 26375 36839
rect 26375 36805 26384 36839
rect 33324 36864 33376 36916
rect 38752 36864 38804 36916
rect 47860 36864 47912 36916
rect 50712 36907 50764 36916
rect 50712 36873 50721 36907
rect 50721 36873 50755 36907
rect 50755 36873 50764 36907
rect 50712 36864 50764 36873
rect 26332 36796 26384 36805
rect 6920 36592 6972 36644
rect 9864 36660 9916 36712
rect 13544 36703 13596 36712
rect 13544 36669 13553 36703
rect 13553 36669 13587 36703
rect 13587 36669 13596 36703
rect 13544 36660 13596 36669
rect 14280 36703 14332 36712
rect 14280 36669 14289 36703
rect 14289 36669 14323 36703
rect 14323 36669 14332 36703
rect 14280 36660 14332 36669
rect 15292 36660 15344 36712
rect 19248 36660 19300 36712
rect 21456 36703 21508 36712
rect 21456 36669 21465 36703
rect 21465 36669 21499 36703
rect 21499 36669 21508 36703
rect 21456 36660 21508 36669
rect 21824 36703 21876 36712
rect 21824 36669 21833 36703
rect 21833 36669 21867 36703
rect 21867 36669 21876 36703
rect 21824 36660 21876 36669
rect 9772 36592 9824 36644
rect 16672 36592 16724 36644
rect 5080 36524 5132 36576
rect 13636 36567 13688 36576
rect 13636 36533 13645 36567
rect 13645 36533 13679 36567
rect 13679 36533 13688 36567
rect 13636 36524 13688 36533
rect 16028 36567 16080 36576
rect 16028 36533 16037 36567
rect 16037 36533 16071 36567
rect 16071 36533 16080 36567
rect 16028 36524 16080 36533
rect 24768 36524 24820 36576
rect 26608 36660 26660 36712
rect 32680 36703 32732 36712
rect 26056 36635 26108 36644
rect 26056 36601 26065 36635
rect 26065 36601 26099 36635
rect 26099 36601 26108 36635
rect 26056 36592 26108 36601
rect 26332 36592 26384 36644
rect 30380 36592 30432 36644
rect 32680 36669 32689 36703
rect 32689 36669 32723 36703
rect 32723 36669 32732 36703
rect 32680 36660 32732 36669
rect 33232 36660 33284 36712
rect 33692 36660 33744 36712
rect 32220 36592 32272 36644
rect 32588 36592 32640 36644
rect 37096 36592 37148 36644
rect 37648 36703 37700 36712
rect 37648 36669 37657 36703
rect 37657 36669 37691 36703
rect 37691 36669 37700 36703
rect 37648 36660 37700 36669
rect 38108 36660 38160 36712
rect 38384 36703 38436 36712
rect 38384 36669 38393 36703
rect 38393 36669 38427 36703
rect 38427 36669 38436 36703
rect 38384 36660 38436 36669
rect 37740 36592 37792 36644
rect 42156 36703 42208 36712
rect 42156 36669 42165 36703
rect 42165 36669 42199 36703
rect 42199 36669 42208 36703
rect 42156 36660 42208 36669
rect 48136 36796 48188 36848
rect 51356 36796 51408 36848
rect 51724 36796 51776 36848
rect 50804 36728 50856 36780
rect 59912 36864 59964 36916
rect 60924 36864 60976 36916
rect 64880 36864 64932 36916
rect 65248 36864 65300 36916
rect 65340 36839 65392 36848
rect 65340 36805 65349 36839
rect 65349 36805 65383 36839
rect 65383 36805 65392 36839
rect 65340 36796 65392 36805
rect 66076 36839 66128 36848
rect 66076 36805 66085 36839
rect 66085 36805 66119 36839
rect 66119 36805 66128 36839
rect 66076 36796 66128 36805
rect 78772 36907 78824 36916
rect 78772 36873 78781 36907
rect 78781 36873 78815 36907
rect 78815 36873 78824 36907
rect 78772 36864 78824 36873
rect 79140 36864 79192 36916
rect 79876 36864 79928 36916
rect 84752 36907 84804 36916
rect 84752 36873 84761 36907
rect 84761 36873 84795 36907
rect 84795 36873 84804 36907
rect 84752 36864 84804 36873
rect 85396 36864 85448 36916
rect 85948 36907 86000 36916
rect 46756 36660 46808 36712
rect 43720 36592 43772 36644
rect 51724 36703 51776 36712
rect 51724 36669 51733 36703
rect 51733 36669 51767 36703
rect 51767 36669 51776 36703
rect 51724 36660 51776 36669
rect 58440 36703 58492 36712
rect 25872 36567 25924 36576
rect 25872 36533 25881 36567
rect 25881 36533 25915 36567
rect 25915 36533 25924 36567
rect 25872 36524 25924 36533
rect 36636 36524 36688 36576
rect 37372 36567 37424 36576
rect 37372 36533 37381 36567
rect 37381 36533 37415 36567
rect 37415 36533 37424 36567
rect 37372 36524 37424 36533
rect 48504 36567 48556 36576
rect 48504 36533 48513 36567
rect 48513 36533 48547 36567
rect 48547 36533 48556 36567
rect 48504 36524 48556 36533
rect 52368 36524 52420 36576
rect 53104 36567 53156 36576
rect 53104 36533 53113 36567
rect 53113 36533 53147 36567
rect 53147 36533 53156 36567
rect 53104 36524 53156 36533
rect 58440 36669 58449 36703
rect 58449 36669 58483 36703
rect 58483 36669 58492 36703
rect 58440 36660 58492 36669
rect 62028 36728 62080 36780
rect 64420 36703 64472 36712
rect 63132 36592 63184 36644
rect 59912 36567 59964 36576
rect 59912 36533 59921 36567
rect 59921 36533 59955 36567
rect 59955 36533 59964 36567
rect 59912 36524 59964 36533
rect 64420 36669 64429 36703
rect 64429 36669 64463 36703
rect 64463 36669 64472 36703
rect 64420 36660 64472 36669
rect 64604 36703 64656 36712
rect 64604 36669 64613 36703
rect 64613 36669 64647 36703
rect 64647 36669 64656 36703
rect 64604 36660 64656 36669
rect 65248 36660 65300 36712
rect 66444 36771 66496 36780
rect 66444 36737 66453 36771
rect 66453 36737 66487 36771
rect 66487 36737 66496 36771
rect 66444 36728 66496 36737
rect 71136 36771 71188 36780
rect 71136 36737 71145 36771
rect 71145 36737 71179 36771
rect 71179 36737 71188 36771
rect 71136 36728 71188 36737
rect 65984 36703 66036 36712
rect 65984 36669 65993 36703
rect 65993 36669 66027 36703
rect 66027 36669 66036 36703
rect 65984 36660 66036 36669
rect 66168 36660 66220 36712
rect 75920 36703 75972 36712
rect 65432 36592 65484 36644
rect 68652 36592 68704 36644
rect 68100 36524 68152 36576
rect 72424 36567 72476 36576
rect 72424 36533 72433 36567
rect 72433 36533 72467 36567
rect 72467 36533 72476 36567
rect 72424 36524 72476 36533
rect 75920 36669 75929 36703
rect 75929 36669 75963 36703
rect 75963 36669 75972 36703
rect 75920 36660 75972 36669
rect 79784 36796 79836 36848
rect 79968 36796 80020 36848
rect 85488 36796 85540 36848
rect 80336 36728 80388 36780
rect 85948 36873 85957 36907
rect 85957 36873 85991 36907
rect 85991 36873 86000 36907
rect 85948 36864 86000 36873
rect 86592 36864 86644 36916
rect 86776 36864 86828 36916
rect 81440 36703 81492 36712
rect 72792 36592 72844 36644
rect 73344 36524 73396 36576
rect 75000 36524 75052 36576
rect 79692 36592 79744 36644
rect 81440 36669 81449 36703
rect 81449 36669 81483 36703
rect 81483 36669 81492 36703
rect 81440 36660 81492 36669
rect 84108 36524 84160 36576
rect 86960 36660 87012 36712
rect 87880 36592 87932 36644
rect 88432 36703 88484 36712
rect 88432 36669 88441 36703
rect 88441 36669 88475 36703
rect 88475 36669 88484 36703
rect 88432 36660 88484 36669
rect 88340 36635 88392 36644
rect 88340 36601 88349 36635
rect 88349 36601 88383 36635
rect 88383 36601 88392 36635
rect 88340 36592 88392 36601
rect 88708 36592 88760 36644
rect 85304 36524 85356 36576
rect 87972 36567 88024 36576
rect 87972 36533 87981 36567
rect 87981 36533 88015 36567
rect 88015 36533 88024 36567
rect 87972 36524 88024 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 81046 36422 81098 36474
rect 81110 36422 81162 36474
rect 81174 36422 81226 36474
rect 81238 36422 81290 36474
rect 4804 36320 4856 36372
rect 16672 36320 16724 36372
rect 17132 36363 17184 36372
rect 17132 36329 17141 36363
rect 17141 36329 17175 36363
rect 17175 36329 17184 36363
rect 17132 36320 17184 36329
rect 18420 36320 18472 36372
rect 24492 36320 24544 36372
rect 3240 36252 3292 36304
rect 26884 36252 26936 36304
rect 5264 36227 5316 36236
rect 5264 36193 5273 36227
rect 5273 36193 5307 36227
rect 5307 36193 5316 36227
rect 5264 36184 5316 36193
rect 9680 36184 9732 36236
rect 15292 36227 15344 36236
rect 15292 36193 15301 36227
rect 15301 36193 15335 36227
rect 15335 36193 15344 36227
rect 15292 36184 15344 36193
rect 15200 36116 15252 36168
rect 16212 36184 16264 36236
rect 17500 36184 17552 36236
rect 19892 36184 19944 36236
rect 21456 36184 21508 36236
rect 21916 36227 21968 36236
rect 16672 36116 16724 36168
rect 19340 36116 19392 36168
rect 9772 36048 9824 36100
rect 10324 36048 10376 36100
rect 21916 36193 21925 36227
rect 21925 36193 21959 36227
rect 21959 36193 21968 36227
rect 21916 36184 21968 36193
rect 22284 36184 22336 36236
rect 26332 36184 26384 36236
rect 26516 36227 26568 36236
rect 26516 36193 26525 36227
rect 26525 36193 26559 36227
rect 26559 36193 26568 36227
rect 26516 36184 26568 36193
rect 33140 36184 33192 36236
rect 37280 36252 37332 36304
rect 34152 36184 34204 36236
rect 37648 36320 37700 36372
rect 68560 36363 68612 36372
rect 47860 36295 47912 36304
rect 37740 36227 37792 36236
rect 37740 36193 37749 36227
rect 37749 36193 37783 36227
rect 37783 36193 37792 36227
rect 37740 36184 37792 36193
rect 15200 35980 15252 36032
rect 17500 36023 17552 36032
rect 17500 35989 17509 36023
rect 17509 35989 17543 36023
rect 17543 35989 17552 36023
rect 17500 35980 17552 35989
rect 24492 36116 24544 36168
rect 38108 36184 38160 36236
rect 47860 36261 47869 36295
rect 47869 36261 47903 36295
rect 47903 36261 47912 36295
rect 47860 36252 47912 36261
rect 48136 36295 48188 36304
rect 48136 36261 48145 36295
rect 48145 36261 48179 36295
rect 48179 36261 48188 36295
rect 48136 36252 48188 36261
rect 52368 36252 52420 36304
rect 32588 36048 32640 36100
rect 33232 36048 33284 36100
rect 22284 35980 22336 36032
rect 25504 35980 25556 36032
rect 25872 35980 25924 36032
rect 26424 35980 26476 36032
rect 32680 35980 32732 36032
rect 38292 36048 38344 36100
rect 44916 36116 44968 36168
rect 51356 36184 51408 36236
rect 68560 36329 68569 36363
rect 68569 36329 68603 36363
rect 68603 36329 68612 36363
rect 68560 36320 68612 36329
rect 68652 36320 68704 36372
rect 57704 36184 57756 36236
rect 64420 36252 64472 36304
rect 66996 36295 67048 36304
rect 66996 36261 67005 36295
rect 67005 36261 67039 36295
rect 67039 36261 67048 36295
rect 66996 36252 67048 36261
rect 62028 36184 62080 36236
rect 67640 36227 67692 36236
rect 67640 36193 67649 36227
rect 67649 36193 67683 36227
rect 67683 36193 67692 36227
rect 67640 36184 67692 36193
rect 68008 36227 68060 36236
rect 68008 36193 68017 36227
rect 68017 36193 68051 36227
rect 68051 36193 68060 36227
rect 68008 36184 68060 36193
rect 34152 36023 34204 36032
rect 34152 35989 34161 36023
rect 34161 35989 34195 36023
rect 34195 35989 34204 36023
rect 34152 35980 34204 35989
rect 38384 35980 38436 36032
rect 47032 36048 47084 36100
rect 46756 36023 46808 36032
rect 46756 35989 46765 36023
rect 46765 35989 46799 36023
rect 46799 35989 46808 36023
rect 46756 35980 46808 35989
rect 48504 35980 48556 36032
rect 50988 36116 51040 36168
rect 56968 36116 57020 36168
rect 67732 36159 67784 36168
rect 67732 36125 67741 36159
rect 67741 36125 67775 36159
rect 67775 36125 67784 36159
rect 67732 36116 67784 36125
rect 67916 36159 67968 36168
rect 67916 36125 67925 36159
rect 67925 36125 67959 36159
rect 67959 36125 67968 36159
rect 67916 36116 67968 36125
rect 58072 36023 58124 36032
rect 58072 35989 58081 36023
rect 58081 35989 58115 36023
rect 58115 35989 58124 36023
rect 58072 35980 58124 35989
rect 62764 35980 62816 36032
rect 68652 35980 68704 36032
rect 73344 36184 73396 36236
rect 76012 36320 76064 36372
rect 85948 36320 86000 36372
rect 86868 36320 86920 36372
rect 71964 36116 72016 36168
rect 75184 36184 75236 36236
rect 75368 36227 75420 36236
rect 75368 36193 75377 36227
rect 75377 36193 75411 36227
rect 75411 36193 75420 36227
rect 75368 36184 75420 36193
rect 79876 36184 79928 36236
rect 80428 36184 80480 36236
rect 85856 36252 85908 36304
rect 86776 36295 86828 36304
rect 86776 36261 86785 36295
rect 86785 36261 86819 36295
rect 86819 36261 86828 36295
rect 86776 36252 86828 36261
rect 87328 36295 87380 36304
rect 87328 36261 87337 36295
rect 87337 36261 87371 36295
rect 87371 36261 87380 36295
rect 87328 36252 87380 36261
rect 88708 36227 88760 36236
rect 75828 36159 75880 36168
rect 75828 36125 75837 36159
rect 75837 36125 75871 36159
rect 75871 36125 75880 36159
rect 75828 36116 75880 36125
rect 88064 36116 88116 36168
rect 77208 36048 77260 36100
rect 72884 36023 72936 36032
rect 72884 35989 72893 36023
rect 72893 35989 72927 36023
rect 72927 35989 72936 36023
rect 72884 35980 72936 35989
rect 73344 36023 73396 36032
rect 73344 35989 73353 36023
rect 73353 35989 73387 36023
rect 73387 35989 73396 36023
rect 73344 35980 73396 35989
rect 76656 35980 76708 36032
rect 79508 35980 79560 36032
rect 80244 36023 80296 36032
rect 80244 35989 80253 36023
rect 80253 35989 80287 36023
rect 80287 35989 80296 36023
rect 80244 35980 80296 35989
rect 85764 36048 85816 36100
rect 87972 36048 88024 36100
rect 86316 35980 86368 36032
rect 88708 36193 88717 36227
rect 88717 36193 88751 36227
rect 88751 36193 88760 36227
rect 88708 36184 88760 36193
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 65686 35878 65738 35930
rect 65750 35878 65802 35930
rect 65814 35878 65866 35930
rect 65878 35878 65930 35930
rect 96406 35878 96458 35930
rect 96470 35878 96522 35930
rect 96534 35878 96586 35930
rect 96598 35878 96650 35930
rect 4068 35776 4120 35828
rect 17776 35776 17828 35828
rect 17868 35776 17920 35828
rect 20628 35776 20680 35828
rect 21916 35776 21968 35828
rect 26056 35776 26108 35828
rect 26700 35776 26752 35828
rect 38292 35776 38344 35828
rect 38384 35776 38436 35828
rect 62764 35776 62816 35828
rect 65984 35776 66036 35828
rect 66812 35776 66864 35828
rect 68008 35776 68060 35828
rect 71688 35776 71740 35828
rect 75920 35776 75972 35828
rect 77024 35776 77076 35828
rect 81348 35819 81400 35828
rect 81348 35785 81357 35819
rect 81357 35785 81391 35819
rect 81391 35785 81400 35819
rect 81348 35776 81400 35785
rect 6000 35751 6052 35760
rect 6000 35717 6009 35751
rect 6009 35717 6043 35751
rect 6043 35717 6052 35751
rect 6000 35708 6052 35717
rect 9404 35708 9456 35760
rect 27620 35708 27672 35760
rect 29368 35708 29420 35760
rect 2596 35683 2648 35692
rect 2596 35649 2605 35683
rect 2605 35649 2639 35683
rect 2639 35649 2648 35683
rect 2596 35640 2648 35649
rect 3056 35640 3108 35692
rect 4896 35640 4948 35692
rect 5264 35640 5316 35692
rect 4712 35572 4764 35624
rect 13636 35640 13688 35692
rect 9312 35572 9364 35624
rect 13544 35572 13596 35624
rect 16028 35640 16080 35692
rect 21088 35640 21140 35692
rect 21824 35640 21876 35692
rect 31944 35640 31996 35692
rect 16120 35615 16172 35624
rect 3148 35436 3200 35488
rect 4160 35479 4212 35488
rect 4160 35445 4169 35479
rect 4169 35445 4203 35479
rect 4203 35445 4212 35479
rect 4160 35436 4212 35445
rect 7288 35436 7340 35488
rect 12716 35504 12768 35556
rect 15200 35547 15252 35556
rect 15200 35513 15209 35547
rect 15209 35513 15243 35547
rect 15243 35513 15252 35547
rect 16120 35581 16129 35615
rect 16129 35581 16163 35615
rect 16163 35581 16172 35615
rect 16120 35572 16172 35581
rect 15200 35504 15252 35513
rect 19892 35572 19944 35624
rect 21364 35572 21416 35624
rect 26332 35615 26384 35624
rect 26332 35581 26341 35615
rect 26341 35581 26375 35615
rect 26375 35581 26384 35615
rect 26332 35572 26384 35581
rect 26608 35572 26660 35624
rect 26884 35615 26936 35624
rect 26884 35581 26893 35615
rect 26893 35581 26927 35615
rect 26927 35581 26936 35615
rect 26884 35572 26936 35581
rect 16672 35504 16724 35556
rect 24768 35504 24820 35556
rect 26240 35504 26292 35556
rect 27068 35572 27120 35624
rect 32036 35615 32088 35624
rect 27252 35504 27304 35556
rect 32036 35581 32045 35615
rect 32045 35581 32079 35615
rect 32079 35581 32088 35615
rect 32036 35572 32088 35581
rect 32588 35572 32640 35624
rect 38844 35708 38896 35760
rect 47032 35751 47084 35760
rect 41236 35640 41288 35692
rect 34152 35615 34204 35624
rect 34152 35581 34161 35615
rect 34161 35581 34195 35615
rect 34195 35581 34204 35615
rect 34152 35572 34204 35581
rect 37372 35572 37424 35624
rect 43720 35615 43772 35624
rect 9864 35436 9916 35488
rect 13452 35479 13504 35488
rect 13452 35445 13461 35479
rect 13461 35445 13495 35479
rect 13495 35445 13504 35479
rect 13452 35436 13504 35445
rect 16488 35479 16540 35488
rect 16488 35445 16497 35479
rect 16497 35445 16531 35479
rect 16531 35445 16540 35479
rect 16488 35436 16540 35445
rect 16764 35436 16816 35488
rect 20536 35479 20588 35488
rect 20536 35445 20545 35479
rect 20545 35445 20579 35479
rect 20579 35445 20588 35479
rect 20536 35436 20588 35445
rect 20628 35436 20680 35488
rect 27068 35436 27120 35488
rect 27160 35479 27212 35488
rect 27160 35445 27169 35479
rect 27169 35445 27203 35479
rect 27203 35445 27212 35479
rect 42432 35504 42484 35556
rect 27160 35436 27212 35445
rect 28080 35436 28132 35488
rect 33508 35479 33560 35488
rect 33508 35445 33517 35479
rect 33517 35445 33551 35479
rect 33551 35445 33560 35479
rect 33508 35436 33560 35445
rect 33784 35436 33836 35488
rect 39764 35436 39816 35488
rect 43720 35581 43729 35615
rect 43729 35581 43763 35615
rect 43763 35581 43772 35615
rect 43720 35572 43772 35581
rect 47032 35717 47041 35751
rect 47041 35717 47075 35751
rect 47075 35717 47084 35751
rect 47032 35708 47084 35717
rect 51172 35708 51224 35760
rect 51908 35708 51960 35760
rect 45192 35640 45244 35692
rect 46756 35640 46808 35692
rect 46204 35572 46256 35624
rect 57060 35640 57112 35692
rect 58072 35640 58124 35692
rect 62028 35640 62080 35692
rect 53104 35572 53156 35624
rect 63132 35615 63184 35624
rect 43536 35504 43588 35556
rect 49700 35504 49752 35556
rect 56600 35504 56652 35556
rect 56876 35504 56928 35556
rect 43260 35436 43312 35488
rect 44364 35436 44416 35488
rect 63132 35581 63141 35615
rect 63141 35581 63175 35615
rect 63175 35581 63184 35615
rect 63132 35572 63184 35581
rect 67640 35640 67692 35692
rect 85488 35751 85540 35760
rect 85488 35717 85497 35751
rect 85497 35717 85531 35751
rect 85531 35717 85540 35751
rect 85488 35708 85540 35717
rect 71964 35683 72016 35692
rect 71964 35649 71973 35683
rect 71973 35649 72007 35683
rect 72007 35649 72016 35683
rect 71964 35640 72016 35649
rect 75368 35640 75420 35692
rect 75828 35683 75880 35692
rect 75828 35649 75837 35683
rect 75837 35649 75871 35683
rect 75871 35649 75880 35683
rect 75828 35640 75880 35649
rect 80244 35640 80296 35692
rect 85304 35640 85356 35692
rect 85856 35683 85908 35692
rect 59452 35436 59504 35488
rect 60924 35436 60976 35488
rect 63224 35479 63276 35488
rect 63224 35445 63233 35479
rect 63233 35445 63267 35479
rect 63267 35445 63276 35479
rect 63224 35436 63276 35445
rect 65524 35436 65576 35488
rect 66812 35615 66864 35624
rect 66812 35581 66821 35615
rect 66821 35581 66855 35615
rect 66855 35581 66864 35615
rect 66812 35572 66864 35581
rect 65984 35504 66036 35556
rect 72148 35572 72200 35624
rect 72884 35572 72936 35624
rect 74172 35547 74224 35556
rect 74172 35513 74178 35547
rect 74178 35513 74212 35547
rect 74212 35513 74224 35547
rect 74172 35504 74224 35513
rect 72148 35479 72200 35488
rect 72148 35445 72157 35479
rect 72157 35445 72191 35479
rect 72191 35445 72200 35479
rect 72148 35436 72200 35445
rect 75000 35479 75052 35488
rect 75000 35445 75009 35479
rect 75009 35445 75043 35479
rect 75043 35445 75052 35479
rect 75000 35436 75052 35445
rect 77300 35479 77352 35488
rect 77300 35445 77309 35479
rect 77309 35445 77343 35479
rect 77343 35445 77352 35479
rect 81440 35572 81492 35624
rect 85856 35649 85865 35683
rect 85865 35649 85899 35683
rect 85899 35649 85908 35683
rect 85856 35640 85908 35649
rect 88340 35683 88392 35692
rect 88340 35649 88349 35683
rect 88349 35649 88383 35683
rect 88383 35649 88392 35683
rect 88340 35640 88392 35649
rect 87880 35615 87932 35624
rect 87880 35581 87889 35615
rect 87889 35581 87923 35615
rect 87923 35581 87932 35615
rect 87880 35572 87932 35581
rect 88064 35615 88116 35624
rect 88064 35581 88073 35615
rect 88073 35581 88107 35615
rect 88107 35581 88116 35615
rect 88064 35572 88116 35581
rect 86776 35504 86828 35556
rect 77300 35436 77352 35445
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 81046 35334 81098 35386
rect 81110 35334 81162 35386
rect 81174 35334 81226 35386
rect 81238 35334 81290 35386
rect 3148 35232 3200 35284
rect 5540 35232 5592 35284
rect 3516 35164 3568 35216
rect 17316 35232 17368 35284
rect 18144 35232 18196 35284
rect 21088 35275 21140 35284
rect 21088 35241 21097 35275
rect 21097 35241 21131 35275
rect 21131 35241 21140 35275
rect 21088 35232 21140 35241
rect 21364 35275 21416 35284
rect 21364 35241 21373 35275
rect 21373 35241 21407 35275
rect 21407 35241 21416 35275
rect 21364 35232 21416 35241
rect 32496 35232 32548 35284
rect 32680 35275 32732 35284
rect 32680 35241 32689 35275
rect 32689 35241 32723 35275
rect 32723 35241 32732 35275
rect 32680 35232 32732 35241
rect 32956 35275 33008 35284
rect 32956 35241 32965 35275
rect 32965 35241 32999 35275
rect 32999 35241 33008 35275
rect 32956 35232 33008 35241
rect 26516 35207 26568 35216
rect 4896 35096 4948 35148
rect 5540 35096 5592 35148
rect 6092 35139 6144 35148
rect 6092 35105 6101 35139
rect 6101 35105 6135 35139
rect 6135 35105 6144 35139
rect 6092 35096 6144 35105
rect 6920 35096 6972 35148
rect 13912 35096 13964 35148
rect 26516 35173 26525 35207
rect 26525 35173 26559 35207
rect 26559 35173 26568 35207
rect 26516 35164 26568 35173
rect 26884 35164 26936 35216
rect 56600 35232 56652 35284
rect 58440 35232 58492 35284
rect 79508 35275 79560 35284
rect 79508 35241 79517 35275
rect 79517 35241 79551 35275
rect 79551 35241 79560 35275
rect 79508 35232 79560 35241
rect 87880 35232 87932 35284
rect 36268 35164 36320 35216
rect 21364 35096 21416 35148
rect 26608 35096 26660 35148
rect 27160 35139 27212 35148
rect 27160 35105 27169 35139
rect 27169 35105 27203 35139
rect 27203 35105 27212 35139
rect 27160 35096 27212 35105
rect 28080 35096 28132 35148
rect 31668 35096 31720 35148
rect 32404 35096 32456 35148
rect 38476 35164 38528 35216
rect 39580 35164 39632 35216
rect 39672 35164 39724 35216
rect 42616 35164 42668 35216
rect 43812 35164 43864 35216
rect 16488 35028 16540 35080
rect 26700 35028 26752 35080
rect 5080 34960 5132 35012
rect 3792 34892 3844 34944
rect 26884 34960 26936 35012
rect 27252 35071 27304 35080
rect 27252 35037 27261 35071
rect 27261 35037 27295 35071
rect 27295 35037 27304 35071
rect 27436 35071 27488 35080
rect 27252 35028 27304 35037
rect 27436 35037 27445 35071
rect 27445 35037 27479 35071
rect 27479 35037 27488 35071
rect 27436 35028 27488 35037
rect 42432 35096 42484 35148
rect 42984 35096 43036 35148
rect 45560 35164 45612 35216
rect 38476 35071 38528 35080
rect 38476 35037 38485 35071
rect 38485 35037 38519 35071
rect 38519 35037 38528 35071
rect 38476 35028 38528 35037
rect 38752 35071 38804 35080
rect 38752 35037 38761 35071
rect 38761 35037 38795 35071
rect 38795 35037 38804 35071
rect 38752 35028 38804 35037
rect 55220 35164 55272 35216
rect 64788 35164 64840 35216
rect 52552 35096 52604 35148
rect 56968 35139 57020 35148
rect 56968 35105 56977 35139
rect 56977 35105 57011 35139
rect 57011 35105 57020 35139
rect 56968 35096 57020 35105
rect 63224 35096 63276 35148
rect 67916 35139 67968 35148
rect 67916 35105 67925 35139
rect 67925 35105 67959 35139
rect 67959 35105 67968 35139
rect 67916 35096 67968 35105
rect 68560 35096 68612 35148
rect 72884 35096 72936 35148
rect 75000 35139 75052 35148
rect 75000 35105 75009 35139
rect 75009 35105 75043 35139
rect 75043 35105 75052 35139
rect 75000 35096 75052 35105
rect 77024 35139 77076 35148
rect 75552 35071 75604 35080
rect 75552 35037 75561 35071
rect 75561 35037 75595 35071
rect 75595 35037 75604 35071
rect 75552 35028 75604 35037
rect 28080 35003 28132 35012
rect 28080 34969 28089 35003
rect 28089 34969 28123 35003
rect 28123 34969 28132 35003
rect 28080 34960 28132 34969
rect 37188 34960 37240 35012
rect 37648 34960 37700 35012
rect 39580 34960 39632 35012
rect 72148 35003 72200 35012
rect 72148 34969 72157 35003
rect 72157 34969 72191 35003
rect 72191 34969 72200 35003
rect 72148 34960 72200 34969
rect 75184 34960 75236 35012
rect 13912 34935 13964 34944
rect 13912 34901 13921 34935
rect 13921 34901 13955 34935
rect 13955 34901 13964 34935
rect 13912 34892 13964 34901
rect 14188 34935 14240 34944
rect 14188 34901 14197 34935
rect 14197 34901 14231 34935
rect 14231 34901 14240 34935
rect 14188 34892 14240 34901
rect 17224 34935 17276 34944
rect 17224 34901 17233 34935
rect 17233 34901 17267 34935
rect 17267 34901 17276 34935
rect 17224 34892 17276 34901
rect 20536 34892 20588 34944
rect 21916 34892 21968 34944
rect 32496 34892 32548 34944
rect 37372 34892 37424 34944
rect 37464 34892 37516 34944
rect 43260 34892 43312 34944
rect 43812 34892 43864 34944
rect 67732 34892 67784 34944
rect 68008 34935 68060 34944
rect 68008 34901 68017 34935
rect 68017 34901 68051 34935
rect 68051 34901 68060 34935
rect 68008 34892 68060 34901
rect 77024 35105 77033 35139
rect 77033 35105 77067 35139
rect 77067 35105 77076 35139
rect 77024 35096 77076 35105
rect 77208 35096 77260 35148
rect 87328 35096 87380 35148
rect 75828 34892 75880 34944
rect 76840 34892 76892 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 65686 34790 65738 34842
rect 65750 34790 65802 34842
rect 65814 34790 65866 34842
rect 65878 34790 65930 34842
rect 96406 34790 96458 34842
rect 96470 34790 96522 34842
rect 96534 34790 96586 34842
rect 96598 34790 96650 34842
rect 4896 34527 4948 34536
rect 4896 34493 4905 34527
rect 4905 34493 4939 34527
rect 4939 34493 4948 34527
rect 4896 34484 4948 34493
rect 19340 34688 19392 34740
rect 21824 34731 21876 34740
rect 7288 34663 7340 34672
rect 7288 34629 7297 34663
rect 7297 34629 7331 34663
rect 7331 34629 7340 34663
rect 7288 34620 7340 34629
rect 14188 34620 14240 34672
rect 15752 34620 15804 34672
rect 16672 34620 16724 34672
rect 7104 34527 7156 34536
rect 7104 34493 7113 34527
rect 7113 34493 7147 34527
rect 7147 34493 7156 34527
rect 7104 34484 7156 34493
rect 21824 34697 21833 34731
rect 21833 34697 21867 34731
rect 21867 34697 21876 34731
rect 21824 34688 21876 34697
rect 22008 34688 22060 34740
rect 21088 34620 21140 34672
rect 13820 34484 13872 34536
rect 15752 34527 15804 34536
rect 15752 34493 15761 34527
rect 15761 34493 15795 34527
rect 15795 34493 15804 34527
rect 15752 34484 15804 34493
rect 15844 34484 15896 34536
rect 16120 34484 16172 34536
rect 16212 34527 16264 34536
rect 16212 34493 16221 34527
rect 16221 34493 16255 34527
rect 16255 34493 16264 34527
rect 16212 34484 16264 34493
rect 16580 34484 16632 34536
rect 19892 34484 19944 34536
rect 20536 34484 20588 34536
rect 21088 34484 21140 34536
rect 25596 34552 25648 34604
rect 27436 34688 27488 34740
rect 27620 34688 27672 34740
rect 37280 34688 37332 34740
rect 38844 34688 38896 34740
rect 39672 34731 39724 34740
rect 39672 34697 39681 34731
rect 39681 34697 39715 34731
rect 39715 34697 39724 34731
rect 39672 34688 39724 34697
rect 49148 34688 49200 34740
rect 51448 34731 51500 34740
rect 51448 34697 51457 34731
rect 51457 34697 51491 34731
rect 51491 34697 51500 34731
rect 51448 34688 51500 34697
rect 27712 34620 27764 34672
rect 25688 34484 25740 34536
rect 25964 34552 26016 34604
rect 41604 34620 41656 34672
rect 44272 34663 44324 34672
rect 44272 34629 44281 34663
rect 44281 34629 44315 34663
rect 44315 34629 44324 34663
rect 44272 34620 44324 34629
rect 44364 34620 44416 34672
rect 52552 34620 52604 34672
rect 32404 34552 32456 34604
rect 32956 34552 33008 34604
rect 26148 34484 26200 34536
rect 5264 34416 5316 34468
rect 9036 34416 9088 34468
rect 6368 34348 6420 34400
rect 13176 34391 13228 34400
rect 13176 34357 13185 34391
rect 13185 34357 13219 34391
rect 13219 34357 13228 34391
rect 13176 34348 13228 34357
rect 15568 34416 15620 34468
rect 37280 34484 37332 34536
rect 37372 34527 37424 34536
rect 37372 34493 37381 34527
rect 37381 34493 37415 34527
rect 37415 34493 37424 34527
rect 38292 34552 38344 34604
rect 46940 34552 46992 34604
rect 56968 34688 57020 34740
rect 57060 34688 57112 34740
rect 59452 34595 59504 34604
rect 59452 34561 59461 34595
rect 59461 34561 59495 34595
rect 59495 34561 59504 34595
rect 59452 34552 59504 34561
rect 59728 34595 59780 34604
rect 59728 34561 59737 34595
rect 59737 34561 59771 34595
rect 59771 34561 59780 34595
rect 59728 34552 59780 34561
rect 59912 34552 59964 34604
rect 60924 34620 60976 34672
rect 63040 34688 63092 34740
rect 68100 34731 68152 34740
rect 68100 34697 68109 34731
rect 68109 34697 68143 34731
rect 68143 34697 68152 34731
rect 68100 34688 68152 34697
rect 68928 34688 68980 34740
rect 75736 34688 75788 34740
rect 77024 34688 77076 34740
rect 62580 34620 62632 34672
rect 68284 34663 68336 34672
rect 37372 34484 37424 34493
rect 38108 34484 38160 34536
rect 38200 34484 38252 34536
rect 39212 34484 39264 34536
rect 39672 34484 39724 34536
rect 39764 34484 39816 34536
rect 41512 34484 41564 34536
rect 42892 34527 42944 34536
rect 42892 34493 42901 34527
rect 42901 34493 42935 34527
rect 42935 34493 42944 34527
rect 42892 34484 42944 34493
rect 43260 34527 43312 34536
rect 43260 34493 43269 34527
rect 43269 34493 43303 34527
rect 43303 34493 43312 34527
rect 43260 34484 43312 34493
rect 43720 34527 43772 34536
rect 43720 34493 43729 34527
rect 43729 34493 43763 34527
rect 43763 34493 43772 34527
rect 43720 34484 43772 34493
rect 43812 34527 43864 34536
rect 43812 34493 43821 34527
rect 43821 34493 43855 34527
rect 43855 34493 43864 34527
rect 43812 34484 43864 34493
rect 43996 34484 44048 34536
rect 49700 34484 49752 34536
rect 52828 34484 52880 34536
rect 57704 34484 57756 34536
rect 62396 34484 62448 34536
rect 63040 34484 63092 34536
rect 68284 34629 68293 34663
rect 68293 34629 68327 34663
rect 68327 34629 68336 34663
rect 68284 34620 68336 34629
rect 68652 34620 68704 34672
rect 75000 34620 75052 34672
rect 68100 34552 68152 34604
rect 65984 34484 66036 34536
rect 16672 34348 16724 34400
rect 25780 34348 25832 34400
rect 27528 34391 27580 34400
rect 27528 34357 27537 34391
rect 27537 34357 27571 34391
rect 27571 34357 27580 34391
rect 27528 34348 27580 34357
rect 59544 34416 59596 34468
rect 36268 34348 36320 34400
rect 36452 34391 36504 34400
rect 36452 34357 36461 34391
rect 36461 34357 36495 34391
rect 36495 34357 36504 34391
rect 36452 34348 36504 34357
rect 37372 34348 37424 34400
rect 38200 34348 38252 34400
rect 39396 34391 39448 34400
rect 39396 34357 39405 34391
rect 39405 34357 39439 34391
rect 39439 34357 39448 34391
rect 39396 34348 39448 34357
rect 39488 34348 39540 34400
rect 54576 34348 54628 34400
rect 56048 34348 56100 34400
rect 65524 34416 65576 34468
rect 68836 34484 68888 34536
rect 68928 34484 68980 34536
rect 85396 34620 85448 34672
rect 77116 34552 77168 34604
rect 75828 34527 75880 34536
rect 75828 34493 75837 34527
rect 75837 34493 75871 34527
rect 75871 34493 75880 34527
rect 75828 34484 75880 34493
rect 77024 34527 77076 34536
rect 77024 34493 77033 34527
rect 77033 34493 77067 34527
rect 77067 34493 77076 34527
rect 77024 34484 77076 34493
rect 85028 34484 85080 34536
rect 85488 34484 85540 34536
rect 89812 34484 89864 34536
rect 62396 34391 62448 34400
rect 62396 34357 62405 34391
rect 62405 34357 62439 34391
rect 62439 34357 62448 34391
rect 62396 34348 62448 34357
rect 68744 34348 68796 34400
rect 76840 34459 76892 34468
rect 76840 34425 76849 34459
rect 76849 34425 76883 34459
rect 76883 34425 76892 34459
rect 76840 34416 76892 34425
rect 87144 34416 87196 34468
rect 88524 34459 88576 34468
rect 88524 34425 88533 34459
rect 88533 34425 88567 34459
rect 88567 34425 88576 34459
rect 88524 34416 88576 34425
rect 69756 34391 69808 34400
rect 69756 34357 69765 34391
rect 69765 34357 69799 34391
rect 69799 34357 69808 34391
rect 69756 34348 69808 34357
rect 70124 34391 70176 34400
rect 70124 34357 70133 34391
rect 70133 34357 70167 34391
rect 70167 34357 70176 34391
rect 70124 34348 70176 34357
rect 75828 34348 75880 34400
rect 76288 34348 76340 34400
rect 88340 34348 88392 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 81046 34246 81098 34298
rect 81110 34246 81162 34298
rect 81174 34246 81226 34298
rect 81238 34246 81290 34298
rect 2780 34144 2832 34196
rect 4896 34144 4948 34196
rect 6092 34144 6144 34196
rect 9312 34187 9364 34196
rect 9312 34153 9321 34187
rect 9321 34153 9355 34187
rect 9355 34153 9364 34187
rect 9312 34144 9364 34153
rect 11704 34144 11756 34196
rect 13820 34144 13872 34196
rect 18972 34144 19024 34196
rect 72424 34144 72476 34196
rect 75184 34187 75236 34196
rect 16672 34119 16724 34128
rect 4528 34051 4580 34060
rect 4528 34017 4537 34051
rect 4537 34017 4571 34051
rect 4571 34017 4580 34051
rect 4528 34008 4580 34017
rect 7104 34008 7156 34060
rect 9588 34008 9640 34060
rect 4896 33940 4948 33992
rect 11704 33983 11756 33992
rect 11704 33949 11713 33983
rect 11713 33949 11747 33983
rect 11747 33949 11756 33983
rect 11704 33940 11756 33949
rect 13176 34008 13228 34060
rect 15568 34051 15620 34060
rect 15568 34017 15577 34051
rect 15577 34017 15611 34051
rect 15611 34017 15620 34051
rect 15568 34008 15620 34017
rect 16672 34085 16681 34119
rect 16681 34085 16715 34119
rect 16715 34085 16724 34119
rect 16672 34076 16724 34085
rect 16488 34008 16540 34060
rect 27068 34076 27120 34128
rect 16856 34008 16908 34060
rect 18420 34051 18472 34060
rect 18052 33940 18104 33992
rect 18420 34017 18429 34051
rect 18429 34017 18463 34051
rect 18463 34017 18472 34051
rect 18420 34008 18472 34017
rect 21364 34008 21416 34060
rect 25412 34051 25464 34060
rect 25412 34017 25421 34051
rect 25421 34017 25455 34051
rect 25455 34017 25464 34051
rect 25412 34008 25464 34017
rect 26332 34008 26384 34060
rect 27160 34008 27212 34060
rect 27344 34008 27396 34060
rect 27620 34076 27672 34128
rect 37188 34119 37240 34128
rect 29276 34008 29328 34060
rect 32128 34051 32180 34060
rect 32128 34017 32137 34051
rect 32137 34017 32171 34051
rect 32171 34017 32180 34051
rect 32128 34008 32180 34017
rect 16396 33872 16448 33924
rect 21916 33915 21968 33924
rect 21916 33881 21925 33915
rect 21925 33881 21959 33915
rect 21959 33881 21968 33915
rect 21916 33872 21968 33881
rect 26056 33940 26108 33992
rect 26240 33983 26292 33992
rect 26240 33949 26249 33983
rect 26249 33949 26283 33983
rect 26283 33949 26292 33983
rect 26240 33940 26292 33949
rect 35532 33940 35584 33992
rect 27804 33872 27856 33924
rect 36452 33872 36504 33924
rect 37188 34085 37197 34119
rect 37197 34085 37231 34119
rect 37231 34085 37240 34119
rect 37188 34076 37240 34085
rect 38752 34076 38804 34128
rect 50988 34076 51040 34128
rect 56784 34119 56836 34128
rect 56784 34085 56793 34119
rect 56793 34085 56827 34119
rect 56827 34085 56836 34119
rect 56784 34076 56836 34085
rect 38844 34008 38896 34060
rect 39396 34008 39448 34060
rect 4988 33804 5040 33856
rect 13912 33804 13964 33856
rect 16488 33847 16540 33856
rect 16488 33813 16497 33847
rect 16497 33813 16531 33847
rect 16531 33813 16540 33847
rect 16488 33804 16540 33813
rect 17224 33804 17276 33856
rect 17960 33804 18012 33856
rect 19892 33804 19944 33856
rect 27712 33847 27764 33856
rect 27712 33813 27721 33847
rect 27721 33813 27755 33847
rect 27755 33813 27764 33847
rect 27712 33804 27764 33813
rect 31208 33804 31260 33856
rect 32036 33804 32088 33856
rect 32864 33804 32916 33856
rect 42892 33804 42944 33856
rect 44272 34008 44324 34060
rect 43812 33940 43864 33992
rect 45560 33940 45612 33992
rect 49240 33872 49292 33924
rect 50160 34008 50212 34060
rect 50712 34008 50764 34060
rect 55496 34051 55548 34060
rect 55496 34017 55505 34051
rect 55505 34017 55539 34051
rect 55539 34017 55548 34051
rect 56048 34051 56100 34060
rect 55496 34008 55548 34017
rect 56048 34017 56057 34051
rect 56057 34017 56091 34051
rect 56091 34017 56100 34051
rect 56048 34008 56100 34017
rect 54576 33983 54628 33992
rect 54576 33949 54585 33983
rect 54585 33949 54619 33983
rect 54619 33949 54628 33983
rect 54576 33940 54628 33949
rect 56692 33983 56744 33992
rect 56692 33949 56701 33983
rect 56701 33949 56735 33983
rect 56735 33949 56744 33983
rect 57520 34008 57572 34060
rect 57704 34051 57756 34060
rect 57704 34017 57713 34051
rect 57713 34017 57747 34051
rect 57747 34017 57756 34051
rect 57704 34008 57756 34017
rect 63132 34076 63184 34128
rect 65984 34076 66036 34128
rect 75184 34153 75193 34187
rect 75193 34153 75227 34187
rect 75227 34153 75236 34187
rect 75184 34144 75236 34153
rect 75736 34144 75788 34196
rect 82912 34144 82964 34196
rect 87972 34187 88024 34196
rect 87972 34153 87981 34187
rect 87981 34153 88015 34187
rect 88015 34153 88024 34187
rect 87972 34144 88024 34153
rect 77116 34076 77168 34128
rect 85028 34119 85080 34128
rect 56692 33940 56744 33949
rect 46848 33804 46900 33856
rect 60924 33940 60976 33992
rect 61292 33940 61344 33992
rect 58440 33872 58492 33924
rect 57704 33804 57756 33856
rect 58532 33847 58584 33856
rect 58532 33813 58541 33847
rect 58541 33813 58575 33847
rect 58575 33813 58584 33847
rect 58532 33804 58584 33813
rect 58624 33847 58676 33856
rect 58624 33813 58633 33847
rect 58633 33813 58667 33847
rect 58667 33813 58676 33847
rect 67640 33940 67692 33992
rect 73252 34051 73304 34060
rect 73252 34017 73261 34051
rect 73261 34017 73295 34051
rect 73295 34017 73304 34051
rect 73252 34008 73304 34017
rect 74448 34008 74500 34060
rect 75552 34008 75604 34060
rect 85028 34085 85037 34119
rect 85037 34085 85071 34119
rect 85071 34085 85080 34119
rect 85028 34076 85080 34085
rect 87144 34051 87196 34060
rect 87144 34017 87153 34051
rect 87153 34017 87187 34051
rect 87187 34017 87196 34051
rect 87144 34008 87196 34017
rect 87420 34008 87472 34060
rect 88432 34051 88484 34060
rect 88432 34017 88441 34051
rect 88441 34017 88475 34051
rect 88475 34017 88484 34051
rect 88432 34008 88484 34017
rect 88524 34051 88576 34060
rect 88524 34017 88533 34051
rect 88533 34017 88567 34051
rect 88567 34017 88576 34051
rect 89812 34051 89864 34060
rect 88524 34008 88576 34017
rect 89812 34017 89821 34051
rect 89821 34017 89855 34051
rect 89855 34017 89864 34051
rect 89812 34008 89864 34017
rect 68560 33983 68612 33992
rect 68560 33949 68569 33983
rect 68569 33949 68603 33983
rect 68603 33949 68612 33983
rect 68560 33940 68612 33949
rect 74264 33983 74316 33992
rect 74264 33949 74273 33983
rect 74273 33949 74307 33983
rect 74307 33949 74316 33983
rect 75736 33983 75788 33992
rect 74264 33940 74316 33949
rect 75736 33949 75745 33983
rect 75745 33949 75779 33983
rect 75779 33949 75788 33983
rect 75736 33940 75788 33949
rect 78680 33940 78732 33992
rect 73988 33872 74040 33924
rect 76840 33872 76892 33924
rect 77208 33872 77260 33924
rect 85488 33940 85540 33992
rect 88340 33872 88392 33924
rect 75552 33847 75604 33856
rect 58624 33804 58676 33813
rect 75552 33813 75576 33847
rect 75576 33813 75604 33847
rect 75552 33804 75604 33813
rect 75828 33804 75880 33856
rect 77484 33847 77536 33856
rect 77484 33813 77493 33847
rect 77493 33813 77527 33847
rect 77527 33813 77536 33847
rect 77484 33804 77536 33813
rect 83188 33847 83240 33856
rect 83188 33813 83197 33847
rect 83197 33813 83231 33847
rect 83231 33813 83240 33847
rect 83188 33804 83240 33813
rect 87236 33847 87288 33856
rect 87236 33813 87245 33847
rect 87245 33813 87279 33847
rect 87279 33813 87288 33847
rect 87236 33804 87288 33813
rect 88524 33804 88576 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 65686 33702 65738 33754
rect 65750 33702 65802 33754
rect 65814 33702 65866 33754
rect 65878 33702 65930 33754
rect 96406 33702 96458 33754
rect 96470 33702 96522 33754
rect 96534 33702 96586 33754
rect 96598 33702 96650 33754
rect 4712 33600 4764 33652
rect 22744 33600 22796 33652
rect 46940 33600 46992 33652
rect 49240 33643 49292 33652
rect 49240 33609 49249 33643
rect 49249 33609 49283 33643
rect 49283 33609 49292 33643
rect 49240 33600 49292 33609
rect 50804 33600 50856 33652
rect 50988 33600 51040 33652
rect 9312 33532 9364 33584
rect 12900 33532 12952 33584
rect 14924 33532 14976 33584
rect 17316 33575 17368 33584
rect 17316 33541 17325 33575
rect 17325 33541 17359 33575
rect 17359 33541 17368 33575
rect 17316 33532 17368 33541
rect 18972 33575 19024 33584
rect 18972 33541 18981 33575
rect 18981 33541 19015 33575
rect 19015 33541 19024 33575
rect 18972 33532 19024 33541
rect 24676 33532 24728 33584
rect 26056 33532 26108 33584
rect 32128 33575 32180 33584
rect 32128 33541 32137 33575
rect 32137 33541 32171 33575
rect 32171 33541 32180 33575
rect 32128 33532 32180 33541
rect 33140 33575 33192 33584
rect 33140 33541 33149 33575
rect 33149 33541 33183 33575
rect 33183 33541 33192 33575
rect 33140 33532 33192 33541
rect 36268 33532 36320 33584
rect 38752 33532 38804 33584
rect 3608 33464 3660 33516
rect 3976 33464 4028 33516
rect 19248 33464 19300 33516
rect 19340 33464 19392 33516
rect 32864 33464 32916 33516
rect 35532 33464 35584 33516
rect 38660 33464 38712 33516
rect 49240 33464 49292 33516
rect 54576 33600 54628 33652
rect 56876 33643 56928 33652
rect 56876 33609 56885 33643
rect 56885 33609 56919 33643
rect 56919 33609 56928 33643
rect 56876 33600 56928 33609
rect 57520 33600 57572 33652
rect 58624 33600 58676 33652
rect 7104 33396 7156 33448
rect 9312 33439 9364 33448
rect 9312 33405 9321 33439
rect 9321 33405 9355 33439
rect 9355 33405 9364 33439
rect 9312 33396 9364 33405
rect 14924 33396 14976 33448
rect 16212 33396 16264 33448
rect 16672 33396 16724 33448
rect 17316 33396 17368 33448
rect 18052 33439 18104 33448
rect 18052 33405 18061 33439
rect 18061 33405 18095 33439
rect 18095 33405 18104 33439
rect 18052 33396 18104 33405
rect 18328 33439 18380 33448
rect 18328 33405 18337 33439
rect 18337 33405 18371 33439
rect 18371 33405 18380 33439
rect 18328 33396 18380 33405
rect 19892 33439 19944 33448
rect 19892 33405 19901 33439
rect 19901 33405 19935 33439
rect 19935 33405 19944 33439
rect 19892 33396 19944 33405
rect 21364 33396 21416 33448
rect 24860 33396 24912 33448
rect 8944 33328 8996 33380
rect 4160 33303 4212 33312
rect 4160 33269 4169 33303
rect 4169 33269 4203 33303
rect 4203 33269 4212 33303
rect 4160 33260 4212 33269
rect 8024 33260 8076 33312
rect 9220 33260 9272 33312
rect 10784 33260 10836 33312
rect 16396 33260 16448 33312
rect 16488 33260 16540 33312
rect 17960 33260 18012 33312
rect 18328 33260 18380 33312
rect 18512 33303 18564 33312
rect 18512 33269 18521 33303
rect 18521 33269 18555 33303
rect 18555 33269 18564 33303
rect 18512 33260 18564 33269
rect 19984 33303 20036 33312
rect 19984 33269 19993 33303
rect 19993 33269 20027 33303
rect 20027 33269 20036 33303
rect 19984 33260 20036 33269
rect 24124 33328 24176 33380
rect 24676 33328 24728 33380
rect 26056 33396 26108 33448
rect 27620 33396 27672 33448
rect 30564 33439 30616 33448
rect 30564 33405 30573 33439
rect 30573 33405 30607 33439
rect 30607 33405 30616 33439
rect 30564 33396 30616 33405
rect 30840 33439 30892 33448
rect 30840 33405 30849 33439
rect 30849 33405 30883 33439
rect 30883 33405 30892 33439
rect 30840 33396 30892 33405
rect 33232 33396 33284 33448
rect 35440 33439 35492 33448
rect 35440 33405 35449 33439
rect 35449 33405 35483 33439
rect 35483 33405 35492 33439
rect 35440 33396 35492 33405
rect 37372 33396 37424 33448
rect 38292 33439 38344 33448
rect 38292 33405 38301 33439
rect 38301 33405 38335 33439
rect 38335 33405 38344 33439
rect 38292 33396 38344 33405
rect 27252 33260 27304 33312
rect 27528 33303 27580 33312
rect 27528 33269 27537 33303
rect 27537 33269 27571 33303
rect 27571 33269 27580 33303
rect 27528 33260 27580 33269
rect 27712 33328 27764 33380
rect 30656 33328 30708 33380
rect 38568 33328 38620 33380
rect 41880 33396 41932 33448
rect 46848 33396 46900 33448
rect 38844 33328 38896 33380
rect 32128 33260 32180 33312
rect 32312 33303 32364 33312
rect 32312 33269 32321 33303
rect 32321 33269 32355 33303
rect 32355 33269 32364 33303
rect 32312 33260 32364 33269
rect 33232 33260 33284 33312
rect 38292 33260 38344 33312
rect 42340 33260 42392 33312
rect 51172 33396 51224 33448
rect 55496 33532 55548 33584
rect 51448 33371 51500 33380
rect 51448 33337 51457 33371
rect 51457 33337 51491 33371
rect 51491 33337 51500 33371
rect 51448 33328 51500 33337
rect 51816 33371 51868 33380
rect 51816 33337 51825 33371
rect 51825 33337 51859 33371
rect 51859 33337 51868 33371
rect 51816 33328 51868 33337
rect 52828 33439 52880 33448
rect 52828 33405 52837 33439
rect 52837 33405 52871 33439
rect 52871 33405 52880 33439
rect 52828 33396 52880 33405
rect 53012 33439 53064 33448
rect 53012 33405 53021 33439
rect 53021 33405 53055 33439
rect 53055 33405 53064 33439
rect 53012 33396 53064 33405
rect 54576 33396 54628 33448
rect 58440 33532 58492 33584
rect 57520 33439 57572 33448
rect 57520 33405 57529 33439
rect 57529 33405 57563 33439
rect 57563 33405 57572 33439
rect 57520 33396 57572 33405
rect 57060 33371 57112 33380
rect 53012 33260 53064 33312
rect 57060 33337 57069 33371
rect 57069 33337 57103 33371
rect 57103 33337 57112 33371
rect 57060 33328 57112 33337
rect 58072 33328 58124 33380
rect 58256 33396 58308 33448
rect 68008 33600 68060 33652
rect 69480 33600 69532 33652
rect 85488 33643 85540 33652
rect 85488 33609 85497 33643
rect 85497 33609 85531 33643
rect 85531 33609 85540 33643
rect 85488 33600 85540 33609
rect 87144 33600 87196 33652
rect 89812 33643 89864 33652
rect 89812 33609 89821 33643
rect 89821 33609 89855 33643
rect 89855 33609 89864 33643
rect 89812 33600 89864 33609
rect 61660 33532 61712 33584
rect 69664 33532 69716 33584
rect 62580 33464 62632 33516
rect 69756 33464 69808 33516
rect 77484 33464 77536 33516
rect 61108 33396 61160 33448
rect 61384 33439 61436 33448
rect 61384 33405 61393 33439
rect 61393 33405 61427 33439
rect 61427 33405 61436 33439
rect 61384 33396 61436 33405
rect 69296 33439 69348 33448
rect 69296 33405 69305 33439
rect 69305 33405 69339 33439
rect 69339 33405 69348 33439
rect 69296 33396 69348 33405
rect 75920 33396 75972 33448
rect 77300 33396 77352 33448
rect 77760 33439 77812 33448
rect 77760 33405 77769 33439
rect 77769 33405 77803 33439
rect 77803 33405 77812 33439
rect 83188 33464 83240 33516
rect 88524 33507 88576 33516
rect 77760 33396 77812 33405
rect 81532 33396 81584 33448
rect 85672 33396 85724 33448
rect 63132 33328 63184 33380
rect 58532 33260 58584 33312
rect 75552 33328 75604 33380
rect 88524 33473 88533 33507
rect 88533 33473 88567 33507
rect 88567 33473 88576 33507
rect 88524 33464 88576 33473
rect 86776 33371 86828 33380
rect 86776 33337 86785 33371
rect 86785 33337 86819 33371
rect 86819 33337 86828 33371
rect 86776 33328 86828 33337
rect 77392 33303 77444 33312
rect 77392 33269 77401 33303
rect 77401 33269 77435 33303
rect 77435 33269 77444 33303
rect 77392 33260 77444 33269
rect 82268 33303 82320 33312
rect 82268 33269 82277 33303
rect 82277 33269 82311 33303
rect 82311 33269 82320 33303
rect 82268 33260 82320 33269
rect 86684 33303 86736 33312
rect 86684 33269 86693 33303
rect 86693 33269 86727 33303
rect 86727 33269 86736 33303
rect 86684 33260 86736 33269
rect 87972 33260 88024 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 50326 33158 50378 33210
rect 50390 33158 50442 33210
rect 50454 33158 50506 33210
rect 50518 33158 50570 33210
rect 81046 33158 81098 33210
rect 81110 33158 81162 33210
rect 81174 33158 81226 33210
rect 81238 33158 81290 33210
rect 3792 33056 3844 33108
rect 7564 33056 7616 33108
rect 8944 33099 8996 33108
rect 8944 33065 8953 33099
rect 8953 33065 8987 33099
rect 8987 33065 8996 33099
rect 8944 33056 8996 33065
rect 8024 32963 8076 32972
rect 8024 32929 8033 32963
rect 8033 32929 8067 32963
rect 8067 32929 8076 32963
rect 8024 32920 8076 32929
rect 8944 32920 8996 32972
rect 62028 33056 62080 33108
rect 11704 32988 11756 33040
rect 18420 32988 18472 33040
rect 24860 32988 24912 33040
rect 25320 32988 25372 33040
rect 27712 32988 27764 33040
rect 29276 33031 29328 33040
rect 29276 32997 29285 33031
rect 29285 32997 29319 33031
rect 29319 32997 29328 33031
rect 29276 32988 29328 32997
rect 8668 32895 8720 32904
rect 8668 32861 8677 32895
rect 8677 32861 8711 32895
rect 8711 32861 8720 32895
rect 8668 32852 8720 32861
rect 10416 32895 10468 32904
rect 10416 32861 10425 32895
rect 10425 32861 10459 32895
rect 10459 32861 10468 32895
rect 10416 32852 10468 32861
rect 16856 32852 16908 32904
rect 16672 32759 16724 32768
rect 16672 32725 16681 32759
rect 16681 32725 16715 32759
rect 16715 32725 16724 32759
rect 19616 32963 19668 32972
rect 19616 32929 19625 32963
rect 19625 32929 19659 32963
rect 19659 32929 19668 32963
rect 19616 32920 19668 32929
rect 21548 32920 21600 32972
rect 30840 32988 30892 33040
rect 25228 32852 25280 32904
rect 26148 32852 26200 32904
rect 20628 32784 20680 32836
rect 23756 32784 23808 32836
rect 16672 32716 16724 32725
rect 24308 32716 24360 32768
rect 30564 32920 30616 32972
rect 31576 32988 31628 33040
rect 32128 32988 32180 33040
rect 31392 32920 31444 32972
rect 33140 32988 33192 33040
rect 49148 33031 49200 33040
rect 49148 32997 49157 33031
rect 49157 32997 49191 33031
rect 49191 32997 49200 33031
rect 49148 32988 49200 32997
rect 31208 32827 31260 32836
rect 31208 32793 31217 32827
rect 31217 32793 31251 32827
rect 31251 32793 31260 32827
rect 31208 32784 31260 32793
rect 37924 32920 37976 32972
rect 41972 32920 42024 32972
rect 49700 32920 49752 32972
rect 51448 32988 51500 33040
rect 43444 32852 43496 32904
rect 43812 32895 43864 32904
rect 43812 32861 43821 32895
rect 43821 32861 43855 32895
rect 43855 32861 43864 32895
rect 43812 32852 43864 32861
rect 44088 32895 44140 32904
rect 44088 32861 44097 32895
rect 44097 32861 44131 32895
rect 44131 32861 44140 32895
rect 44088 32852 44140 32861
rect 50160 32852 50212 32904
rect 51172 32920 51224 32972
rect 55864 32920 55916 32972
rect 61568 32920 61620 32972
rect 61844 32963 61896 32972
rect 61844 32929 61853 32963
rect 61853 32929 61887 32963
rect 61887 32929 61896 32963
rect 61844 32920 61896 32929
rect 62028 32963 62080 32972
rect 62028 32929 62037 32963
rect 62037 32929 62071 32963
rect 62071 32929 62080 32963
rect 62028 32920 62080 32929
rect 50988 32852 51040 32904
rect 53380 32852 53432 32904
rect 56692 32852 56744 32904
rect 62396 32920 62448 32972
rect 63040 32920 63092 32972
rect 67916 33056 67968 33108
rect 68744 33099 68796 33108
rect 68744 33065 68753 33099
rect 68753 33065 68787 33099
rect 68787 33065 68796 33099
rect 68744 33056 68796 33065
rect 75552 33099 75604 33108
rect 75552 33065 75561 33099
rect 75561 33065 75595 33099
rect 75595 33065 75604 33099
rect 75552 33056 75604 33065
rect 77760 33099 77812 33108
rect 77760 33065 77769 33099
rect 77769 33065 77803 33099
rect 77803 33065 77812 33099
rect 77760 33056 77812 33065
rect 85212 33056 85264 33108
rect 66996 33031 67048 33040
rect 66996 32997 67005 33031
rect 67005 32997 67039 33031
rect 67039 32997 67048 33031
rect 66996 32988 67048 32997
rect 69296 32988 69348 33040
rect 76012 32988 76064 33040
rect 67456 32963 67508 32972
rect 67456 32929 67465 32963
rect 67465 32929 67499 32963
rect 67499 32929 67508 32963
rect 67916 32963 67968 32972
rect 67456 32920 67508 32929
rect 67916 32929 67925 32963
rect 67925 32929 67959 32963
rect 67959 32929 67968 32963
rect 67916 32920 67968 32929
rect 68100 32963 68152 32972
rect 68100 32929 68109 32963
rect 68109 32929 68143 32963
rect 68143 32929 68152 32963
rect 68100 32920 68152 32929
rect 73988 32963 74040 32972
rect 73988 32929 73997 32963
rect 73997 32929 74031 32963
rect 74031 32929 74040 32963
rect 73988 32920 74040 32929
rect 74264 32963 74316 32972
rect 74264 32929 74273 32963
rect 74273 32929 74307 32963
rect 74307 32929 74316 32963
rect 74264 32920 74316 32929
rect 74448 32963 74500 32972
rect 74448 32929 74457 32963
rect 74457 32929 74491 32963
rect 74491 32929 74500 32963
rect 74448 32920 74500 32929
rect 37188 32784 37240 32836
rect 42340 32827 42392 32836
rect 42340 32793 42349 32827
rect 42349 32793 42383 32827
rect 42383 32793 42392 32827
rect 42340 32784 42392 32793
rect 68836 32852 68888 32904
rect 31852 32716 31904 32768
rect 37924 32759 37976 32768
rect 37924 32725 37933 32759
rect 37933 32725 37967 32759
rect 37967 32725 37976 32759
rect 37924 32716 37976 32725
rect 41788 32716 41840 32768
rect 41972 32759 42024 32768
rect 41972 32725 41981 32759
rect 41981 32725 42015 32759
rect 42015 32725 42024 32759
rect 41972 32716 42024 32725
rect 42432 32716 42484 32768
rect 74264 32784 74316 32836
rect 63224 32716 63276 32768
rect 63500 32759 63552 32768
rect 63500 32725 63509 32759
rect 63509 32725 63543 32759
rect 63543 32725 63552 32759
rect 63500 32716 63552 32725
rect 66996 32716 67048 32768
rect 68100 32716 68152 32768
rect 69940 32716 69992 32768
rect 77392 32920 77444 32972
rect 82268 32988 82320 33040
rect 82544 32988 82596 33040
rect 80520 32963 80572 32972
rect 80520 32929 80529 32963
rect 80529 32929 80563 32963
rect 80563 32929 80572 32963
rect 80520 32920 80572 32929
rect 82360 32920 82412 32972
rect 82452 32852 82504 32904
rect 85028 32852 85080 32904
rect 88432 33056 88484 33108
rect 85672 33031 85724 33040
rect 85672 32997 85681 33031
rect 85681 32997 85715 33031
rect 85715 32997 85724 33031
rect 85672 32988 85724 32997
rect 87236 32988 87288 33040
rect 86684 32963 86736 32972
rect 86684 32929 86693 32963
rect 86693 32929 86727 32963
rect 86727 32929 86736 32963
rect 86684 32920 86736 32929
rect 86776 32963 86828 32972
rect 86776 32929 86785 32963
rect 86785 32929 86819 32963
rect 86819 32929 86828 32963
rect 86776 32920 86828 32929
rect 88340 32920 88392 32972
rect 75184 32784 75236 32836
rect 82084 32784 82136 32836
rect 82544 32716 82596 32768
rect 85580 32759 85632 32768
rect 85580 32725 85589 32759
rect 85589 32725 85623 32759
rect 85623 32725 85632 32759
rect 85580 32716 85632 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 65686 32614 65738 32666
rect 65750 32614 65802 32666
rect 65814 32614 65866 32666
rect 65878 32614 65930 32666
rect 96406 32614 96458 32666
rect 96470 32614 96522 32666
rect 96534 32614 96586 32666
rect 96598 32614 96650 32666
rect 3792 32512 3844 32564
rect 6552 32444 6604 32496
rect 9956 32512 10008 32564
rect 10784 32512 10836 32564
rect 15844 32487 15896 32496
rect 3148 32419 3200 32428
rect 3148 32385 3157 32419
rect 3157 32385 3191 32419
rect 3191 32385 3200 32419
rect 3148 32376 3200 32385
rect 8484 32419 8536 32428
rect 8484 32385 8493 32419
rect 8493 32385 8527 32419
rect 8527 32385 8536 32419
rect 8484 32376 8536 32385
rect 2964 32308 3016 32360
rect 8024 32351 8076 32360
rect 8024 32317 8033 32351
rect 8033 32317 8067 32351
rect 8067 32317 8076 32351
rect 8024 32308 8076 32317
rect 9404 32376 9456 32428
rect 15844 32453 15853 32487
rect 15853 32453 15887 32487
rect 15887 32453 15896 32487
rect 15844 32444 15896 32453
rect 16856 32487 16908 32496
rect 16856 32453 16865 32487
rect 16865 32453 16899 32487
rect 16899 32453 16908 32487
rect 16856 32444 16908 32453
rect 19616 32444 19668 32496
rect 21364 32487 21416 32496
rect 10048 32419 10100 32428
rect 10048 32385 10057 32419
rect 10057 32385 10091 32419
rect 10091 32385 10100 32419
rect 10048 32376 10100 32385
rect 9956 32351 10008 32360
rect 9956 32317 9965 32351
rect 9965 32317 9999 32351
rect 9999 32317 10008 32351
rect 9956 32308 10008 32317
rect 15660 32351 15712 32360
rect 15660 32317 15669 32351
rect 15669 32317 15703 32351
rect 15703 32317 15712 32351
rect 15660 32308 15712 32317
rect 18512 32308 18564 32360
rect 19984 32351 20036 32360
rect 16672 32240 16724 32292
rect 17960 32240 18012 32292
rect 19984 32317 19993 32351
rect 19993 32317 20027 32351
rect 20027 32317 20036 32351
rect 19984 32308 20036 32317
rect 21364 32453 21373 32487
rect 21373 32453 21407 32487
rect 21407 32453 21416 32487
rect 21364 32444 21416 32453
rect 21548 32487 21600 32496
rect 21548 32453 21557 32487
rect 21557 32453 21591 32487
rect 21591 32453 21600 32487
rect 21548 32444 21600 32453
rect 25596 32444 25648 32496
rect 25228 32376 25280 32428
rect 26056 32419 26108 32428
rect 26056 32385 26065 32419
rect 26065 32385 26099 32419
rect 26099 32385 26108 32419
rect 26056 32376 26108 32385
rect 27160 32444 27212 32496
rect 29368 32444 29420 32496
rect 31392 32444 31444 32496
rect 36176 32555 36228 32564
rect 36176 32521 36185 32555
rect 36185 32521 36219 32555
rect 36219 32521 36228 32555
rect 36176 32512 36228 32521
rect 37188 32512 37240 32564
rect 44088 32512 44140 32564
rect 53564 32512 53616 32564
rect 53656 32512 53708 32564
rect 62304 32512 62356 32564
rect 69940 32512 69992 32564
rect 41604 32444 41656 32496
rect 42432 32487 42484 32496
rect 42432 32453 42441 32487
rect 42441 32453 42475 32487
rect 42475 32453 42484 32487
rect 42432 32444 42484 32453
rect 42984 32487 43036 32496
rect 42984 32453 42993 32487
rect 42993 32453 43027 32487
rect 43027 32453 43036 32487
rect 42984 32444 43036 32453
rect 31576 32419 31628 32428
rect 31576 32385 31585 32419
rect 31585 32385 31619 32419
rect 31619 32385 31628 32419
rect 31576 32376 31628 32385
rect 31852 32419 31904 32428
rect 31852 32385 31861 32419
rect 31861 32385 31895 32419
rect 31895 32385 31904 32419
rect 31852 32376 31904 32385
rect 34336 32376 34388 32428
rect 40960 32419 41012 32428
rect 25596 32351 25648 32360
rect 25596 32317 25605 32351
rect 25605 32317 25639 32351
rect 25639 32317 25648 32351
rect 25596 32308 25648 32317
rect 26332 32308 26384 32360
rect 27068 32351 27120 32360
rect 21732 32283 21784 32292
rect 21732 32249 21741 32283
rect 21741 32249 21775 32283
rect 21775 32249 21784 32283
rect 21732 32240 21784 32249
rect 2872 32172 2924 32224
rect 4712 32215 4764 32224
rect 4712 32181 4721 32215
rect 4721 32181 4755 32215
rect 4755 32181 4764 32215
rect 4712 32172 4764 32181
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 22284 32172 22336 32224
rect 27068 32317 27077 32351
rect 27077 32317 27111 32351
rect 27111 32317 27120 32351
rect 27068 32308 27120 32317
rect 27160 32308 27212 32360
rect 33232 32351 33284 32360
rect 33232 32317 33241 32351
rect 33241 32317 33275 32351
rect 33275 32317 33284 32351
rect 33232 32308 33284 32317
rect 36176 32308 36228 32360
rect 40960 32385 40969 32419
rect 40969 32385 41003 32419
rect 41003 32385 41012 32419
rect 40960 32376 41012 32385
rect 61660 32487 61712 32496
rect 61660 32453 61669 32487
rect 61669 32453 61703 32487
rect 61703 32453 61712 32487
rect 61660 32444 61712 32453
rect 69664 32487 69716 32496
rect 69664 32453 69673 32487
rect 69673 32453 69707 32487
rect 69707 32453 69716 32487
rect 69664 32444 69716 32453
rect 54300 32419 54352 32428
rect 54300 32385 54309 32419
rect 54309 32385 54343 32419
rect 54343 32385 54352 32419
rect 54300 32376 54352 32385
rect 54852 32376 54904 32428
rect 57060 32376 57112 32428
rect 67088 32376 67140 32428
rect 67456 32376 67508 32428
rect 37924 32308 37976 32360
rect 41604 32351 41656 32360
rect 41604 32317 41613 32351
rect 41613 32317 41647 32351
rect 41647 32317 41656 32351
rect 41604 32308 41656 32317
rect 42340 32308 42392 32360
rect 42984 32308 43036 32360
rect 44364 32351 44416 32360
rect 44364 32317 44373 32351
rect 44373 32317 44407 32351
rect 44407 32317 44416 32351
rect 44364 32308 44416 32317
rect 48044 32308 48096 32360
rect 53472 32308 53524 32360
rect 53748 32351 53800 32360
rect 53748 32317 53757 32351
rect 53757 32317 53791 32351
rect 53791 32317 53800 32351
rect 53748 32308 53800 32317
rect 55036 32308 55088 32360
rect 41236 32240 41288 32292
rect 31576 32172 31628 32224
rect 35072 32215 35124 32224
rect 35072 32181 35081 32215
rect 35081 32181 35115 32215
rect 35115 32181 35124 32215
rect 35072 32172 35124 32181
rect 36544 32215 36596 32224
rect 36544 32181 36553 32215
rect 36553 32181 36587 32215
rect 36587 32181 36596 32215
rect 36544 32172 36596 32181
rect 36636 32172 36688 32224
rect 41972 32172 42024 32224
rect 42708 32240 42760 32292
rect 55864 32240 55916 32292
rect 42800 32172 42852 32224
rect 44548 32172 44600 32224
rect 48504 32172 48556 32224
rect 55036 32215 55088 32224
rect 55036 32181 55045 32215
rect 55045 32181 55079 32215
rect 55079 32181 55088 32215
rect 55036 32172 55088 32181
rect 60280 32172 60332 32224
rect 61844 32308 61896 32360
rect 63500 32308 63552 32360
rect 62028 32240 62080 32292
rect 62120 32172 62172 32224
rect 62396 32215 62448 32224
rect 62396 32181 62405 32215
rect 62405 32181 62439 32215
rect 62439 32181 62448 32215
rect 62396 32172 62448 32181
rect 67548 32172 67600 32224
rect 69296 32351 69348 32360
rect 69296 32317 69305 32351
rect 69305 32317 69339 32351
rect 69339 32317 69348 32351
rect 86960 32512 87012 32564
rect 76012 32444 76064 32496
rect 85580 32444 85632 32496
rect 69296 32308 69348 32317
rect 80520 32376 80572 32428
rect 81532 32419 81584 32428
rect 81532 32385 81541 32419
rect 81541 32385 81575 32419
rect 81575 32385 81584 32419
rect 81532 32376 81584 32385
rect 82084 32419 82136 32428
rect 82084 32385 82093 32419
rect 82093 32385 82127 32419
rect 82127 32385 82136 32419
rect 82084 32376 82136 32385
rect 82544 32419 82596 32428
rect 82544 32385 82553 32419
rect 82553 32385 82587 32419
rect 82587 32385 82596 32419
rect 82544 32376 82596 32385
rect 74264 32308 74316 32360
rect 82452 32308 82504 32360
rect 75920 32283 75972 32292
rect 75920 32249 75929 32283
rect 75929 32249 75963 32283
rect 75963 32249 75972 32283
rect 75920 32240 75972 32249
rect 82728 32240 82780 32292
rect 75552 32215 75604 32224
rect 75552 32181 75561 32215
rect 75561 32181 75595 32215
rect 75595 32181 75604 32215
rect 75552 32172 75604 32181
rect 80888 32172 80940 32224
rect 85396 32172 85448 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 50326 32070 50378 32122
rect 50390 32070 50442 32122
rect 50454 32070 50506 32122
rect 50518 32070 50570 32122
rect 81046 32070 81098 32122
rect 81110 32070 81162 32122
rect 81174 32070 81226 32122
rect 81238 32070 81290 32122
rect 11704 31968 11756 32020
rect 32956 31968 33008 32020
rect 36636 31968 36688 32020
rect 40960 32011 41012 32020
rect 40960 31977 40969 32011
rect 40969 31977 41003 32011
rect 41003 31977 41012 32011
rect 40960 31968 41012 31977
rect 42708 31968 42760 32020
rect 42800 32011 42852 32020
rect 42800 31977 42809 32011
rect 42809 31977 42843 32011
rect 42843 31977 42852 32011
rect 42800 31968 42852 31977
rect 44364 31968 44416 32020
rect 52368 31968 52420 32020
rect 53748 31968 53800 32020
rect 54852 32011 54904 32020
rect 54852 31977 54861 32011
rect 54861 31977 54895 32011
rect 54895 31977 54904 32011
rect 54852 31968 54904 31977
rect 55036 31968 55088 32020
rect 62304 31968 62356 32020
rect 62396 31968 62448 32020
rect 16120 31900 16172 31952
rect 17040 31875 17092 31884
rect 17040 31841 17049 31875
rect 17049 31841 17083 31875
rect 17083 31841 17092 31875
rect 17040 31832 17092 31841
rect 17408 31875 17460 31884
rect 11244 31807 11296 31816
rect 11244 31773 11253 31807
rect 11253 31773 11287 31807
rect 11287 31773 11296 31807
rect 11244 31764 11296 31773
rect 15384 31764 15436 31816
rect 16580 31807 16632 31816
rect 12440 31696 12492 31748
rect 16580 31773 16589 31807
rect 16589 31773 16623 31807
rect 16623 31773 16632 31807
rect 16580 31764 16632 31773
rect 17408 31841 17417 31875
rect 17417 31841 17451 31875
rect 17451 31841 17460 31875
rect 17408 31832 17460 31841
rect 41512 31900 41564 31952
rect 17960 31807 18012 31816
rect 17960 31773 17969 31807
rect 17969 31773 18003 31807
rect 18003 31773 18012 31807
rect 17960 31764 18012 31773
rect 19984 31832 20036 31884
rect 25412 31764 25464 31816
rect 27068 31764 27120 31816
rect 35072 31832 35124 31884
rect 41236 31875 41288 31884
rect 41236 31841 41245 31875
rect 41245 31841 41279 31875
rect 41279 31841 41288 31875
rect 41880 31875 41932 31884
rect 41236 31832 41288 31841
rect 41880 31841 41885 31875
rect 41885 31841 41919 31875
rect 41919 31841 41932 31875
rect 41880 31832 41932 31841
rect 44548 31900 44600 31952
rect 56232 31900 56284 31952
rect 40960 31764 41012 31816
rect 18236 31739 18288 31748
rect 12992 31628 13044 31680
rect 18236 31705 18245 31739
rect 18245 31705 18279 31739
rect 18279 31705 18288 31739
rect 18236 31696 18288 31705
rect 17408 31628 17460 31680
rect 19432 31628 19484 31680
rect 21364 31696 21416 31748
rect 34796 31696 34848 31748
rect 41880 31696 41932 31748
rect 53196 31832 53248 31884
rect 53380 31832 53432 31884
rect 42708 31764 42760 31816
rect 43352 31807 43404 31816
rect 43352 31773 43361 31807
rect 43361 31773 43395 31807
rect 43395 31773 43404 31807
rect 43352 31764 43404 31773
rect 48320 31764 48372 31816
rect 53656 31764 53708 31816
rect 54944 31696 54996 31748
rect 67548 31900 67600 31952
rect 67180 31832 67232 31884
rect 74448 32011 74500 32020
rect 74448 31977 74457 32011
rect 74457 31977 74491 32011
rect 74491 31977 74500 32011
rect 74448 31968 74500 31977
rect 76012 32011 76064 32020
rect 76012 31977 76021 32011
rect 76021 31977 76055 32011
rect 76055 31977 76064 32011
rect 76012 31968 76064 31977
rect 75184 31900 75236 31952
rect 69020 31832 69072 31884
rect 75552 31832 75604 31884
rect 75736 31832 75788 31884
rect 80888 31968 80940 32020
rect 81440 31968 81492 32020
rect 78680 31832 78732 31884
rect 79784 31832 79836 31884
rect 82268 31900 82320 31952
rect 85396 31875 85448 31884
rect 85396 31841 85405 31875
rect 85405 31841 85439 31875
rect 85439 31841 85448 31875
rect 85396 31832 85448 31841
rect 66904 31807 66956 31816
rect 66904 31773 66913 31807
rect 66913 31773 66947 31807
rect 66947 31773 66956 31807
rect 66904 31764 66956 31773
rect 67272 31807 67324 31816
rect 67272 31773 67281 31807
rect 67281 31773 67315 31807
rect 67315 31773 67324 31807
rect 67272 31764 67324 31773
rect 80888 31807 80940 31816
rect 80888 31773 80897 31807
rect 80897 31773 80931 31807
rect 80931 31773 80940 31807
rect 80888 31764 80940 31773
rect 82820 31764 82872 31816
rect 86960 31875 87012 31884
rect 86960 31841 86969 31875
rect 86969 31841 87003 31875
rect 87003 31841 87012 31875
rect 86960 31832 87012 31841
rect 87696 31832 87748 31884
rect 88248 31875 88300 31884
rect 88248 31841 88257 31875
rect 88257 31841 88291 31875
rect 88291 31841 88300 31875
rect 88248 31832 88300 31841
rect 50160 31628 50212 31680
rect 53196 31628 53248 31680
rect 54116 31628 54168 31680
rect 55404 31628 55456 31680
rect 67272 31628 67324 31680
rect 67548 31628 67600 31680
rect 68468 31671 68520 31680
rect 68468 31637 68477 31671
rect 68477 31637 68511 31671
rect 68511 31637 68520 31671
rect 68468 31628 68520 31637
rect 69020 31671 69072 31680
rect 69020 31637 69029 31671
rect 69029 31637 69063 31671
rect 69063 31637 69072 31671
rect 69020 31628 69072 31637
rect 80520 31628 80572 31680
rect 85120 31628 85172 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 65686 31526 65738 31578
rect 65750 31526 65802 31578
rect 65814 31526 65866 31578
rect 65878 31526 65930 31578
rect 96406 31526 96458 31578
rect 96470 31526 96522 31578
rect 96534 31526 96586 31578
rect 96598 31526 96650 31578
rect 17500 31424 17552 31476
rect 17960 31424 18012 31476
rect 4068 31356 4120 31408
rect 23664 31356 23716 31408
rect 7012 31288 7064 31340
rect 16120 31331 16172 31340
rect 16120 31297 16129 31331
rect 16129 31297 16163 31331
rect 16163 31297 16172 31331
rect 16120 31288 16172 31297
rect 16396 31288 16448 31340
rect 22744 31288 22796 31340
rect 25504 31356 25556 31408
rect 35256 31399 35308 31408
rect 35256 31365 35265 31399
rect 35265 31365 35299 31399
rect 35299 31365 35308 31399
rect 35256 31356 35308 31365
rect 41972 31399 42024 31408
rect 25412 31288 25464 31340
rect 35164 31288 35216 31340
rect 2964 31220 3016 31272
rect 4712 31220 4764 31272
rect 15660 31220 15712 31272
rect 17684 31220 17736 31272
rect 18328 31220 18380 31272
rect 24676 31263 24728 31272
rect 24676 31229 24685 31263
rect 24685 31229 24719 31263
rect 24719 31229 24728 31263
rect 24676 31220 24728 31229
rect 24952 31220 25004 31272
rect 15568 31195 15620 31204
rect 15568 31161 15577 31195
rect 15577 31161 15611 31195
rect 15611 31161 15620 31195
rect 15568 31152 15620 31161
rect 16488 31152 16540 31204
rect 17040 31152 17092 31204
rect 22744 31152 22796 31204
rect 24032 31195 24084 31204
rect 24032 31161 24041 31195
rect 24041 31161 24075 31195
rect 24075 31161 24084 31195
rect 24032 31152 24084 31161
rect 3516 31084 3568 31136
rect 4712 31127 4764 31136
rect 4712 31093 4721 31127
rect 4721 31093 4755 31127
rect 4755 31093 4764 31127
rect 4712 31084 4764 31093
rect 9588 31084 9640 31136
rect 12900 31084 12952 31136
rect 18328 31084 18380 31136
rect 24952 31084 25004 31136
rect 29460 31220 29512 31272
rect 41972 31365 41981 31399
rect 41981 31365 42015 31399
rect 42015 31365 42024 31399
rect 41972 31356 42024 31365
rect 35624 31288 35676 31340
rect 41236 31288 41288 31340
rect 41788 31288 41840 31340
rect 35900 31220 35952 31272
rect 36728 31263 36780 31272
rect 36728 31229 36737 31263
rect 36737 31229 36771 31263
rect 36771 31229 36780 31263
rect 36728 31220 36780 31229
rect 25412 31152 25464 31204
rect 29000 31084 29052 31136
rect 29460 31084 29512 31136
rect 30656 31084 30708 31136
rect 40776 31220 40828 31272
rect 38108 31195 38160 31204
rect 38108 31161 38117 31195
rect 38117 31161 38151 31195
rect 38151 31161 38160 31195
rect 38108 31152 38160 31161
rect 55404 31356 55456 31408
rect 61936 31424 61988 31476
rect 62120 31467 62172 31476
rect 62120 31433 62129 31467
rect 62129 31433 62163 31467
rect 62163 31433 62172 31467
rect 62120 31424 62172 31433
rect 63224 31467 63276 31476
rect 63224 31433 63233 31467
rect 63233 31433 63267 31467
rect 63267 31433 63276 31467
rect 63224 31424 63276 31433
rect 63592 31467 63644 31476
rect 63592 31433 63601 31467
rect 63601 31433 63635 31467
rect 63635 31433 63644 31467
rect 63592 31424 63644 31433
rect 68468 31424 68520 31476
rect 68836 31467 68888 31476
rect 68836 31433 68845 31467
rect 68845 31433 68879 31467
rect 68879 31433 68888 31467
rect 68836 31424 68888 31433
rect 75736 31467 75788 31476
rect 75736 31433 75745 31467
rect 75745 31433 75779 31467
rect 75779 31433 75788 31467
rect 75736 31424 75788 31433
rect 66904 31356 66956 31408
rect 68376 31356 68428 31408
rect 73620 31356 73672 31408
rect 43260 31288 43312 31340
rect 54944 31288 54996 31340
rect 37924 31084 37976 31136
rect 42064 31084 42116 31136
rect 42432 31084 42484 31136
rect 52368 31220 52420 31272
rect 53656 31263 53708 31272
rect 53656 31229 53665 31263
rect 53665 31229 53699 31263
rect 53699 31229 53708 31263
rect 53656 31220 53708 31229
rect 53840 31220 53892 31272
rect 54116 31263 54168 31272
rect 54116 31229 54125 31263
rect 54125 31229 54159 31263
rect 54159 31229 54168 31263
rect 54116 31220 54168 31229
rect 55036 31220 55088 31272
rect 59268 31220 59320 31272
rect 60464 31220 60516 31272
rect 60832 31263 60884 31272
rect 60832 31229 60841 31263
rect 60841 31229 60875 31263
rect 60875 31229 60884 31263
rect 60832 31220 60884 31229
rect 49240 31152 49292 31204
rect 57336 31152 57388 31204
rect 60280 31195 60332 31204
rect 60280 31161 60289 31195
rect 60289 31161 60323 31195
rect 60323 31161 60332 31195
rect 62120 31220 62172 31272
rect 60280 31152 60332 31161
rect 61936 31152 61988 31204
rect 62212 31152 62264 31204
rect 62396 31152 62448 31204
rect 67456 31152 67508 31204
rect 72516 31152 72568 31204
rect 45008 31084 45060 31136
rect 46940 31127 46992 31136
rect 46940 31093 46949 31127
rect 46949 31093 46983 31127
rect 46983 31093 46992 31127
rect 46940 31084 46992 31093
rect 53288 31084 53340 31136
rect 58440 31084 58492 31136
rect 60464 31127 60516 31136
rect 60464 31093 60473 31127
rect 60473 31093 60507 31127
rect 60507 31093 60516 31127
rect 60464 31084 60516 31093
rect 60832 31084 60884 31136
rect 62028 31084 62080 31136
rect 67180 31084 67232 31136
rect 69020 31084 69072 31136
rect 73620 31084 73672 31136
rect 76012 31424 76064 31476
rect 79600 31424 79652 31476
rect 82728 31356 82780 31408
rect 84200 31467 84252 31476
rect 84200 31433 84209 31467
rect 84209 31433 84243 31467
rect 84243 31433 84252 31467
rect 85120 31467 85172 31476
rect 84200 31424 84252 31433
rect 85120 31433 85129 31467
rect 85129 31433 85163 31467
rect 85163 31433 85172 31467
rect 85120 31424 85172 31433
rect 79784 31263 79836 31272
rect 79784 31229 79793 31263
rect 79793 31229 79827 31263
rect 79827 31229 79836 31263
rect 79784 31220 79836 31229
rect 79876 31220 79928 31272
rect 82360 31263 82412 31272
rect 82360 31229 82369 31263
rect 82369 31229 82403 31263
rect 82403 31229 82412 31263
rect 82360 31220 82412 31229
rect 82728 31263 82780 31272
rect 82728 31229 82737 31263
rect 82737 31229 82771 31263
rect 82771 31229 82780 31263
rect 82728 31220 82780 31229
rect 85028 31356 85080 31408
rect 87420 31263 87472 31272
rect 85396 31152 85448 31204
rect 87420 31229 87429 31263
rect 87429 31229 87463 31263
rect 87463 31229 87472 31263
rect 87420 31220 87472 31229
rect 87696 31263 87748 31272
rect 87696 31229 87705 31263
rect 87705 31229 87739 31263
rect 87739 31229 87748 31263
rect 87696 31220 87748 31229
rect 86684 31152 86736 31204
rect 88616 31152 88668 31204
rect 87420 31084 87472 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 50326 30982 50378 31034
rect 50390 30982 50442 31034
rect 50454 30982 50506 31034
rect 50518 30982 50570 31034
rect 81046 30982 81098 31034
rect 81110 30982 81162 31034
rect 81174 30982 81226 31034
rect 81238 30982 81290 31034
rect 11244 30812 11296 30864
rect 7748 30744 7800 30796
rect 12900 30880 12952 30932
rect 12992 30923 13044 30932
rect 12992 30889 13001 30923
rect 13001 30889 13035 30923
rect 13035 30889 13044 30923
rect 12992 30880 13044 30889
rect 17960 30880 18012 30932
rect 18236 30923 18288 30932
rect 18236 30889 18245 30923
rect 18245 30889 18279 30923
rect 18279 30889 18288 30923
rect 18236 30880 18288 30889
rect 25320 30880 25372 30932
rect 31024 30880 31076 30932
rect 31576 30880 31628 30932
rect 35164 30880 35216 30932
rect 11796 30787 11848 30796
rect 11796 30753 11805 30787
rect 11805 30753 11839 30787
rect 11839 30753 11848 30787
rect 12348 30812 12400 30864
rect 12440 30812 12492 30864
rect 12532 30812 12584 30864
rect 34796 30812 34848 30864
rect 36728 30855 36780 30864
rect 11796 30744 11848 30753
rect 12624 30787 12676 30796
rect 4712 30676 4764 30728
rect 11152 30676 11204 30728
rect 12624 30753 12633 30787
rect 12633 30753 12667 30787
rect 12667 30753 12676 30787
rect 12624 30744 12676 30753
rect 16120 30744 16172 30796
rect 16580 30744 16632 30796
rect 19984 30744 20036 30796
rect 24032 30787 24084 30796
rect 24032 30753 24041 30787
rect 24041 30753 24075 30787
rect 24075 30753 24084 30787
rect 24032 30744 24084 30753
rect 25320 30744 25372 30796
rect 35624 30787 35676 30796
rect 35624 30753 35633 30787
rect 35633 30753 35667 30787
rect 35667 30753 35676 30787
rect 35624 30744 35676 30753
rect 36360 30787 36412 30796
rect 36360 30753 36369 30787
rect 36369 30753 36403 30787
rect 36403 30753 36412 30787
rect 36360 30744 36412 30753
rect 16488 30719 16540 30728
rect 16488 30685 16497 30719
rect 16497 30685 16531 30719
rect 16531 30685 16540 30719
rect 16488 30676 16540 30685
rect 29092 30719 29144 30728
rect 29092 30685 29101 30719
rect 29101 30685 29135 30719
rect 29135 30685 29144 30719
rect 29092 30676 29144 30685
rect 29276 30676 29328 30728
rect 36728 30821 36737 30855
rect 36737 30821 36771 30855
rect 36771 30821 36780 30855
rect 36728 30812 36780 30821
rect 57336 30880 57388 30932
rect 41604 30812 41656 30864
rect 41788 30812 41840 30864
rect 37188 30744 37240 30796
rect 37556 30676 37608 30728
rect 12532 30608 12584 30660
rect 4068 30540 4120 30592
rect 6644 30583 6696 30592
rect 6644 30549 6653 30583
rect 6653 30549 6687 30583
rect 6687 30549 6696 30583
rect 6644 30540 6696 30549
rect 11704 30540 11756 30592
rect 15384 30608 15436 30660
rect 30656 30651 30708 30660
rect 30656 30617 30665 30651
rect 30665 30617 30699 30651
rect 30699 30617 30708 30651
rect 30656 30608 30708 30617
rect 17408 30540 17460 30592
rect 19892 30540 19944 30592
rect 24124 30583 24176 30592
rect 24124 30549 24133 30583
rect 24133 30549 24167 30583
rect 24167 30549 24176 30583
rect 24124 30540 24176 30549
rect 36360 30540 36412 30592
rect 37464 30583 37516 30592
rect 37464 30549 37473 30583
rect 37473 30549 37507 30583
rect 37507 30549 37516 30583
rect 37464 30540 37516 30549
rect 38016 30676 38068 30728
rect 38660 30744 38712 30796
rect 40960 30787 41012 30796
rect 40960 30753 40969 30787
rect 40969 30753 41003 30787
rect 41003 30753 41012 30787
rect 40960 30744 41012 30753
rect 41696 30787 41748 30796
rect 40776 30719 40828 30728
rect 40776 30685 40785 30719
rect 40785 30685 40819 30719
rect 40819 30685 40828 30719
rect 40776 30676 40828 30685
rect 38292 30608 38344 30660
rect 40500 30651 40552 30660
rect 40500 30617 40509 30651
rect 40509 30617 40543 30651
rect 40543 30617 40552 30651
rect 40500 30608 40552 30617
rect 41696 30753 41705 30787
rect 41705 30753 41739 30787
rect 41739 30753 41748 30787
rect 41696 30744 41748 30753
rect 41880 30787 41932 30796
rect 41880 30753 41889 30787
rect 41889 30753 41923 30787
rect 41923 30753 41932 30787
rect 42432 30787 42484 30796
rect 41880 30744 41932 30753
rect 42432 30753 42441 30787
rect 42441 30753 42475 30787
rect 42475 30753 42484 30787
rect 42432 30744 42484 30753
rect 43168 30744 43220 30796
rect 43536 30744 43588 30796
rect 49240 30787 49292 30796
rect 43628 30676 43680 30728
rect 41604 30608 41656 30660
rect 48504 30676 48556 30728
rect 46940 30608 46992 30660
rect 38660 30540 38712 30592
rect 43260 30540 43312 30592
rect 43444 30583 43496 30592
rect 43444 30549 43453 30583
rect 43453 30549 43487 30583
rect 43487 30549 43496 30583
rect 43444 30540 43496 30549
rect 43536 30540 43588 30592
rect 47492 30608 47544 30660
rect 49240 30753 49249 30787
rect 49249 30753 49283 30787
rect 49283 30753 49292 30787
rect 49240 30744 49292 30753
rect 54024 30744 54076 30796
rect 56232 30787 56284 30796
rect 56232 30753 56241 30787
rect 56241 30753 56275 30787
rect 56275 30753 56284 30787
rect 56232 30744 56284 30753
rect 58716 30744 58768 30796
rect 54116 30676 54168 30728
rect 56600 30719 56652 30728
rect 56600 30685 56609 30719
rect 56609 30685 56643 30719
rect 56643 30685 56652 30719
rect 56600 30676 56652 30685
rect 57796 30651 57848 30660
rect 57796 30617 57805 30651
rect 57805 30617 57839 30651
rect 57839 30617 57848 30651
rect 57796 30608 57848 30617
rect 59176 30880 59228 30932
rect 60924 30676 60976 30728
rect 62212 30880 62264 30932
rect 67456 30923 67508 30932
rect 62396 30855 62448 30864
rect 61660 30744 61712 30796
rect 61936 30787 61988 30796
rect 61936 30753 61941 30787
rect 61941 30753 61975 30787
rect 61975 30753 61988 30787
rect 61936 30744 61988 30753
rect 62396 30821 62405 30855
rect 62405 30821 62439 30855
rect 62439 30821 62448 30855
rect 62396 30812 62448 30821
rect 67456 30889 67465 30923
rect 67465 30889 67499 30923
rect 67499 30889 67508 30923
rect 67456 30880 67508 30889
rect 67548 30880 67600 30932
rect 66996 30787 67048 30796
rect 66996 30753 67005 30787
rect 67005 30753 67039 30787
rect 67039 30753 67048 30787
rect 66996 30744 67048 30753
rect 67732 30744 67784 30796
rect 68008 30676 68060 30728
rect 69480 30880 69532 30932
rect 69756 30880 69808 30932
rect 84660 30880 84712 30932
rect 85120 30880 85172 30932
rect 87972 30923 88024 30932
rect 70032 30812 70084 30864
rect 72516 30812 72568 30864
rect 69204 30787 69256 30796
rect 69204 30753 69213 30787
rect 69213 30753 69247 30787
rect 69247 30753 69256 30787
rect 69204 30744 69256 30753
rect 73712 30787 73764 30796
rect 73712 30753 73721 30787
rect 73721 30753 73755 30787
rect 73755 30753 73764 30787
rect 73712 30744 73764 30753
rect 73160 30676 73212 30728
rect 74264 30787 74316 30796
rect 74264 30753 74273 30787
rect 74273 30753 74307 30787
rect 74307 30753 74316 30787
rect 76012 30812 76064 30864
rect 82820 30812 82872 30864
rect 83188 30812 83240 30864
rect 83924 30812 83976 30864
rect 87972 30889 87981 30923
rect 87981 30889 88015 30923
rect 88015 30889 88024 30923
rect 87972 30880 88024 30889
rect 88248 30880 88300 30932
rect 74264 30744 74316 30753
rect 79600 30787 79652 30796
rect 79600 30753 79609 30787
rect 79609 30753 79643 30787
rect 79643 30753 79652 30787
rect 79876 30787 79928 30796
rect 79600 30744 79652 30753
rect 79876 30753 79885 30787
rect 79885 30753 79919 30787
rect 79919 30753 79928 30787
rect 80888 30787 80940 30796
rect 79876 30744 79928 30753
rect 79784 30676 79836 30728
rect 69664 30608 69716 30660
rect 80888 30753 80897 30787
rect 80897 30753 80931 30787
rect 80931 30753 80940 30787
rect 80888 30744 80940 30753
rect 84200 30787 84252 30796
rect 84200 30753 84209 30787
rect 84209 30753 84243 30787
rect 84243 30753 84252 30787
rect 86592 30787 86644 30796
rect 84200 30744 84252 30753
rect 86592 30753 86601 30787
rect 86601 30753 86635 30787
rect 86635 30753 86644 30787
rect 86592 30744 86644 30753
rect 88616 30787 88668 30796
rect 88616 30753 88625 30787
rect 88625 30753 88659 30787
rect 88659 30753 88668 30787
rect 88616 30744 88668 30753
rect 80704 30719 80756 30728
rect 80704 30685 80713 30719
rect 80713 30685 80747 30719
rect 80747 30685 80756 30719
rect 83924 30719 83976 30728
rect 80704 30676 80756 30685
rect 83924 30685 83933 30719
rect 83933 30685 83967 30719
rect 83967 30685 83976 30719
rect 83924 30676 83976 30685
rect 82360 30608 82412 30660
rect 47216 30540 47268 30592
rect 48780 30583 48832 30592
rect 48780 30549 48789 30583
rect 48789 30549 48823 30583
rect 48823 30549 48832 30583
rect 48780 30540 48832 30549
rect 50160 30540 50212 30592
rect 54668 30583 54720 30592
rect 54668 30549 54677 30583
rect 54677 30549 54711 30583
rect 54711 30549 54720 30583
rect 54668 30540 54720 30549
rect 59084 30540 59136 30592
rect 59176 30583 59228 30592
rect 59176 30549 59185 30583
rect 59185 30549 59219 30583
rect 59219 30549 59228 30583
rect 59176 30540 59228 30549
rect 60372 30540 60424 30592
rect 61660 30540 61712 30592
rect 61936 30540 61988 30592
rect 66996 30540 67048 30592
rect 67732 30583 67784 30592
rect 67732 30549 67741 30583
rect 67741 30549 67775 30583
rect 67775 30549 67784 30583
rect 67732 30540 67784 30549
rect 68008 30583 68060 30592
rect 68008 30549 68017 30583
rect 68017 30549 68051 30583
rect 68051 30549 68060 30583
rect 68008 30540 68060 30549
rect 69756 30540 69808 30592
rect 70032 30583 70084 30592
rect 70032 30549 70041 30583
rect 70041 30549 70075 30583
rect 70075 30549 70084 30583
rect 70032 30540 70084 30549
rect 73160 30583 73212 30592
rect 73160 30549 73169 30583
rect 73169 30549 73203 30583
rect 73203 30549 73212 30583
rect 73160 30540 73212 30549
rect 79232 30540 79284 30592
rect 85304 30583 85356 30592
rect 85304 30549 85313 30583
rect 85313 30549 85347 30583
rect 85347 30549 85356 30583
rect 85304 30540 85356 30549
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 65686 30438 65738 30490
rect 65750 30438 65802 30490
rect 65814 30438 65866 30490
rect 65878 30438 65930 30490
rect 96406 30438 96458 30490
rect 96470 30438 96522 30490
rect 96534 30438 96586 30490
rect 96598 30438 96650 30490
rect 3608 30336 3660 30388
rect 4896 30336 4948 30388
rect 10692 30336 10744 30388
rect 16488 30336 16540 30388
rect 31024 30379 31076 30388
rect 31024 30345 31033 30379
rect 31033 30345 31067 30379
rect 31067 30345 31076 30379
rect 31024 30336 31076 30345
rect 37464 30336 37516 30388
rect 3884 30268 3936 30320
rect 20076 30268 20128 30320
rect 2964 30200 3016 30252
rect 4712 30200 4764 30252
rect 9588 30132 9640 30184
rect 18512 30200 18564 30252
rect 26792 30268 26844 30320
rect 29276 30268 29328 30320
rect 9956 30064 10008 30116
rect 3148 29996 3200 30048
rect 4436 30039 4488 30048
rect 4436 30005 4445 30039
rect 4445 30005 4479 30039
rect 4479 30005 4488 30039
rect 4436 29996 4488 30005
rect 7748 30039 7800 30048
rect 7748 30005 7757 30039
rect 7757 30005 7791 30039
rect 7791 30005 7800 30039
rect 7748 29996 7800 30005
rect 9680 29996 9732 30048
rect 10692 29996 10744 30048
rect 11152 30132 11204 30184
rect 12624 30132 12676 30184
rect 15568 30132 15620 30184
rect 19984 30132 20036 30184
rect 22468 30200 22520 30252
rect 24676 30200 24728 30252
rect 24768 30175 24820 30184
rect 11704 29996 11756 30048
rect 11888 30039 11940 30048
rect 11888 30005 11897 30039
rect 11897 30005 11931 30039
rect 11931 30005 11940 30039
rect 11888 29996 11940 30005
rect 15568 30039 15620 30048
rect 15568 30005 15577 30039
rect 15577 30005 15611 30039
rect 15611 30005 15620 30039
rect 15568 29996 15620 30005
rect 19984 30039 20036 30048
rect 19984 30005 19993 30039
rect 19993 30005 20027 30039
rect 20027 30005 20036 30039
rect 19984 29996 20036 30005
rect 20812 29996 20864 30048
rect 20904 29996 20956 30048
rect 22284 30107 22336 30116
rect 22284 30073 22293 30107
rect 22293 30073 22327 30107
rect 22327 30073 22336 30107
rect 22284 30064 22336 30073
rect 24768 30141 24777 30175
rect 24777 30141 24811 30175
rect 24811 30141 24820 30175
rect 24768 30132 24820 30141
rect 24952 30175 25004 30184
rect 24952 30141 24961 30175
rect 24961 30141 24995 30175
rect 24995 30141 25004 30175
rect 24952 30132 25004 30141
rect 26332 30132 26384 30184
rect 27160 30175 27212 30184
rect 22468 30039 22520 30048
rect 22468 30005 22477 30039
rect 22477 30005 22511 30039
rect 22511 30005 22520 30039
rect 22468 29996 22520 30005
rect 23296 29996 23348 30048
rect 23664 29996 23716 30048
rect 27160 30141 27169 30175
rect 27169 30141 27203 30175
rect 27203 30141 27212 30175
rect 27160 30132 27212 30141
rect 27252 30132 27304 30184
rect 27804 30175 27856 30184
rect 27804 30141 27809 30175
rect 27809 30141 27843 30175
rect 27843 30141 27856 30175
rect 27804 30132 27856 30141
rect 27252 29996 27304 30048
rect 29000 30200 29052 30252
rect 29092 30200 29144 30252
rect 37556 30311 37608 30320
rect 37556 30277 37565 30311
rect 37565 30277 37599 30311
rect 37599 30277 37608 30311
rect 37556 30268 37608 30277
rect 43168 30311 43220 30320
rect 43168 30277 43177 30311
rect 43177 30277 43211 30311
rect 43211 30277 43220 30311
rect 43168 30268 43220 30277
rect 48780 30311 48832 30320
rect 48780 30277 48789 30311
rect 48789 30277 48823 30311
rect 48823 30277 48832 30311
rect 48780 30268 48832 30277
rect 54024 30336 54076 30388
rect 60464 30336 60516 30388
rect 60924 30336 60976 30388
rect 29368 30132 29420 30184
rect 29644 30132 29696 30184
rect 52644 30200 52696 30252
rect 35716 30132 35768 30184
rect 37280 30132 37332 30184
rect 37464 30175 37516 30184
rect 37464 30141 37473 30175
rect 37473 30141 37507 30175
rect 37507 30141 37516 30175
rect 37464 30132 37516 30141
rect 37924 30132 37976 30184
rect 38016 30132 38068 30184
rect 41604 30175 41656 30184
rect 41604 30141 41613 30175
rect 41613 30141 41647 30175
rect 41647 30141 41656 30175
rect 41604 30132 41656 30141
rect 42248 30132 42300 30184
rect 43352 30175 43404 30184
rect 43352 30141 43361 30175
rect 43361 30141 43395 30175
rect 43395 30141 43404 30175
rect 43352 30132 43404 30141
rect 43628 30175 43680 30184
rect 43628 30141 43637 30175
rect 43637 30141 43671 30175
rect 43671 30141 43680 30175
rect 43628 30132 43680 30141
rect 44732 30132 44784 30184
rect 45468 30132 45520 30184
rect 46940 30175 46992 30184
rect 46940 30141 46949 30175
rect 46949 30141 46983 30175
rect 46983 30141 46992 30175
rect 46940 30132 46992 30141
rect 47216 30175 47268 30184
rect 47216 30141 47225 30175
rect 47225 30141 47259 30175
rect 47259 30141 47268 30175
rect 47216 30132 47268 30141
rect 47308 30132 47360 30184
rect 48780 30132 48832 30184
rect 45008 30107 45060 30116
rect 28724 30039 28776 30048
rect 28724 30005 28733 30039
rect 28733 30005 28767 30039
rect 28767 30005 28776 30039
rect 28724 29996 28776 30005
rect 29828 29996 29880 30048
rect 30840 30039 30892 30048
rect 30840 30005 30849 30039
rect 30849 30005 30883 30039
rect 30883 30005 30892 30039
rect 37004 30039 37056 30048
rect 30840 29996 30892 30005
rect 37004 30005 37013 30039
rect 37013 30005 37047 30039
rect 37047 30005 37056 30039
rect 37004 29996 37056 30005
rect 37924 30039 37976 30048
rect 37924 30005 37933 30039
rect 37933 30005 37967 30039
rect 37967 30005 37976 30039
rect 37924 29996 37976 30005
rect 45008 30073 45017 30107
rect 45017 30073 45051 30107
rect 45051 30073 45060 30107
rect 45008 30064 45060 30073
rect 46848 30064 46900 30116
rect 58716 30200 58768 30252
rect 59176 30200 59228 30252
rect 53012 30175 53064 30184
rect 53012 30141 53021 30175
rect 53021 30141 53055 30175
rect 53055 30141 53064 30175
rect 53012 30132 53064 30141
rect 53288 30132 53340 30184
rect 56784 30132 56836 30184
rect 48320 30039 48372 30048
rect 48320 30005 48329 30039
rect 48329 30005 48363 30039
rect 48363 30005 48372 30039
rect 48320 29996 48372 30005
rect 52000 29996 52052 30048
rect 56600 29996 56652 30048
rect 57796 30132 57848 30184
rect 59452 30132 59504 30184
rect 60372 30175 60424 30184
rect 60372 30141 60381 30175
rect 60381 30141 60415 30175
rect 60415 30141 60424 30175
rect 60372 30132 60424 30141
rect 60188 30064 60240 30116
rect 59360 29996 59412 30048
rect 60004 30039 60056 30048
rect 60004 30005 60013 30039
rect 60013 30005 60047 30039
rect 60047 30005 60056 30039
rect 60004 29996 60056 30005
rect 60648 29996 60700 30048
rect 61108 30268 61160 30320
rect 61936 30311 61988 30320
rect 61936 30277 61945 30311
rect 61945 30277 61979 30311
rect 61979 30277 61988 30311
rect 61936 30268 61988 30277
rect 67732 30336 67784 30388
rect 69664 30336 69716 30388
rect 70032 30336 70084 30388
rect 80704 30336 80756 30388
rect 84660 30379 84712 30388
rect 84660 30345 84669 30379
rect 84669 30345 84703 30379
rect 84703 30345 84712 30379
rect 84660 30336 84712 30345
rect 85304 30336 85356 30388
rect 62028 30175 62080 30184
rect 60832 30064 60884 30116
rect 62028 30141 62037 30175
rect 62037 30141 62071 30175
rect 62071 30141 62080 30175
rect 62028 30132 62080 30141
rect 66076 30200 66128 30252
rect 71596 30268 71648 30320
rect 85120 30268 85172 30320
rect 67088 30132 67140 30184
rect 68836 30132 68888 30184
rect 73160 30200 73212 30252
rect 74356 30175 74408 30184
rect 74356 30141 74365 30175
rect 74365 30141 74399 30175
rect 74399 30141 74408 30175
rect 74356 30132 74408 30141
rect 80060 30175 80112 30184
rect 75920 30064 75972 30116
rect 80060 30141 80069 30175
rect 80069 30141 80103 30175
rect 80103 30141 80112 30175
rect 80060 30132 80112 30141
rect 84660 30132 84712 30184
rect 85396 30132 85448 30184
rect 86592 30200 86644 30252
rect 86684 30175 86736 30184
rect 86684 30141 86693 30175
rect 86693 30141 86727 30175
rect 86727 30141 86736 30175
rect 86684 30132 86736 30141
rect 88248 30132 88300 30184
rect 86960 30107 87012 30116
rect 86960 30073 86969 30107
rect 86969 30073 87003 30107
rect 87003 30073 87012 30107
rect 86960 30064 87012 30073
rect 66076 30039 66128 30048
rect 66076 30005 66085 30039
rect 66085 30005 66119 30039
rect 66119 30005 66128 30039
rect 66076 29996 66128 30005
rect 67916 29996 67968 30048
rect 68836 30039 68888 30048
rect 68836 30005 68845 30039
rect 68845 30005 68879 30039
rect 68879 30005 68888 30039
rect 68836 29996 68888 30005
rect 73160 29996 73212 30048
rect 80520 29996 80572 30048
rect 87052 30039 87104 30048
rect 87052 30005 87061 30039
rect 87061 30005 87095 30039
rect 87095 30005 87104 30039
rect 87052 29996 87104 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 50326 29894 50378 29946
rect 50390 29894 50442 29946
rect 50454 29894 50506 29946
rect 50518 29894 50570 29946
rect 81046 29894 81098 29946
rect 81110 29894 81162 29946
rect 81174 29894 81226 29946
rect 81238 29894 81290 29946
rect 4436 29792 4488 29844
rect 13452 29792 13504 29844
rect 15384 29792 15436 29844
rect 17960 29835 18012 29844
rect 17960 29801 17969 29835
rect 17969 29801 18003 29835
rect 18003 29801 18012 29835
rect 17960 29792 18012 29801
rect 18236 29792 18288 29844
rect 19248 29792 19300 29844
rect 27160 29792 27212 29844
rect 6644 29724 6696 29776
rect 7748 29724 7800 29776
rect 4712 29699 4764 29708
rect 4712 29665 4721 29699
rect 4721 29665 4755 29699
rect 4755 29665 4764 29699
rect 4712 29656 4764 29665
rect 8484 29656 8536 29708
rect 9680 29699 9732 29708
rect 9680 29665 9689 29699
rect 9689 29665 9723 29699
rect 9723 29665 9732 29699
rect 9956 29699 10008 29708
rect 9680 29656 9732 29665
rect 9956 29665 9965 29699
rect 9965 29665 9999 29699
rect 9999 29665 10008 29699
rect 9956 29656 10008 29665
rect 11888 29656 11940 29708
rect 15568 29656 15620 29708
rect 16120 29656 16172 29708
rect 18328 29724 18380 29776
rect 23664 29724 23716 29776
rect 26792 29767 26844 29776
rect 26792 29733 26801 29767
rect 26801 29733 26835 29767
rect 26835 29733 26844 29767
rect 26792 29724 26844 29733
rect 19984 29656 20036 29708
rect 24124 29656 24176 29708
rect 27804 29792 27856 29844
rect 29368 29792 29420 29844
rect 29828 29792 29880 29844
rect 36544 29792 36596 29844
rect 37464 29792 37516 29844
rect 40960 29835 41012 29844
rect 40960 29801 40969 29835
rect 40969 29801 41003 29835
rect 41003 29801 41012 29835
rect 40960 29792 41012 29801
rect 41788 29792 41840 29844
rect 42064 29792 42116 29844
rect 42248 29835 42300 29844
rect 42248 29801 42257 29835
rect 42257 29801 42291 29835
rect 42291 29801 42300 29835
rect 42248 29792 42300 29801
rect 42800 29792 42852 29844
rect 43444 29792 43496 29844
rect 47492 29792 47544 29844
rect 52644 29792 52696 29844
rect 53012 29792 53064 29844
rect 19248 29588 19300 29640
rect 24032 29588 24084 29640
rect 26148 29588 26200 29640
rect 26884 29588 26936 29640
rect 27804 29656 27856 29708
rect 28724 29699 28776 29708
rect 28724 29665 28733 29699
rect 28733 29665 28767 29699
rect 28767 29665 28776 29699
rect 28724 29656 28776 29665
rect 30840 29724 30892 29776
rect 45284 29724 45336 29776
rect 28172 29588 28224 29640
rect 37004 29656 37056 29708
rect 37280 29656 37332 29708
rect 38292 29656 38344 29708
rect 40960 29656 41012 29708
rect 41236 29699 41288 29708
rect 41236 29665 41245 29699
rect 41245 29665 41279 29699
rect 41279 29665 41288 29699
rect 41236 29656 41288 29665
rect 41788 29699 41840 29708
rect 41788 29665 41797 29699
rect 41797 29665 41831 29699
rect 41831 29665 41840 29699
rect 41788 29656 41840 29665
rect 42800 29656 42852 29708
rect 42248 29588 42300 29640
rect 44180 29588 44232 29640
rect 46848 29724 46900 29776
rect 47032 29699 47084 29708
rect 47032 29665 47041 29699
rect 47041 29665 47075 29699
rect 47075 29665 47084 29699
rect 47032 29656 47084 29665
rect 2780 29520 2832 29572
rect 3240 29520 3292 29572
rect 17316 29520 17368 29572
rect 4068 29452 4120 29504
rect 9680 29452 9732 29504
rect 24584 29520 24636 29572
rect 18696 29452 18748 29504
rect 24768 29452 24820 29504
rect 26332 29452 26384 29504
rect 26424 29452 26476 29504
rect 29276 29452 29328 29504
rect 29460 29520 29512 29572
rect 40500 29520 40552 29572
rect 45376 29588 45428 29640
rect 45560 29588 45612 29640
rect 50988 29656 51040 29708
rect 52736 29656 52788 29708
rect 52000 29631 52052 29640
rect 52000 29597 52009 29631
rect 52009 29597 52043 29631
rect 52043 29597 52052 29631
rect 52000 29588 52052 29597
rect 53104 29656 53156 29708
rect 60556 29792 60608 29844
rect 67640 29792 67692 29844
rect 53196 29588 53248 29640
rect 54668 29588 54720 29640
rect 48044 29563 48096 29572
rect 48044 29529 48053 29563
rect 48053 29529 48087 29563
rect 48087 29529 48096 29563
rect 48044 29520 48096 29529
rect 48136 29520 48188 29572
rect 55496 29699 55548 29708
rect 55496 29665 55505 29699
rect 55505 29665 55539 29699
rect 55539 29665 55548 29699
rect 55496 29656 55548 29665
rect 56784 29699 56836 29708
rect 56784 29665 56793 29699
rect 56793 29665 56827 29699
rect 56827 29665 56836 29699
rect 56784 29656 56836 29665
rect 57888 29699 57940 29708
rect 57888 29665 57897 29699
rect 57897 29665 57931 29699
rect 57931 29665 57940 29699
rect 58440 29699 58492 29708
rect 57888 29656 57940 29665
rect 58440 29665 58449 29699
rect 58449 29665 58483 29699
rect 58483 29665 58492 29699
rect 58440 29656 58492 29665
rect 61292 29724 61344 29776
rect 60556 29656 60608 29708
rect 67916 29699 67968 29708
rect 59636 29588 59688 29640
rect 60188 29631 60240 29640
rect 60188 29597 60197 29631
rect 60197 29597 60231 29631
rect 60231 29597 60240 29631
rect 60188 29588 60240 29597
rect 67640 29631 67692 29640
rect 67640 29597 67649 29631
rect 67649 29597 67683 29631
rect 67683 29597 67692 29631
rect 67640 29588 67692 29597
rect 67916 29665 67925 29699
rect 67925 29665 67959 29699
rect 67959 29665 67968 29699
rect 67916 29656 67968 29665
rect 69480 29792 69532 29844
rect 73160 29835 73212 29844
rect 73160 29801 73169 29835
rect 73169 29801 73203 29835
rect 73203 29801 73212 29835
rect 73160 29792 73212 29801
rect 74356 29792 74408 29844
rect 80060 29792 80112 29844
rect 80704 29792 80756 29844
rect 79232 29699 79284 29708
rect 79232 29665 79241 29699
rect 79241 29665 79275 29699
rect 79275 29665 79284 29699
rect 79232 29656 79284 29665
rect 80520 29699 80572 29708
rect 80520 29665 80529 29699
rect 80529 29665 80563 29699
rect 80563 29665 80572 29699
rect 80520 29656 80572 29665
rect 71596 29631 71648 29640
rect 71596 29597 71605 29631
rect 71605 29597 71639 29631
rect 71639 29597 71648 29631
rect 71596 29588 71648 29597
rect 55312 29563 55364 29572
rect 55312 29529 55321 29563
rect 55321 29529 55355 29563
rect 55355 29529 55364 29563
rect 59084 29563 59136 29572
rect 55312 29520 55364 29529
rect 59084 29529 59093 29563
rect 59093 29529 59127 29563
rect 59127 29529 59136 29563
rect 59084 29520 59136 29529
rect 59544 29563 59596 29572
rect 59544 29529 59553 29563
rect 59553 29529 59587 29563
rect 59587 29529 59596 29563
rect 59544 29520 59596 29529
rect 35900 29452 35952 29504
rect 41604 29452 41656 29504
rect 43352 29452 43404 29504
rect 45376 29495 45428 29504
rect 45376 29461 45385 29495
rect 45385 29461 45419 29495
rect 45419 29461 45428 29495
rect 45376 29452 45428 29461
rect 46204 29452 46256 29504
rect 48872 29452 48924 29504
rect 48964 29452 49016 29504
rect 53564 29452 53616 29504
rect 58716 29452 58768 29504
rect 58992 29452 59044 29504
rect 59176 29495 59228 29504
rect 59176 29461 59185 29495
rect 59185 29461 59219 29495
rect 59219 29461 59228 29495
rect 59176 29452 59228 29461
rect 59728 29495 59780 29504
rect 59728 29461 59737 29495
rect 59737 29461 59771 29495
rect 59771 29461 59780 29495
rect 59728 29452 59780 29461
rect 59912 29495 59964 29504
rect 59912 29461 59921 29495
rect 59921 29461 59955 29495
rect 59955 29461 59964 29495
rect 59912 29452 59964 29461
rect 75920 29588 75972 29640
rect 82912 29520 82964 29572
rect 83924 29520 83976 29572
rect 87144 29563 87196 29572
rect 87144 29529 87153 29563
rect 87153 29529 87187 29563
rect 87187 29529 87196 29563
rect 87144 29520 87196 29529
rect 61292 29452 61344 29504
rect 61568 29495 61620 29504
rect 61568 29461 61577 29495
rect 61577 29461 61611 29495
rect 61611 29461 61620 29495
rect 61568 29452 61620 29461
rect 67916 29452 67968 29504
rect 68836 29452 68888 29504
rect 86316 29495 86368 29504
rect 86316 29461 86325 29495
rect 86325 29461 86359 29495
rect 86359 29461 86368 29495
rect 86316 29452 86368 29461
rect 86500 29495 86552 29504
rect 86500 29461 86509 29495
rect 86509 29461 86543 29495
rect 86543 29461 86552 29495
rect 86500 29452 86552 29461
rect 86592 29452 86644 29504
rect 87236 29495 87288 29504
rect 87236 29461 87245 29495
rect 87245 29461 87279 29495
rect 87279 29461 87288 29495
rect 87236 29452 87288 29461
rect 87420 29495 87472 29504
rect 87420 29461 87429 29495
rect 87429 29461 87463 29495
rect 87463 29461 87472 29495
rect 87420 29452 87472 29461
rect 87604 29495 87656 29504
rect 87604 29461 87613 29495
rect 87613 29461 87647 29495
rect 87647 29461 87656 29495
rect 87604 29452 87656 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 65686 29350 65738 29402
rect 65750 29350 65802 29402
rect 65814 29350 65866 29402
rect 65878 29350 65930 29402
rect 96406 29350 96458 29402
rect 96470 29350 96522 29402
rect 96534 29350 96586 29402
rect 96598 29350 96650 29402
rect 2596 29112 2648 29164
rect 4712 29248 4764 29300
rect 4896 29248 4948 29300
rect 3056 29155 3108 29164
rect 3056 29121 3065 29155
rect 3065 29121 3099 29155
rect 3099 29121 3108 29155
rect 3056 29112 3108 29121
rect 3424 29112 3476 29164
rect 11888 29112 11940 29164
rect 23020 29248 23072 29300
rect 23112 29248 23164 29300
rect 46204 29248 46256 29300
rect 47032 29248 47084 29300
rect 55496 29248 55548 29300
rect 56784 29248 56836 29300
rect 66076 29248 66128 29300
rect 20904 29180 20956 29232
rect 12348 29044 12400 29096
rect 14924 29044 14976 29096
rect 13268 28976 13320 29028
rect 14004 28976 14056 29028
rect 16580 29044 16632 29096
rect 19340 29044 19392 29096
rect 20720 29112 20772 29164
rect 24584 29180 24636 29232
rect 25044 29180 25096 29232
rect 25320 29180 25372 29232
rect 25504 29180 25556 29232
rect 52000 29180 52052 29232
rect 52644 29180 52696 29232
rect 60004 29180 60056 29232
rect 63500 29180 63552 29232
rect 69480 29180 69532 29232
rect 17500 28976 17552 29028
rect 14832 28951 14884 28960
rect 14832 28917 14841 28951
rect 14841 28917 14875 28951
rect 14875 28917 14884 28951
rect 14832 28908 14884 28917
rect 14924 28951 14976 28960
rect 14924 28917 14933 28951
rect 14933 28917 14967 28951
rect 14967 28917 14976 28951
rect 20444 28976 20496 29028
rect 14924 28908 14976 28917
rect 25044 29044 25096 29096
rect 25136 29044 25188 29096
rect 20904 28976 20956 29028
rect 20812 28908 20864 28960
rect 23296 28908 23348 28960
rect 23940 28908 23992 28960
rect 25596 29112 25648 29164
rect 25412 29044 25464 29096
rect 29460 29044 29512 29096
rect 35440 29112 35492 29164
rect 42800 29112 42852 29164
rect 45376 29112 45428 29164
rect 53840 29112 53892 29164
rect 59268 29112 59320 29164
rect 61568 29112 61620 29164
rect 73620 29112 73672 29164
rect 50988 28976 51040 29028
rect 57796 28976 57848 29028
rect 59728 28976 59780 29028
rect 53564 28908 53616 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 4620 28704 4672 28756
rect 9588 28704 9640 28756
rect 3976 28636 4028 28688
rect 15108 28704 15160 28756
rect 15384 28747 15436 28756
rect 15384 28713 15393 28747
rect 15393 28713 15427 28747
rect 15427 28713 15436 28747
rect 15384 28704 15436 28713
rect 19340 28704 19392 28756
rect 20904 28704 20956 28756
rect 4620 28568 4672 28620
rect 2964 28500 3016 28552
rect 5080 28500 5132 28552
rect 8300 28568 8352 28620
rect 10692 28568 10744 28620
rect 13820 28611 13872 28620
rect 13820 28577 13829 28611
rect 13829 28577 13863 28611
rect 13863 28577 13872 28611
rect 13820 28568 13872 28577
rect 13912 28611 13964 28620
rect 13912 28577 13921 28611
rect 13921 28577 13955 28611
rect 13955 28577 13964 28611
rect 13912 28568 13964 28577
rect 14004 28500 14056 28552
rect 14096 28500 14148 28552
rect 8208 28432 8260 28484
rect 14832 28568 14884 28620
rect 15752 28611 15804 28620
rect 15752 28577 15761 28611
rect 15761 28577 15795 28611
rect 15795 28577 15804 28611
rect 15752 28568 15804 28577
rect 17868 28568 17920 28620
rect 15292 28500 15344 28552
rect 23664 28500 23716 28552
rect 37924 28432 37976 28484
rect 4620 28364 4672 28416
rect 8300 28407 8352 28416
rect 8300 28373 8309 28407
rect 8309 28373 8343 28407
rect 8343 28373 8352 28407
rect 8300 28364 8352 28373
rect 9864 28407 9916 28416
rect 9864 28373 9873 28407
rect 9873 28373 9907 28407
rect 9907 28373 9916 28407
rect 9864 28364 9916 28373
rect 12716 28364 12768 28416
rect 25228 28364 25280 28416
rect 26240 28364 26292 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 9588 28160 9640 28212
rect 2596 28067 2648 28076
rect 2596 28033 2605 28067
rect 2605 28033 2639 28067
rect 2639 28033 2648 28067
rect 2596 28024 2648 28033
rect 3516 28024 3568 28076
rect 11060 28160 11112 28212
rect 16396 28160 16448 28212
rect 17868 28160 17920 28212
rect 20260 28203 20312 28212
rect 20260 28169 20269 28203
rect 20269 28169 20303 28203
rect 20303 28169 20312 28203
rect 20260 28160 20312 28169
rect 21180 28203 21232 28212
rect 21180 28169 21189 28203
rect 21189 28169 21223 28203
rect 21223 28169 21232 28203
rect 21180 28160 21232 28169
rect 24952 28160 25004 28212
rect 25596 28160 25648 28212
rect 9864 28092 9916 28144
rect 13820 28092 13872 28144
rect 14924 28092 14976 28144
rect 10692 28067 10744 28076
rect 10692 28033 10701 28067
rect 10701 28033 10735 28067
rect 10735 28033 10744 28067
rect 10692 28024 10744 28033
rect 13912 28024 13964 28076
rect 14464 28024 14516 28076
rect 2964 27820 3016 27872
rect 4896 27820 4948 27872
rect 10140 27956 10192 28008
rect 14280 27956 14332 28008
rect 12624 27888 12676 27940
rect 14004 27888 14056 27940
rect 14464 27931 14516 27940
rect 14464 27897 14473 27931
rect 14473 27897 14507 27931
rect 14507 27897 14516 27931
rect 14464 27888 14516 27897
rect 48320 28092 48372 28144
rect 15200 28024 15252 28076
rect 17868 28024 17920 28076
rect 19340 27999 19392 28008
rect 15752 27888 15804 27940
rect 16120 27931 16172 27940
rect 16120 27897 16129 27931
rect 16129 27897 16163 27931
rect 16163 27897 16172 27931
rect 16120 27888 16172 27897
rect 16764 27888 16816 27940
rect 18144 27888 18196 27940
rect 19340 27965 19349 27999
rect 19349 27965 19383 27999
rect 19383 27965 19392 27999
rect 19340 27956 19392 27965
rect 20260 28024 20312 28076
rect 24768 28067 24820 28076
rect 19984 27999 20036 28008
rect 19984 27965 19993 27999
rect 19993 27965 20027 27999
rect 20027 27965 20036 27999
rect 19984 27956 20036 27965
rect 20812 27956 20864 28008
rect 19892 27888 19944 27940
rect 24768 28033 24777 28067
rect 24777 28033 24811 28067
rect 24811 28033 24820 28067
rect 24768 28024 24820 28033
rect 27528 28024 27580 28076
rect 25044 27956 25096 28008
rect 25596 27999 25648 28008
rect 25596 27965 25605 27999
rect 25605 27965 25639 27999
rect 25639 27965 25648 27999
rect 25596 27956 25648 27965
rect 27436 27956 27488 28008
rect 67916 27888 67968 27940
rect 8208 27820 8260 27872
rect 9680 27820 9732 27872
rect 13820 27820 13872 27872
rect 14372 27863 14424 27872
rect 14372 27829 14381 27863
rect 14381 27829 14415 27863
rect 14415 27829 14424 27863
rect 14372 27820 14424 27829
rect 14924 27820 14976 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 13820 27659 13872 27668
rect 13820 27625 13829 27659
rect 13829 27625 13863 27659
rect 13863 27625 13872 27659
rect 13820 27616 13872 27625
rect 14188 27616 14240 27668
rect 16120 27616 16172 27668
rect 17868 27616 17920 27668
rect 7288 27480 7340 27532
rect 9864 27480 9916 27532
rect 8392 27412 8444 27464
rect 10232 27480 10284 27532
rect 12532 27523 12584 27532
rect 12532 27489 12541 27523
rect 12541 27489 12575 27523
rect 12575 27489 12584 27523
rect 12532 27480 12584 27489
rect 13636 27523 13688 27532
rect 13636 27489 13645 27523
rect 13645 27489 13679 27523
rect 13679 27489 13688 27523
rect 13636 27480 13688 27489
rect 13912 27523 13964 27532
rect 13912 27489 13921 27523
rect 13921 27489 13955 27523
rect 13955 27489 13964 27523
rect 13912 27480 13964 27489
rect 14188 27480 14240 27532
rect 14464 27480 14516 27532
rect 8208 27344 8260 27396
rect 9772 27387 9824 27396
rect 9772 27353 9781 27387
rect 9781 27353 9815 27387
rect 9815 27353 9824 27387
rect 9772 27344 9824 27353
rect 10692 27412 10744 27464
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 15292 27455 15344 27464
rect 15292 27421 15301 27455
rect 15301 27421 15335 27455
rect 15335 27421 15344 27455
rect 15292 27412 15344 27421
rect 15752 27412 15804 27464
rect 16304 27412 16356 27464
rect 13728 27344 13780 27396
rect 15660 27344 15712 27396
rect 9588 27276 9640 27328
rect 12624 27276 12676 27328
rect 13912 27276 13964 27328
rect 25044 27548 25096 27600
rect 19340 27412 19392 27464
rect 20812 27480 20864 27532
rect 23388 27480 23440 27532
rect 24952 27523 25004 27532
rect 24952 27489 24961 27523
rect 24961 27489 24995 27523
rect 24995 27489 25004 27523
rect 24952 27480 25004 27489
rect 25320 27523 25372 27532
rect 25320 27489 25329 27523
rect 25329 27489 25363 27523
rect 25363 27489 25372 27523
rect 25320 27480 25372 27489
rect 35440 27548 35492 27600
rect 26700 27523 26752 27532
rect 26700 27489 26709 27523
rect 26709 27489 26743 27523
rect 26743 27489 26752 27523
rect 26700 27480 26752 27489
rect 27436 27523 27488 27532
rect 27436 27489 27445 27523
rect 27445 27489 27479 27523
rect 27479 27489 27488 27523
rect 27436 27480 27488 27489
rect 23480 27412 23532 27464
rect 25872 27412 25924 27464
rect 26240 27412 26292 27464
rect 50160 27344 50212 27396
rect 20168 27319 20220 27328
rect 20168 27285 20177 27319
rect 20177 27285 20211 27319
rect 20211 27285 20220 27319
rect 20168 27276 20220 27285
rect 25872 27319 25924 27328
rect 25872 27285 25881 27319
rect 25881 27285 25915 27319
rect 25915 27285 25924 27319
rect 25872 27276 25924 27285
rect 26240 27319 26292 27328
rect 26240 27285 26249 27319
rect 26249 27285 26283 27319
rect 26283 27285 26292 27319
rect 26240 27276 26292 27285
rect 26792 27276 26844 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 4988 27072 5040 27124
rect 7288 27115 7340 27124
rect 7288 27081 7297 27115
rect 7297 27081 7331 27115
rect 7331 27081 7340 27115
rect 7288 27072 7340 27081
rect 9864 27072 9916 27124
rect 8300 27047 8352 27056
rect 8300 27013 8309 27047
rect 8309 27013 8343 27047
rect 8343 27013 8352 27047
rect 8300 27004 8352 27013
rect 10692 27072 10744 27124
rect 15936 27072 15988 27124
rect 23940 27072 23992 27124
rect 24584 27072 24636 27124
rect 25872 27072 25924 27124
rect 41880 27072 41932 27124
rect 18604 27004 18656 27056
rect 26148 27004 26200 27056
rect 3424 26732 3476 26784
rect 3700 26732 3752 26784
rect 4252 26800 4304 26852
rect 9864 26911 9916 26920
rect 9864 26877 9873 26911
rect 9873 26877 9907 26911
rect 9907 26877 9916 26911
rect 9864 26868 9916 26877
rect 10140 26911 10192 26920
rect 10140 26877 10149 26911
rect 10149 26877 10183 26911
rect 10183 26877 10192 26911
rect 10140 26868 10192 26877
rect 12532 26936 12584 26988
rect 13728 26868 13780 26920
rect 14004 26868 14056 26920
rect 26792 26979 26844 26988
rect 26792 26945 26801 26979
rect 26801 26945 26835 26979
rect 26835 26945 26844 26979
rect 26792 26936 26844 26945
rect 10692 26800 10744 26852
rect 14832 26911 14884 26920
rect 14832 26877 14841 26911
rect 14841 26877 14875 26911
rect 14875 26877 14884 26911
rect 14832 26868 14884 26877
rect 15108 26868 15160 26920
rect 15752 26868 15804 26920
rect 23664 26911 23716 26920
rect 23664 26877 23673 26911
rect 23673 26877 23707 26911
rect 23707 26877 23716 26911
rect 23664 26868 23716 26877
rect 4528 26775 4580 26784
rect 4528 26741 4537 26775
rect 4537 26741 4571 26775
rect 4571 26741 4580 26775
rect 4528 26732 4580 26741
rect 7932 26775 7984 26784
rect 7932 26741 7941 26775
rect 7941 26741 7975 26775
rect 7975 26741 7984 26775
rect 7932 26732 7984 26741
rect 8024 26775 8076 26784
rect 8024 26741 8033 26775
rect 8033 26741 8067 26775
rect 8067 26741 8076 26775
rect 8024 26732 8076 26741
rect 8300 26732 8352 26784
rect 9772 26732 9824 26784
rect 14832 26732 14884 26784
rect 24860 26732 24912 26784
rect 28080 26775 28132 26784
rect 28080 26741 28089 26775
rect 28089 26741 28123 26775
rect 28123 26741 28132 26775
rect 28080 26732 28132 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 5816 26528 5868 26580
rect 6552 26571 6604 26580
rect 6552 26537 6561 26571
rect 6561 26537 6595 26571
rect 6595 26537 6604 26571
rect 6552 26528 6604 26537
rect 8392 26571 8444 26580
rect 8392 26537 8401 26571
rect 8401 26537 8435 26571
rect 8435 26537 8444 26571
rect 8392 26528 8444 26537
rect 10140 26528 10192 26580
rect 4252 26503 4304 26512
rect 4252 26469 4261 26503
rect 4261 26469 4295 26503
rect 4295 26469 4304 26503
rect 4252 26460 4304 26469
rect 4528 26460 4580 26512
rect 10600 26460 10652 26512
rect 15752 26460 15804 26512
rect 5172 26392 5224 26444
rect 5816 26435 5868 26444
rect 5816 26401 5825 26435
rect 5825 26401 5859 26435
rect 5859 26401 5868 26435
rect 5816 26392 5868 26401
rect 8300 26392 8352 26444
rect 10692 26435 10744 26444
rect 10692 26401 10701 26435
rect 10701 26401 10735 26435
rect 10735 26401 10744 26435
rect 10692 26392 10744 26401
rect 19340 26460 19392 26512
rect 22836 26460 22888 26512
rect 23296 26460 23348 26512
rect 27436 26528 27488 26580
rect 28172 26528 28224 26580
rect 17408 26392 17460 26444
rect 22376 26392 22428 26444
rect 23388 26435 23440 26444
rect 23388 26401 23397 26435
rect 23397 26401 23431 26435
rect 23431 26401 23440 26435
rect 23388 26392 23440 26401
rect 63500 26528 63552 26580
rect 24768 26435 24820 26444
rect 24768 26401 24777 26435
rect 24777 26401 24811 26435
rect 24811 26401 24820 26435
rect 24768 26392 24820 26401
rect 28080 26392 28132 26444
rect 4620 26324 4672 26376
rect 4712 26324 4764 26376
rect 5356 26324 5408 26376
rect 17868 26324 17920 26376
rect 18788 26367 18840 26376
rect 18788 26333 18794 26367
rect 18794 26333 18840 26367
rect 18788 26324 18840 26333
rect 19432 26324 19484 26376
rect 22744 26367 22796 26376
rect 22744 26333 22753 26367
rect 22753 26333 22787 26367
rect 22787 26333 22796 26367
rect 22744 26324 22796 26333
rect 28172 26324 28224 26376
rect 4988 26299 5040 26308
rect 4988 26265 4997 26299
rect 4997 26265 5031 26299
rect 5031 26265 5040 26299
rect 4988 26256 5040 26265
rect 11612 26256 11664 26308
rect 57888 26460 57940 26512
rect 5172 26231 5224 26240
rect 5172 26197 5181 26231
rect 5181 26197 5215 26231
rect 5215 26197 5224 26231
rect 5172 26188 5224 26197
rect 8024 26231 8076 26240
rect 8024 26197 8033 26231
rect 8033 26197 8067 26231
rect 8067 26197 8076 26231
rect 8024 26188 8076 26197
rect 8300 26188 8352 26240
rect 17500 26231 17552 26240
rect 17500 26197 17509 26231
rect 17509 26197 17543 26231
rect 17543 26197 17552 26231
rect 17500 26188 17552 26197
rect 56692 26256 56744 26308
rect 55128 26188 55180 26240
rect 56600 26188 56652 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 9864 25984 9916 26036
rect 15936 26027 15988 26036
rect 15936 25993 15945 26027
rect 15945 25993 15979 26027
rect 15979 25993 15988 26027
rect 15936 25984 15988 25993
rect 18420 26027 18472 26036
rect 18420 25993 18429 26027
rect 18429 25993 18463 26027
rect 18463 25993 18472 26027
rect 18420 25984 18472 25993
rect 18788 26027 18840 26036
rect 18788 25993 18797 26027
rect 18797 25993 18831 26027
rect 18831 25993 18840 26027
rect 18788 25984 18840 25993
rect 3884 25916 3936 25968
rect 9956 25916 10008 25968
rect 12716 25916 12768 25968
rect 4804 25848 4856 25900
rect 15936 25780 15988 25832
rect 18604 25823 18656 25832
rect 18604 25789 18613 25823
rect 18613 25789 18647 25823
rect 18647 25789 18656 25823
rect 18604 25780 18656 25789
rect 18972 25780 19024 25832
rect 3792 25644 3844 25696
rect 4436 25687 4488 25696
rect 4436 25653 4445 25687
rect 4445 25653 4479 25687
rect 4479 25653 4488 25687
rect 4436 25644 4488 25653
rect 7932 25687 7984 25696
rect 7932 25653 7941 25687
rect 7941 25653 7975 25687
rect 7975 25653 7984 25687
rect 7932 25644 7984 25653
rect 15844 25644 15896 25696
rect 16212 25687 16264 25696
rect 16212 25653 16221 25687
rect 16221 25653 16255 25687
rect 16255 25653 16264 25687
rect 16212 25644 16264 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 11612 25440 11664 25492
rect 4436 25304 4488 25356
rect 4896 25304 4948 25356
rect 12164 25372 12216 25424
rect 12808 25304 12860 25356
rect 22376 25440 22428 25492
rect 23112 25483 23164 25492
rect 23112 25449 23121 25483
rect 23121 25449 23155 25483
rect 23155 25449 23164 25483
rect 23112 25440 23164 25449
rect 24308 25440 24360 25492
rect 17408 25372 17460 25424
rect 16212 25304 16264 25356
rect 6092 25236 6144 25288
rect 11060 25279 11112 25288
rect 11060 25245 11069 25279
rect 11069 25245 11103 25279
rect 11103 25245 11112 25279
rect 11060 25236 11112 25245
rect 15844 25279 15896 25288
rect 15844 25245 15853 25279
rect 15853 25245 15887 25279
rect 15887 25245 15896 25279
rect 15844 25236 15896 25245
rect 11520 25168 11572 25220
rect 14740 25168 14792 25220
rect 17500 25304 17552 25356
rect 19064 25304 19116 25356
rect 20996 25304 21048 25356
rect 22376 25347 22428 25356
rect 22376 25313 22385 25347
rect 22385 25313 22419 25347
rect 22419 25313 22428 25347
rect 22376 25304 22428 25313
rect 22836 25304 22888 25356
rect 24124 25304 24176 25356
rect 24768 25440 24820 25492
rect 24768 25304 24820 25356
rect 25136 25347 25188 25356
rect 25136 25313 25145 25347
rect 25145 25313 25179 25347
rect 25179 25313 25188 25347
rect 25136 25304 25188 25313
rect 26700 25440 26752 25492
rect 19432 25236 19484 25288
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 24032 25236 24084 25288
rect 24308 25279 24360 25288
rect 24308 25245 24317 25279
rect 24317 25245 24351 25279
rect 24351 25245 24360 25279
rect 24308 25236 24360 25245
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 12164 25100 12216 25152
rect 12716 25143 12768 25152
rect 12716 25109 12725 25143
rect 12725 25109 12759 25143
rect 12759 25109 12768 25143
rect 12716 25100 12768 25109
rect 13544 25100 13596 25152
rect 19340 25100 19392 25152
rect 19616 25143 19668 25152
rect 19616 25109 19625 25143
rect 19625 25109 19659 25143
rect 19659 25109 19668 25143
rect 19616 25100 19668 25109
rect 24676 25100 24728 25152
rect 25412 25143 25464 25152
rect 25412 25109 25421 25143
rect 25421 25109 25455 25143
rect 25455 25109 25464 25143
rect 25412 25100 25464 25109
rect 25964 25168 26016 25220
rect 31760 25168 31812 25220
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 12716 24896 12768 24948
rect 24768 24896 24820 24948
rect 7196 24871 7248 24880
rect 7196 24837 7205 24871
rect 7205 24837 7239 24871
rect 7239 24837 7248 24871
rect 7196 24828 7248 24837
rect 18420 24828 18472 24880
rect 19064 24871 19116 24880
rect 19064 24837 19073 24871
rect 19073 24837 19107 24871
rect 19107 24837 19116 24871
rect 19064 24828 19116 24837
rect 21548 24828 21600 24880
rect 31576 24896 31628 24948
rect 26516 24828 26568 24880
rect 31668 24828 31720 24880
rect 4988 24692 5040 24744
rect 5356 24735 5408 24744
rect 5356 24701 5365 24735
rect 5365 24701 5399 24735
rect 5399 24701 5408 24735
rect 5356 24692 5408 24701
rect 19616 24760 19668 24812
rect 25412 24760 25464 24812
rect 7196 24692 7248 24744
rect 12624 24735 12676 24744
rect 12624 24701 12633 24735
rect 12633 24701 12667 24735
rect 12667 24701 12676 24735
rect 12624 24692 12676 24701
rect 12808 24735 12860 24744
rect 12808 24701 12817 24735
rect 12817 24701 12851 24735
rect 12851 24701 12860 24735
rect 12808 24692 12860 24701
rect 13544 24692 13596 24744
rect 5908 24667 5960 24676
rect 5908 24633 5917 24667
rect 5917 24633 5951 24667
rect 5951 24633 5960 24667
rect 5908 24624 5960 24633
rect 15936 24692 15988 24744
rect 18420 24735 18472 24744
rect 14464 24624 14516 24676
rect 18420 24701 18429 24735
rect 18429 24701 18463 24735
rect 18463 24701 18472 24735
rect 18420 24692 18472 24701
rect 18788 24735 18840 24744
rect 18788 24701 18797 24735
rect 18797 24701 18831 24735
rect 18831 24701 18840 24735
rect 18788 24692 18840 24701
rect 22744 24692 22796 24744
rect 24124 24735 24176 24744
rect 24124 24701 24133 24735
rect 24133 24701 24167 24735
rect 24167 24701 24176 24735
rect 24124 24692 24176 24701
rect 26148 24692 26200 24744
rect 26884 24667 26936 24676
rect 26884 24633 26893 24667
rect 26893 24633 26927 24667
rect 26927 24633 26936 24667
rect 26884 24624 26936 24633
rect 6184 24556 6236 24608
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 18604 24556 18656 24608
rect 23204 24556 23256 24608
rect 24952 24556 25004 24608
rect 25504 24556 25556 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 6092 24352 6144 24404
rect 18420 24352 18472 24404
rect 25136 24352 25188 24404
rect 19432 24284 19484 24336
rect 22468 24284 22520 24336
rect 24676 24327 24728 24336
rect 5632 24216 5684 24268
rect 6920 24216 6972 24268
rect 11520 24259 11572 24268
rect 11520 24225 11529 24259
rect 11529 24225 11563 24259
rect 11563 24225 11572 24259
rect 11520 24216 11572 24225
rect 17500 24216 17552 24268
rect 23204 24259 23256 24268
rect 23204 24225 23213 24259
rect 23213 24225 23247 24259
rect 23247 24225 23256 24259
rect 23204 24216 23256 24225
rect 24676 24293 24685 24327
rect 24685 24293 24719 24327
rect 24719 24293 24728 24327
rect 24676 24284 24728 24293
rect 3332 24148 3384 24200
rect 4068 24148 4120 24200
rect 18052 24148 18104 24200
rect 18788 24148 18840 24200
rect 19432 24148 19484 24200
rect 13544 24080 13596 24132
rect 4804 24055 4856 24064
rect 4804 24021 4813 24055
rect 4813 24021 4847 24055
rect 4847 24021 4856 24055
rect 4804 24012 4856 24021
rect 11152 24055 11204 24064
rect 11152 24021 11161 24055
rect 11161 24021 11195 24055
rect 11195 24021 11204 24055
rect 11152 24012 11204 24021
rect 12716 24012 12768 24064
rect 23940 24259 23992 24268
rect 23940 24225 23949 24259
rect 23949 24225 23983 24259
rect 23983 24225 23992 24259
rect 23940 24216 23992 24225
rect 24584 24216 24636 24268
rect 26884 24216 26936 24268
rect 24124 24080 24176 24132
rect 24584 24012 24636 24064
rect 26884 24055 26936 24064
rect 26884 24021 26893 24055
rect 26893 24021 26927 24055
rect 26927 24021 26936 24055
rect 26884 24012 26936 24021
rect 27436 24012 27488 24064
rect 31576 24012 31628 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 4068 23808 4120 23860
rect 32220 23808 32272 23860
rect 12808 23740 12860 23792
rect 13912 23740 13964 23792
rect 16304 23740 16356 23792
rect 4896 23672 4948 23724
rect 15200 23715 15252 23724
rect 15200 23681 15209 23715
rect 15209 23681 15243 23715
rect 15243 23681 15252 23715
rect 15200 23672 15252 23681
rect 19340 23672 19392 23724
rect 26516 23672 26568 23724
rect 3424 23604 3476 23656
rect 4068 23604 4120 23656
rect 5540 23604 5592 23656
rect 12716 23604 12768 23656
rect 13912 23647 13964 23656
rect 13912 23613 13921 23647
rect 13921 23613 13955 23647
rect 13955 23613 13964 23647
rect 13912 23604 13964 23613
rect 14280 23647 14332 23656
rect 14280 23613 14289 23647
rect 14289 23613 14323 23647
rect 14323 23613 14332 23647
rect 14280 23604 14332 23613
rect 14464 23647 14516 23656
rect 14464 23613 14473 23647
rect 14473 23613 14507 23647
rect 14507 23613 14516 23647
rect 14464 23604 14516 23613
rect 13820 23579 13872 23588
rect 3056 23468 3108 23520
rect 3700 23468 3752 23520
rect 6092 23468 6144 23520
rect 12716 23511 12768 23520
rect 12716 23477 12725 23511
rect 12725 23477 12759 23511
rect 12759 23477 12768 23511
rect 12716 23468 12768 23477
rect 13820 23545 13829 23579
rect 13829 23545 13863 23579
rect 13863 23545 13872 23579
rect 14832 23604 14884 23656
rect 15108 23604 15160 23656
rect 13820 23536 13872 23545
rect 18972 23647 19024 23656
rect 18972 23613 18981 23647
rect 18981 23613 19015 23647
rect 19015 23613 19024 23647
rect 18972 23604 19024 23613
rect 24400 23647 24452 23656
rect 18788 23468 18840 23520
rect 24400 23613 24409 23647
rect 24409 23613 24443 23647
rect 24443 23613 24452 23647
rect 24400 23604 24452 23613
rect 24216 23468 24268 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 4804 23264 4856 23316
rect 5632 23196 5684 23248
rect 5080 23171 5132 23180
rect 5080 23137 5089 23171
rect 5089 23137 5123 23171
rect 5123 23137 5132 23171
rect 5080 23128 5132 23137
rect 6092 23128 6144 23180
rect 5540 23103 5592 23112
rect 3424 22924 3476 22976
rect 5540 23069 5549 23103
rect 5549 23069 5583 23103
rect 5583 23069 5592 23103
rect 5540 23060 5592 23069
rect 12624 23264 12676 23316
rect 13728 23264 13780 23316
rect 22468 23264 22520 23316
rect 24400 23264 24452 23316
rect 24032 23196 24084 23248
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 13728 23128 13780 23180
rect 14280 23128 14332 23180
rect 17500 23128 17552 23180
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 13912 22992 13964 23044
rect 18144 22992 18196 23044
rect 17868 22967 17920 22976
rect 17868 22933 17877 22967
rect 17877 22933 17911 22967
rect 17911 22933 17920 22967
rect 17868 22924 17920 22933
rect 24308 23171 24360 23180
rect 24308 23137 24317 23171
rect 24317 23137 24351 23171
rect 24351 23137 24360 23171
rect 24308 23128 24360 23137
rect 26516 23171 26568 23180
rect 26516 23137 26525 23171
rect 26525 23137 26559 23171
rect 26559 23137 26568 23171
rect 26516 23128 26568 23137
rect 25412 22992 25464 23044
rect 26240 22924 26292 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 8484 22720 8536 22772
rect 9312 22720 9364 22772
rect 13820 22720 13872 22772
rect 17868 22763 17920 22772
rect 17868 22729 17877 22763
rect 17877 22729 17911 22763
rect 17911 22729 17920 22763
rect 17868 22720 17920 22729
rect 5080 22652 5132 22704
rect 8392 22652 8444 22704
rect 13544 22584 13596 22636
rect 4160 22516 4212 22568
rect 8484 22559 8536 22568
rect 8484 22525 8493 22559
rect 8493 22525 8527 22559
rect 8527 22525 8536 22559
rect 8484 22516 8536 22525
rect 13912 22516 13964 22568
rect 14096 22559 14148 22568
rect 14096 22525 14105 22559
rect 14105 22525 14139 22559
rect 14139 22525 14148 22559
rect 14096 22516 14148 22525
rect 14280 22559 14332 22568
rect 14280 22525 14289 22559
rect 14289 22525 14323 22559
rect 14323 22525 14332 22559
rect 14280 22516 14332 22525
rect 14556 22559 14608 22568
rect 14556 22525 14565 22559
rect 14565 22525 14599 22559
rect 14599 22525 14608 22559
rect 14556 22516 14608 22525
rect 15108 22516 15160 22568
rect 17868 22516 17920 22568
rect 18696 22516 18748 22568
rect 18972 22559 19024 22568
rect 18972 22525 18981 22559
rect 18981 22525 19015 22559
rect 19015 22525 19024 22559
rect 18972 22516 19024 22525
rect 19064 22516 19116 22568
rect 23480 22516 23532 22568
rect 23848 22516 23900 22568
rect 3792 22448 3844 22500
rect 8760 22448 8812 22500
rect 24032 22559 24084 22568
rect 24032 22525 24041 22559
rect 24041 22525 24075 22559
rect 24075 22525 24084 22559
rect 24032 22516 24084 22525
rect 25964 22559 26016 22568
rect 24308 22448 24360 22500
rect 25964 22525 25973 22559
rect 25973 22525 26007 22559
rect 26007 22525 26016 22559
rect 25964 22516 26016 22525
rect 3884 22423 3936 22432
rect 3884 22389 3893 22423
rect 3893 22389 3927 22423
rect 3927 22389 3936 22423
rect 3884 22380 3936 22389
rect 8576 22423 8628 22432
rect 8576 22389 8585 22423
rect 8585 22389 8619 22423
rect 8619 22389 8628 22423
rect 8576 22380 8628 22389
rect 18972 22380 19024 22432
rect 24860 22380 24912 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 8024 22219 8076 22228
rect 8024 22185 8033 22219
rect 8033 22185 8067 22219
rect 8067 22185 8076 22219
rect 8024 22176 8076 22185
rect 4160 22083 4212 22092
rect 4160 22049 4169 22083
rect 4169 22049 4203 22083
rect 4203 22049 4212 22083
rect 4160 22040 4212 22049
rect 5080 22040 5132 22092
rect 8576 22040 8628 22092
rect 12164 22083 12216 22092
rect 12164 22049 12173 22083
rect 12173 22049 12207 22083
rect 12207 22049 12216 22083
rect 12164 22040 12216 22049
rect 13176 22108 13228 22160
rect 14096 22040 14148 22092
rect 19064 22176 19116 22228
rect 18604 22040 18656 22092
rect 4620 21836 4672 21888
rect 6552 21836 6604 21888
rect 11060 21904 11112 21956
rect 17868 21972 17920 22024
rect 19156 22083 19208 22092
rect 19156 22049 19165 22083
rect 19165 22049 19199 22083
rect 19199 22049 19208 22083
rect 19156 22040 19208 22049
rect 23664 22176 23716 22228
rect 31576 22176 31628 22228
rect 24124 22083 24176 22092
rect 24124 22049 24133 22083
rect 24133 22049 24167 22083
rect 24167 22049 24176 22083
rect 24124 22040 24176 22049
rect 21180 21972 21232 22024
rect 7472 21836 7524 21888
rect 17960 21904 18012 21956
rect 19156 21904 19208 21956
rect 12716 21836 12768 21888
rect 14096 21836 14148 21888
rect 15108 21836 15160 21888
rect 17868 21836 17920 21888
rect 18236 21836 18288 21888
rect 24216 21836 24268 21888
rect 25412 21879 25464 21888
rect 25412 21845 25421 21879
rect 25421 21845 25455 21879
rect 25455 21845 25464 21879
rect 25412 21836 25464 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 5080 21632 5132 21684
rect 9312 21675 9364 21684
rect 4620 21564 4672 21616
rect 9312 21641 9321 21675
rect 9321 21641 9355 21675
rect 9355 21641 9364 21675
rect 9312 21632 9364 21641
rect 13544 21632 13596 21684
rect 17960 21632 18012 21684
rect 21364 21632 21416 21684
rect 25964 21675 26016 21684
rect 25964 21641 25973 21675
rect 25973 21641 26007 21675
rect 26007 21641 26016 21675
rect 25964 21632 26016 21641
rect 3884 21496 3936 21548
rect 8024 21539 8076 21548
rect 4896 21428 4948 21480
rect 5632 21471 5684 21480
rect 5632 21437 5641 21471
rect 5641 21437 5675 21471
rect 5675 21437 5684 21471
rect 5632 21428 5684 21437
rect 8024 21505 8033 21539
rect 8033 21505 8067 21539
rect 8067 21505 8076 21539
rect 8024 21496 8076 21505
rect 12716 21539 12768 21548
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 24860 21496 24912 21548
rect 11152 21428 11204 21480
rect 21732 21428 21784 21480
rect 14096 21403 14148 21412
rect 14096 21369 14105 21403
rect 14105 21369 14139 21403
rect 14139 21369 14148 21403
rect 14096 21360 14148 21369
rect 4620 21335 4672 21344
rect 4620 21301 4629 21335
rect 4629 21301 4663 21335
rect 4663 21301 4672 21335
rect 4620 21292 4672 21301
rect 10508 21292 10560 21344
rect 15200 21292 15252 21344
rect 15752 21335 15804 21344
rect 15752 21301 15761 21335
rect 15761 21301 15795 21335
rect 15795 21301 15804 21335
rect 15752 21292 15804 21301
rect 24216 21335 24268 21344
rect 24216 21301 24225 21335
rect 24225 21301 24259 21335
rect 24259 21301 24268 21335
rect 24216 21292 24268 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 3792 21088 3844 21140
rect 7472 21088 7524 21140
rect 7564 21088 7616 21140
rect 18236 21088 18288 21140
rect 23664 21063 23716 21072
rect 23664 21029 23673 21063
rect 23673 21029 23707 21063
rect 23707 21029 23716 21063
rect 23664 21020 23716 21029
rect 22284 20927 22336 20936
rect 11060 20816 11112 20868
rect 16212 20816 16264 20868
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 24216 20748 24268 20800
rect 24768 20748 24820 20800
rect 26424 20748 26476 20800
rect 29000 20748 29052 20800
rect 59360 20748 59412 20800
rect 59912 20748 59964 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 3976 20519 4028 20528
rect 3976 20485 3985 20519
rect 3985 20485 4019 20519
rect 4019 20485 4028 20519
rect 3976 20476 4028 20485
rect 5264 20544 5316 20596
rect 15200 20544 15252 20596
rect 16580 20587 16632 20596
rect 14464 20476 14516 20528
rect 15108 20476 15160 20528
rect 16580 20553 16589 20587
rect 16589 20553 16623 20587
rect 16623 20553 16632 20587
rect 16580 20544 16632 20553
rect 23848 20587 23900 20596
rect 23848 20553 23857 20587
rect 23857 20553 23891 20587
rect 23891 20553 23900 20587
rect 23848 20544 23900 20553
rect 2596 20383 2648 20392
rect 2596 20349 2605 20383
rect 2605 20349 2639 20383
rect 2639 20349 2648 20383
rect 2596 20340 2648 20349
rect 5632 20340 5684 20392
rect 14372 20408 14424 20460
rect 15752 20408 15804 20460
rect 15200 20340 15252 20392
rect 15568 20383 15620 20392
rect 15568 20349 15577 20383
rect 15577 20349 15611 20383
rect 15611 20349 15620 20383
rect 15568 20340 15620 20349
rect 17868 20476 17920 20528
rect 17960 20340 18012 20392
rect 27436 20408 27488 20460
rect 23480 20340 23532 20392
rect 23664 20383 23716 20392
rect 23664 20349 23679 20383
rect 23679 20349 23713 20383
rect 23713 20349 23716 20383
rect 23664 20340 23716 20349
rect 26424 20340 26476 20392
rect 4620 20247 4672 20256
rect 4620 20213 4629 20247
rect 4629 20213 4663 20247
rect 4663 20213 4672 20247
rect 4620 20204 4672 20213
rect 6000 20204 6052 20256
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 16580 20272 16632 20324
rect 16764 20272 16816 20324
rect 8392 20204 8444 20256
rect 11428 20204 11480 20256
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 15568 20204 15620 20256
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 18144 20247 18196 20256
rect 18144 20213 18153 20247
rect 18153 20213 18187 20247
rect 18187 20213 18196 20247
rect 18144 20204 18196 20213
rect 22376 20204 22428 20256
rect 23664 20204 23716 20256
rect 27160 20204 27212 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 9128 20000 9180 20052
rect 16120 20000 16172 20052
rect 17960 20043 18012 20052
rect 17960 20009 17969 20043
rect 17969 20009 18003 20043
rect 18003 20009 18012 20043
rect 17960 20000 18012 20009
rect 20444 20043 20496 20052
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 8300 19932 8352 19984
rect 6000 19864 6052 19916
rect 6920 19864 6972 19916
rect 11428 19907 11480 19916
rect 11428 19873 11437 19907
rect 11437 19873 11471 19907
rect 11471 19873 11480 19907
rect 11428 19864 11480 19873
rect 12992 19864 13044 19916
rect 22284 20000 22336 20052
rect 22008 19864 22060 19916
rect 22376 19907 22428 19916
rect 22376 19873 22385 19907
rect 22385 19873 22419 19907
rect 22419 19873 22428 19907
rect 22376 19864 22428 19873
rect 23848 19864 23900 19916
rect 26240 19864 26292 19916
rect 29000 19864 29052 19916
rect 16856 19839 16908 19848
rect 6276 19771 6328 19780
rect 6276 19737 6285 19771
rect 6285 19737 6319 19771
rect 6319 19737 6328 19771
rect 6276 19728 6328 19737
rect 12164 19728 12216 19780
rect 16856 19805 16865 19839
rect 16865 19805 16899 19839
rect 16899 19805 16908 19839
rect 16856 19796 16908 19805
rect 4988 19703 5040 19712
rect 4988 19669 4997 19703
rect 4997 19669 5031 19703
rect 5031 19669 5040 19703
rect 4988 19660 5040 19669
rect 11244 19660 11296 19712
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 20168 19703 20220 19712
rect 12440 19660 12492 19669
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 24952 19660 25004 19712
rect 26608 19703 26660 19712
rect 26608 19669 26617 19703
rect 26617 19669 26651 19703
rect 26651 19669 26660 19703
rect 26608 19660 26660 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 86684 19592 86736 19644
rect 87236 19592 87288 19644
rect 4988 19456 5040 19508
rect 24860 19456 24912 19508
rect 12992 19431 13044 19440
rect 12992 19397 13001 19431
rect 13001 19397 13035 19431
rect 13035 19397 13044 19431
rect 12992 19388 13044 19397
rect 9956 19320 10008 19372
rect 26516 19456 26568 19508
rect 26516 19320 26568 19372
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7840 19116 7892 19168
rect 8300 19295 8352 19304
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 10692 19252 10744 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 24860 19252 24912 19304
rect 27712 19252 27764 19304
rect 17684 19184 17736 19236
rect 25688 19184 25740 19236
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 13728 19116 13780 19168
rect 17040 19159 17092 19168
rect 17040 19125 17049 19159
rect 17049 19125 17083 19159
rect 17083 19125 17092 19159
rect 17040 19116 17092 19125
rect 22008 19116 22060 19168
rect 23572 19116 23624 19168
rect 27252 19116 27304 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 7196 18912 7248 18964
rect 14648 18912 14700 18964
rect 16212 18955 16264 18964
rect 16212 18921 16221 18955
rect 16221 18921 16255 18955
rect 16255 18921 16264 18955
rect 16212 18912 16264 18921
rect 6276 18776 6328 18828
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 16856 18912 16908 18964
rect 12440 18776 12492 18785
rect 4620 18708 4672 18760
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 18972 18844 19024 18896
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 18144 18776 18196 18828
rect 19432 18819 19484 18828
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 23572 18912 23624 18964
rect 23756 18912 23808 18964
rect 25688 18912 25740 18964
rect 27712 18955 27764 18964
rect 22008 18844 22060 18896
rect 24952 18819 25004 18828
rect 18788 18751 18840 18760
rect 10692 18572 10744 18624
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 20260 18708 20312 18760
rect 22836 18708 22888 18760
rect 17224 18640 17276 18692
rect 24952 18785 24961 18819
rect 24961 18785 24995 18819
rect 24995 18785 25004 18819
rect 24952 18776 25004 18785
rect 26608 18776 26660 18828
rect 27712 18921 27721 18955
rect 27721 18921 27755 18955
rect 27755 18921 27764 18955
rect 27712 18912 27764 18921
rect 27160 18819 27212 18828
rect 27160 18785 27169 18819
rect 27169 18785 27203 18819
rect 27203 18785 27212 18819
rect 27160 18776 27212 18785
rect 27252 18819 27304 18828
rect 27252 18785 27261 18819
rect 27261 18785 27295 18819
rect 27295 18785 27304 18819
rect 27252 18776 27304 18785
rect 25136 18640 25188 18692
rect 13728 18615 13780 18624
rect 13728 18581 13737 18615
rect 13737 18581 13771 18615
rect 13771 18581 13780 18615
rect 13728 18572 13780 18581
rect 19156 18572 19208 18624
rect 24952 18572 25004 18624
rect 27252 18572 27304 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 2596 18275 2648 18284
rect 2596 18241 2605 18275
rect 2605 18241 2639 18275
rect 2639 18241 2648 18275
rect 2596 18232 2648 18241
rect 9220 18368 9272 18420
rect 11244 18368 11296 18420
rect 17224 18368 17276 18420
rect 20260 18411 20312 18420
rect 20260 18377 20269 18411
rect 20269 18377 20303 18411
rect 20303 18377 20312 18411
rect 20260 18368 20312 18377
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 9864 18207 9916 18216
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 18788 18164 18840 18216
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 17960 18096 18012 18148
rect 19432 18164 19484 18216
rect 20996 18164 21048 18216
rect 24860 18207 24912 18216
rect 24860 18173 24869 18207
rect 24869 18173 24903 18207
rect 24903 18173 24912 18207
rect 24860 18164 24912 18173
rect 26792 18164 26844 18216
rect 4160 18071 4212 18080
rect 4160 18037 4169 18071
rect 4169 18037 4203 18071
rect 4203 18037 4212 18071
rect 4160 18028 4212 18037
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 13820 18028 13872 18080
rect 24860 18028 24912 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 8024 17756 8076 17808
rect 8208 17756 8260 17808
rect 8116 17620 8168 17672
rect 7748 17484 7800 17536
rect 8116 17484 8168 17536
rect 17960 17688 18012 17740
rect 18236 17688 18288 17740
rect 20168 17824 20220 17876
rect 23940 17824 23992 17876
rect 19340 17756 19392 17808
rect 86684 17756 86736 17808
rect 87604 17756 87656 17808
rect 13360 17620 13412 17672
rect 18604 17663 18656 17672
rect 13084 17552 13136 17604
rect 8576 17484 8628 17536
rect 13544 17484 13596 17536
rect 18236 17484 18288 17536
rect 18604 17629 18613 17663
rect 18613 17629 18647 17663
rect 18647 17629 18656 17663
rect 18604 17620 18656 17629
rect 19432 17552 19484 17604
rect 20260 17484 20312 17536
rect 20812 17484 20864 17536
rect 28080 17688 28132 17740
rect 28908 17688 28960 17740
rect 27344 17484 27396 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 86684 17416 86736 17468
rect 87420 17416 87472 17468
rect 59360 17348 59412 17400
rect 59636 17348 59688 17400
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 9772 17280 9824 17332
rect 9864 17280 9916 17332
rect 10784 17280 10836 17332
rect 13544 17212 13596 17264
rect 17316 17280 17368 17332
rect 13636 17144 13688 17196
rect 7012 17119 7064 17128
rect 3884 17008 3936 17060
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 19432 17187 19484 17196
rect 8576 17008 8628 17060
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 26516 17144 26568 17196
rect 14188 17119 14240 17128
rect 4160 16983 4212 16992
rect 4160 16949 4169 16983
rect 4169 16949 4203 16983
rect 4203 16949 4212 16983
rect 4160 16940 4212 16949
rect 4620 16983 4672 16992
rect 4620 16949 4629 16983
rect 4629 16949 4663 16983
rect 4663 16949 4672 16983
rect 4620 16940 4672 16949
rect 7288 16940 7340 16992
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 15200 17076 15252 17128
rect 20812 17051 20864 17060
rect 20812 17017 20821 17051
rect 20821 17017 20855 17051
rect 20855 17017 20864 17051
rect 20812 17008 20864 17017
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 27344 17119 27396 17128
rect 27344 17085 27353 17119
rect 27353 17085 27387 17119
rect 27387 17085 27396 17119
rect 27344 17076 27396 17085
rect 27252 17008 27304 17060
rect 21640 16940 21692 16992
rect 26792 16940 26844 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 20168 16779 20220 16788
rect 20168 16745 20177 16779
rect 20177 16745 20211 16779
rect 20211 16745 20220 16779
rect 20168 16736 20220 16745
rect 21640 16736 21692 16788
rect 24860 16736 24912 16788
rect 28080 16779 28132 16788
rect 12348 16711 12400 16720
rect 12348 16677 12357 16711
rect 12357 16677 12391 16711
rect 12391 16677 12400 16711
rect 12348 16668 12400 16677
rect 4620 16600 4672 16652
rect 7104 16600 7156 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 13084 16643 13136 16652
rect 12440 16600 12492 16609
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 13268 16600 13320 16652
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 14372 16600 14424 16652
rect 18328 16600 18380 16652
rect 18512 16600 18564 16652
rect 20996 16600 21048 16652
rect 22836 16600 22888 16652
rect 28080 16745 28089 16779
rect 28089 16745 28123 16779
rect 28123 16745 28132 16779
rect 28080 16736 28132 16745
rect 26792 16643 26844 16652
rect 26792 16609 26801 16643
rect 26801 16609 26835 16643
rect 26835 16609 26844 16643
rect 26792 16600 26844 16609
rect 8944 16532 8996 16584
rect 9588 16532 9640 16584
rect 19892 16396 19944 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 8668 16192 8720 16244
rect 8944 16235 8996 16244
rect 8944 16201 8953 16235
rect 8953 16201 8987 16235
rect 8987 16201 8996 16235
rect 8944 16192 8996 16201
rect 7104 16056 7156 16108
rect 12348 16192 12400 16244
rect 2596 16031 2648 16040
rect 2596 15997 2605 16031
rect 2605 15997 2639 16031
rect 2639 15997 2648 16031
rect 2596 15988 2648 15997
rect 4620 15988 4672 16040
rect 7472 16031 7524 16040
rect 7472 15997 7481 16031
rect 7481 15997 7515 16031
rect 7515 15997 7524 16031
rect 7472 15988 7524 15997
rect 21548 16192 21600 16244
rect 23664 16235 23716 16244
rect 23664 16201 23673 16235
rect 23673 16201 23707 16235
rect 23707 16201 23716 16235
rect 23664 16192 23716 16201
rect 24860 16235 24912 16244
rect 24860 16201 24869 16235
rect 24869 16201 24903 16235
rect 24903 16201 24912 16235
rect 24860 16192 24912 16201
rect 26516 16235 26568 16244
rect 26516 16201 26525 16235
rect 26525 16201 26559 16235
rect 26559 16201 26568 16235
rect 26516 16192 26568 16201
rect 28908 16192 28960 16244
rect 19892 16099 19944 16108
rect 19892 16065 19901 16099
rect 19901 16065 19935 16099
rect 19935 16065 19944 16099
rect 19892 16056 19944 16065
rect 4160 15895 4212 15904
rect 4160 15861 4169 15895
rect 4169 15861 4203 15895
rect 4203 15861 4212 15895
rect 4160 15852 4212 15861
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 12624 15852 12676 15904
rect 13912 15852 13964 15904
rect 23664 15988 23716 16040
rect 25228 16031 25280 16040
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 21272 15963 21324 15972
rect 21272 15929 21281 15963
rect 21281 15929 21315 15963
rect 21315 15929 21324 15963
rect 21272 15920 21324 15929
rect 21640 15852 21692 15904
rect 24400 15852 24452 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 7472 15648 7524 15700
rect 20996 15691 21048 15700
rect 20996 15657 21005 15691
rect 21005 15657 21039 15691
rect 21039 15657 21048 15691
rect 20996 15648 21048 15657
rect 21272 15691 21324 15700
rect 21272 15657 21281 15691
rect 21281 15657 21315 15691
rect 21315 15657 21324 15691
rect 21272 15648 21324 15657
rect 25228 15648 25280 15700
rect 7012 15512 7064 15564
rect 9772 15512 9824 15564
rect 24400 15555 24452 15564
rect 24400 15521 24409 15555
rect 24409 15521 24443 15555
rect 24443 15521 24452 15555
rect 24952 15555 25004 15564
rect 24400 15512 24452 15521
rect 24952 15521 24961 15555
rect 24961 15521 24995 15555
rect 24995 15521 25004 15555
rect 24952 15512 25004 15521
rect 26516 15555 26568 15564
rect 26516 15521 26525 15555
rect 26525 15521 26559 15555
rect 26559 15521 26568 15555
rect 26516 15512 26568 15521
rect 6368 15419 6420 15428
rect 6368 15385 6377 15419
rect 6377 15385 6411 15419
rect 6411 15385 6420 15419
rect 18604 15444 18656 15496
rect 6368 15376 6420 15385
rect 18328 15376 18380 15428
rect 25412 15376 25464 15428
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 10416 15104 10468 15156
rect 13912 14968 13964 15020
rect 2596 14900 2648 14952
rect 3976 14900 4028 14952
rect 6368 14900 6420 14952
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 12624 14764 12676 14816
rect 15016 14764 15068 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 21548 14560 21600 14612
rect 14740 14492 14792 14544
rect 18052 14535 18104 14544
rect 18052 14501 18061 14535
rect 18061 14501 18095 14535
rect 18095 14501 18104 14535
rect 18052 14492 18104 14501
rect 12440 14424 12492 14476
rect 20628 14424 20680 14476
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 8392 14288 8444 14340
rect 9036 14288 9088 14340
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 4896 14220 4948 14272
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 20996 14220 21048 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 6184 14016 6236 14068
rect 6828 14016 6880 14068
rect 3700 13948 3752 14000
rect 12624 14016 12676 14068
rect 20628 14016 20680 14068
rect 25412 14059 25464 14068
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 8392 13880 8444 13932
rect 6828 13812 6880 13864
rect 10600 13880 10652 13932
rect 15200 13948 15252 14000
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 12992 13880 13044 13932
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 14740 13812 14792 13864
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 8208 13676 8260 13728
rect 20996 13812 21048 13864
rect 24952 13812 25004 13864
rect 27804 13855 27856 13864
rect 27804 13821 27813 13855
rect 27813 13821 27847 13855
rect 27847 13821 27856 13855
rect 27804 13812 27856 13821
rect 15752 13676 15804 13728
rect 22284 13719 22336 13728
rect 22284 13685 22293 13719
rect 22293 13685 22327 13719
rect 22327 13685 22336 13719
rect 22284 13676 22336 13685
rect 26792 13719 26844 13728
rect 26792 13685 26801 13719
rect 26801 13685 26835 13719
rect 26835 13685 26844 13719
rect 26792 13676 26844 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 6184 13472 6236 13524
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 10508 13515 10560 13524
rect 10508 13481 10517 13515
rect 10517 13481 10551 13515
rect 10551 13481 10560 13515
rect 10508 13472 10560 13481
rect 18052 13472 18104 13524
rect 21640 13472 21692 13524
rect 24308 13472 24360 13524
rect 7288 13404 7340 13456
rect 8484 13336 8536 13388
rect 16672 13404 16724 13456
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 17960 13311 18012 13320
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 9956 13132 10008 13184
rect 15752 13132 15804 13184
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 22284 13336 22336 13388
rect 26792 13379 26844 13388
rect 26792 13345 26801 13379
rect 26801 13345 26835 13379
rect 26835 13345 26844 13379
rect 26792 13336 26844 13345
rect 27620 13132 27672 13184
rect 27804 13132 27856 13184
rect 31760 13132 31812 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 4620 12928 4672 12980
rect 7840 12928 7892 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9772 12928 9824 12980
rect 15200 12928 15252 12980
rect 15752 12971 15804 12980
rect 8208 12903 8260 12912
rect 8208 12869 8217 12903
rect 8217 12869 8251 12903
rect 8251 12869 8260 12903
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 24308 12971 24360 12980
rect 24308 12937 24317 12971
rect 24317 12937 24351 12971
rect 24351 12937 24360 12971
rect 24308 12928 24360 12937
rect 8208 12860 8260 12869
rect 17960 12860 18012 12912
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 4896 12792 4948 12844
rect 9128 12724 9180 12776
rect 14832 12724 14884 12776
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 15752 12724 15804 12776
rect 24860 12724 24912 12776
rect 25044 12724 25096 12776
rect 8392 12699 8444 12708
rect 8392 12665 8401 12699
rect 8401 12665 8435 12699
rect 8435 12665 8444 12699
rect 8392 12656 8444 12665
rect 11152 12699 11204 12708
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 11152 12665 11161 12699
rect 11161 12665 11195 12699
rect 11195 12665 11204 12699
rect 11152 12656 11204 12665
rect 11060 12588 11112 12640
rect 25872 12631 25924 12640
rect 25872 12597 25881 12631
rect 25881 12597 25915 12631
rect 25915 12597 25924 12631
rect 25872 12588 25924 12597
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 10600 12427 10652 12436
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 11060 12384 11112 12436
rect 20260 12384 20312 12436
rect 22836 12427 22888 12436
rect 12532 12316 12584 12368
rect 3332 12248 3384 12300
rect 4988 12248 5040 12300
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 7472 12248 7524 12300
rect 11428 12248 11480 12300
rect 13820 12248 13872 12300
rect 13728 12180 13780 12232
rect 20628 12248 20680 12300
rect 22836 12393 22845 12427
rect 22845 12393 22879 12427
rect 22879 12393 22888 12427
rect 22836 12384 22888 12393
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 20076 12180 20128 12232
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 8392 11840 8444 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 11152 11704 11204 11756
rect 13728 11704 13780 11756
rect 7012 11636 7064 11688
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 17960 11772 18012 11824
rect 19156 11772 19208 11824
rect 17500 11704 17552 11756
rect 20076 11840 20128 11892
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 20996 11747 21048 11756
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 25872 11704 25924 11756
rect 19156 11679 19208 11688
rect 19156 11645 19165 11679
rect 19165 11645 19199 11679
rect 19199 11645 19208 11679
rect 19156 11636 19208 11645
rect 20628 11568 20680 11620
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 4620 11500 4672 11552
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 21640 11543 21692 11552
rect 21640 11509 21649 11543
rect 21649 11509 21683 11543
rect 21683 11509 21692 11543
rect 21640 11500 21692 11509
rect 26424 11500 26476 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 13820 11296 13872 11348
rect 12716 11228 12768 11280
rect 4620 11160 4672 11212
rect 6920 11092 6972 11144
rect 7472 11092 7524 11144
rect 7380 11067 7432 11076
rect 7380 11033 7389 11067
rect 7389 11033 7423 11067
rect 7423 11033 7432 11067
rect 7380 11024 7432 11033
rect 8852 11024 8904 11076
rect 8484 10956 8536 11008
rect 15384 11160 15436 11212
rect 14740 11092 14792 11144
rect 17040 11092 17092 11144
rect 15200 11024 15252 11076
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 18512 11024 18564 11076
rect 14740 10956 14792 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 3976 10752 4028 10804
rect 4620 10684 4672 10736
rect 8392 10752 8444 10804
rect 8852 10752 8904 10804
rect 12624 10752 12676 10804
rect 20628 10752 20680 10804
rect 11244 10684 11296 10736
rect 2596 10659 2648 10668
rect 2596 10625 2605 10659
rect 2605 10625 2639 10659
rect 2639 10625 2648 10659
rect 2596 10616 2648 10625
rect 7840 10616 7892 10668
rect 11428 10616 11480 10668
rect 4620 10548 4672 10600
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 8116 10548 8168 10600
rect 12992 10480 13044 10532
rect 14096 10548 14148 10600
rect 16120 10616 16172 10668
rect 26424 10616 26476 10668
rect 14740 10591 14792 10600
rect 14740 10557 14749 10591
rect 14749 10557 14783 10591
rect 14783 10557 14792 10591
rect 14740 10548 14792 10557
rect 15292 10480 15344 10532
rect 20904 10591 20956 10600
rect 20904 10557 20913 10591
rect 20913 10557 20947 10591
rect 20947 10557 20956 10591
rect 20904 10548 20956 10557
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 26792 10412 26844 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 20904 10208 20956 10260
rect 27620 10208 27672 10260
rect 8392 10072 8444 10124
rect 9864 10072 9916 10124
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 19340 9868 19392 9920
rect 20444 9868 20496 9920
rect 21272 10072 21324 10124
rect 21640 10072 21692 10124
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 22836 10004 22888 10056
rect 25596 9868 25648 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 15292 9707 15344 9716
rect 15292 9673 15301 9707
rect 15301 9673 15335 9707
rect 15335 9673 15344 9707
rect 15292 9664 15344 9673
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 19892 9596 19944 9648
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 8116 9528 8168 9580
rect 13728 9571 13780 9580
rect 13728 9537 13737 9571
rect 13737 9537 13771 9571
rect 13771 9537 13780 9571
rect 13728 9528 13780 9537
rect 17776 9528 17828 9580
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 21272 9571 21324 9580
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 8484 9460 8536 9512
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 17040 9460 17092 9512
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 18052 9435 18104 9444
rect 18052 9401 18061 9435
rect 18061 9401 18095 9435
rect 18095 9401 18104 9435
rect 18052 9392 18104 9401
rect 19064 9503 19116 9512
rect 19064 9469 19073 9503
rect 19073 9469 19107 9503
rect 19107 9469 19116 9503
rect 19064 9460 19116 9469
rect 3516 9324 3568 9376
rect 7748 9324 7800 9376
rect 22192 9324 22244 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 7840 9120 7892 9172
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 7380 9052 7432 9104
rect 19432 9095 19484 9104
rect 19432 9061 19441 9095
rect 19441 9061 19475 9095
rect 19475 9061 19484 9095
rect 19432 9052 19484 9061
rect 17776 9027 17828 9036
rect 4988 8984 5040 8993
rect 17776 8993 17785 9027
rect 17785 8993 17819 9027
rect 17819 8993 17828 9027
rect 17776 8984 17828 8993
rect 18052 9027 18104 9036
rect 18052 8993 18061 9027
rect 18061 8993 18095 9027
rect 18095 8993 18104 9027
rect 18052 8984 18104 8993
rect 5632 8916 5684 8968
rect 19340 8916 19392 8968
rect 22192 8959 22244 8968
rect 22192 8925 22201 8959
rect 22201 8925 22235 8959
rect 22235 8925 22244 8959
rect 22192 8916 22244 8925
rect 22284 8780 22336 8832
rect 23940 8780 23992 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 4988 8576 5040 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 14004 8576 14056 8628
rect 19064 8576 19116 8628
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 7104 8440 7156 8492
rect 7380 8440 7432 8492
rect 9772 8440 9824 8492
rect 11060 8440 11112 8492
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 12624 8372 12676 8424
rect 22192 8372 22244 8424
rect 22284 8372 22336 8424
rect 25596 8372 25648 8424
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 7380 8032 7432 8084
rect 4068 7896 4120 7905
rect 11060 7896 11112 7948
rect 8116 7828 8168 7880
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 4068 7488 4120 7540
rect 8760 7488 8812 7540
rect 9772 7488 9824 7540
rect 15200 7531 15252 7540
rect 15200 7497 15209 7531
rect 15209 7497 15243 7531
rect 15243 7497 15252 7531
rect 15200 7488 15252 7497
rect 3700 7352 3752 7404
rect 7380 7352 7432 7404
rect 8760 7284 8812 7336
rect 13912 7327 13964 7336
rect 9772 7216 9824 7268
rect 12072 7216 12124 7268
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 12532 7148 12584 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 13912 6919 13964 6928
rect 13912 6885 13921 6919
rect 13921 6885 13955 6919
rect 13955 6885 13964 6919
rect 13912 6876 13964 6885
rect 8116 6808 8168 6860
rect 8760 6808 8812 6860
rect 12072 6851 12124 6860
rect 12072 6817 12081 6851
rect 12081 6817 12115 6851
rect 12115 6817 12124 6851
rect 12072 6808 12124 6817
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 3976 6740 4028 6792
rect 6552 6740 6604 6792
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 3884 6400 3936 6452
rect 8576 6264 8628 6316
rect 4160 6060 4212 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 2964 5312 3016 5364
rect 4804 5312 4856 5364
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 25596 5244 25648 5296
rect 29920 5040 29972 5092
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 12072 4768 12124 4820
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 5908 4088 5960 4140
rect 3976 4020 4028 4072
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 4068 3680 4120 3732
rect 11060 3680 11112 3732
rect 3332 3612 3384 3664
rect 7932 3612 7984 3664
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 4712 3179 4764 3188
rect 4712 3145 4721 3179
rect 4721 3145 4755 3179
rect 4755 3145 4764 3179
rect 4712 3136 4764 3145
rect 3976 2932 4028 2984
rect 2780 2796 2832 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 2872 2252 2924 2304
rect 4988 2252 5040 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 3240 1708 3292 1760
rect 8024 1708 8076 1760
rect 3424 688 3476 740
rect 8208 688 8260 740
<< metal2 >>
rect 3974 49736 4030 49745
rect 3974 49671 4030 49680
rect 2778 49056 2834 49065
rect 2778 48991 2834 49000
rect 2792 46714 2820 48991
rect 3988 48346 4016 49671
rect 18142 49248 18198 50048
rect 54482 49248 54538 50048
rect 90822 49248 90878 50048
rect 4068 48408 4120 48414
rect 4066 48376 4068 48385
rect 14924 48408 14976 48414
rect 4120 48376 4122 48385
rect 3976 48340 4028 48346
rect 14924 48350 14976 48356
rect 4066 48311 4122 48320
rect 3976 48282 4028 48288
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 8392 47660 8444 47666
rect 8392 47602 8444 47608
rect 7932 47592 7984 47598
rect 7932 47534 7984 47540
rect 7944 47122 7972 47534
rect 3424 47116 3476 47122
rect 3424 47058 3476 47064
rect 7932 47116 7984 47122
rect 7932 47058 7984 47064
rect 2780 46708 2832 46714
rect 2780 46650 2832 46656
rect 2792 46578 2820 46650
rect 2780 46572 2832 46578
rect 2780 46514 2832 46520
rect 2596 46504 2648 46510
rect 2596 46446 2648 46452
rect 2608 45422 2636 46446
rect 2596 45416 2648 45422
rect 2596 45358 2648 45364
rect 2608 44334 2636 45358
rect 2596 44328 2648 44334
rect 2596 44270 2648 44276
rect 2608 43246 2636 44270
rect 2596 43240 2648 43246
rect 2596 43182 2648 43188
rect 2596 42220 2648 42226
rect 2596 42162 2648 42168
rect 2608 41070 2636 42162
rect 2596 41064 2648 41070
rect 2596 41006 2648 41012
rect 2608 35698 2636 41006
rect 2596 35692 2648 35698
rect 2596 35634 2648 35640
rect 2792 34202 2820 46514
rect 2964 45280 3016 45286
rect 2964 45222 3016 45228
rect 2872 44192 2924 44198
rect 2872 44134 2924 44140
rect 2884 39953 2912 44134
rect 2870 39944 2926 39953
rect 2870 39879 2926 39888
rect 2976 37369 3004 45222
rect 3056 40520 3108 40526
rect 3056 40462 3108 40468
rect 2962 37360 3018 37369
rect 2962 37295 3018 37304
rect 3068 35698 3096 40462
rect 3436 38593 3464 47058
rect 4712 46912 4764 46918
rect 4712 46854 4764 46860
rect 7196 46912 7248 46918
rect 7196 46854 7248 46860
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4724 46374 4752 46854
rect 7208 46510 7236 46854
rect 7196 46504 7248 46510
rect 7196 46446 7248 46452
rect 7944 46458 7972 47058
rect 8404 46578 8432 47602
rect 13728 47592 13780 47598
rect 13728 47534 13780 47540
rect 12072 47456 12124 47462
rect 12072 47398 12124 47404
rect 12084 46986 12112 47398
rect 12072 46980 12124 46986
rect 12072 46922 12124 46928
rect 13360 46980 13412 46986
rect 13360 46922 13412 46928
rect 8392 46572 8444 46578
rect 8392 46514 8444 46520
rect 4160 46368 4212 46374
rect 4160 46310 4212 46316
rect 4712 46368 4764 46374
rect 4712 46310 4764 46316
rect 4172 45914 4200 46310
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4080 45886 4200 45914
rect 4080 45121 4108 45886
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4632 45490 4660 46106
rect 4620 45484 4672 45490
rect 4620 45426 4672 45432
rect 4436 45280 4488 45286
rect 4436 45222 4488 45228
rect 4066 45112 4122 45121
rect 4448 45082 4476 45222
rect 4724 45082 4752 46310
rect 7104 46028 7156 46034
rect 7104 45970 7156 45976
rect 4066 45047 4122 45056
rect 4436 45076 4488 45082
rect 4436 45018 4488 45024
rect 4712 45076 4764 45082
rect 4712 45018 4764 45024
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4724 44538 4752 45018
rect 6920 44872 6972 44878
rect 6920 44814 6972 44820
rect 4712 44532 4764 44538
rect 4712 44474 4764 44480
rect 4620 44192 4672 44198
rect 4620 44134 4672 44140
rect 3974 43888 4030 43897
rect 3974 43823 4030 43832
rect 3700 43716 3752 43722
rect 3700 43658 3752 43664
rect 3608 40996 3660 41002
rect 3608 40938 3660 40944
rect 3516 38752 3568 38758
rect 3516 38694 3568 38700
rect 3422 38584 3478 38593
rect 3422 38519 3478 38528
rect 3424 37800 3476 37806
rect 3528 37788 3556 38694
rect 3476 37760 3556 37788
rect 3424 37742 3476 37748
rect 3332 36576 3384 36582
rect 3332 36518 3384 36524
rect 3240 36304 3292 36310
rect 3240 36246 3292 36252
rect 3056 35692 3108 35698
rect 3056 35634 3108 35640
rect 3148 35488 3200 35494
rect 3068 35436 3148 35442
rect 3068 35430 3200 35436
rect 3068 35414 3188 35430
rect 2780 34196 2832 34202
rect 2780 34138 2832 34144
rect 2964 32360 3016 32366
rect 2964 32302 3016 32308
rect 2872 32224 2924 32230
rect 2872 32166 2924 32172
rect 2780 29572 2832 29578
rect 2780 29514 2832 29520
rect 2596 29164 2648 29170
rect 2596 29106 2648 29112
rect 2608 28082 2636 29106
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2792 24993 2820 29514
rect 2884 28257 2912 32166
rect 2976 31278 3004 32302
rect 2964 31272 3016 31278
rect 2964 31214 3016 31220
rect 2976 30258 3004 31214
rect 2964 30252 3016 30258
rect 2964 30194 3016 30200
rect 3068 29170 3096 35414
rect 3148 35284 3200 35290
rect 3148 35226 3200 35232
rect 3160 32434 3188 35226
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 3148 30048 3200 30054
rect 3148 29990 3200 29996
rect 3056 29164 3108 29170
rect 3056 29106 3108 29112
rect 3054 29064 3110 29073
rect 3054 28999 3110 29008
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2870 28248 2926 28257
rect 2870 28183 2926 28192
rect 2976 27962 3004 28494
rect 2884 27934 3004 27962
rect 2778 24984 2834 24993
rect 2778 24919 2834 24928
rect 2884 22409 2912 27934
rect 2964 27872 3016 27878
rect 2964 27814 3016 27820
rect 2976 24313 3004 27814
rect 2962 24304 3018 24313
rect 2962 24239 3018 24248
rect 3068 23526 3096 28999
rect 3056 23520 3108 23526
rect 3056 23462 3108 23468
rect 2870 22400 2926 22409
rect 2870 22335 2926 22344
rect 3160 21729 3188 29990
rect 3252 29578 3280 36246
rect 3240 29572 3292 29578
rect 3240 29514 3292 29520
rect 3344 29458 3372 36518
rect 3252 29430 3372 29458
rect 3252 26353 3280 29430
rect 3436 29322 3464 37742
rect 3516 35216 3568 35222
rect 3516 35158 3568 35164
rect 3528 31226 3556 35158
rect 3620 33522 3648 40938
rect 3712 34105 3740 43658
rect 3988 43450 4016 43823
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 3976 43444 4028 43450
rect 3976 43386 4028 43392
rect 4066 43208 4122 43217
rect 4066 43143 4122 43152
rect 4080 42906 4108 43143
rect 4068 42900 4120 42906
rect 4068 42842 4120 42848
rect 4068 42628 4120 42634
rect 4068 42570 4120 42576
rect 3974 42528 4030 42537
rect 3974 42463 4030 42472
rect 3988 42362 4016 42463
rect 3976 42356 4028 42362
rect 3976 42298 4028 42304
rect 4080 41857 4108 42570
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4632 42362 4660 44134
rect 4724 43382 4752 44474
rect 6736 44328 6788 44334
rect 6736 44270 6788 44276
rect 4712 43376 4764 43382
rect 4712 43318 4764 43324
rect 4724 43110 4752 43318
rect 4712 43104 4764 43110
rect 4764 43052 4936 43058
rect 4712 43046 4936 43052
rect 4724 43030 4936 43046
rect 4620 42356 4672 42362
rect 4672 42316 4752 42344
rect 4620 42298 4672 42304
rect 4066 41848 4122 41857
rect 4066 41783 4122 41792
rect 4620 41812 4672 41818
rect 4620 41754 4672 41760
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4066 41304 4122 41313
rect 4220 41296 4516 41316
rect 4066 41239 4068 41248
rect 4120 41239 4122 41248
rect 4068 41210 4120 41216
rect 3976 41132 4028 41138
rect 3976 41074 4028 41080
rect 3884 40180 3936 40186
rect 3884 40122 3936 40128
rect 3792 39636 3844 39642
rect 3792 39578 3844 39584
rect 3804 39273 3832 39578
rect 3790 39264 3846 39273
rect 3790 39199 3846 39208
rect 3792 37664 3844 37670
rect 3792 37606 3844 37612
rect 3804 36718 3832 37606
rect 3792 36712 3844 36718
rect 3896 36689 3924 40122
rect 3792 36654 3844 36660
rect 3882 36680 3938 36689
rect 3882 36615 3938 36624
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 3698 34096 3754 34105
rect 3698 34031 3754 34040
rect 3608 33516 3660 33522
rect 3608 33458 3660 33464
rect 3804 33266 3832 34886
rect 3988 34785 4016 41074
rect 4632 41070 4660 41754
rect 4724 41206 4752 42316
rect 4804 42152 4856 42158
rect 4804 42094 4856 42100
rect 4712 41200 4764 41206
rect 4712 41142 4764 41148
rect 4620 41064 4672 41070
rect 4620 41006 4672 41012
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4816 40118 4844 42094
rect 4804 40112 4856 40118
rect 4804 40054 4856 40060
rect 4804 39976 4856 39982
rect 4908 39930 4936 43030
rect 6748 42838 6776 44270
rect 6932 43994 6960 44814
rect 7012 44736 7064 44742
rect 7012 44678 7064 44684
rect 6920 43988 6972 43994
rect 6920 43930 6972 43936
rect 6736 42832 6788 42838
rect 6736 42774 6788 42780
rect 6828 41608 6880 41614
rect 6828 41550 6880 41556
rect 6840 41070 6868 41550
rect 7024 41274 7052 44678
rect 7116 43858 7144 45970
rect 7208 45082 7236 46446
rect 7944 46430 8064 46458
rect 7932 46368 7984 46374
rect 7932 46310 7984 46316
rect 7196 45076 7248 45082
rect 7196 45018 7248 45024
rect 7840 44532 7892 44538
rect 7840 44474 7892 44480
rect 7852 43994 7880 44474
rect 7840 43988 7892 43994
rect 7840 43930 7892 43936
rect 7104 43852 7156 43858
rect 7104 43794 7156 43800
rect 7116 42770 7144 43794
rect 7564 43104 7616 43110
rect 7564 43046 7616 43052
rect 7104 42764 7156 42770
rect 7104 42706 7156 42712
rect 7116 42362 7144 42706
rect 7104 42356 7156 42362
rect 7104 42298 7156 42304
rect 7288 42152 7340 42158
rect 7288 42094 7340 42100
rect 7300 41682 7328 42094
rect 7288 41676 7340 41682
rect 7288 41618 7340 41624
rect 7012 41268 7064 41274
rect 7012 41210 7064 41216
rect 5540 41064 5592 41070
rect 5540 41006 5592 41012
rect 6828 41064 6880 41070
rect 6828 41006 6880 41012
rect 5552 40662 5580 41006
rect 5540 40656 5592 40662
rect 5540 40598 5592 40604
rect 6840 40594 6868 41006
rect 7012 40928 7064 40934
rect 7012 40870 7064 40876
rect 6828 40588 6880 40594
rect 6828 40530 6880 40536
rect 4988 40112 5040 40118
rect 4988 40054 5040 40060
rect 4856 39924 4936 39930
rect 4804 39918 4936 39924
rect 4816 39902 4936 39918
rect 4620 39500 4672 39506
rect 4620 39442 4672 39448
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4632 39098 4660 39442
rect 4712 39296 4764 39302
rect 4712 39238 4764 39244
rect 4620 39092 4672 39098
rect 4620 39034 4672 39040
rect 4620 38888 4672 38894
rect 4620 38830 4672 38836
rect 4068 38548 4120 38554
rect 4068 38490 4120 38496
rect 4080 38049 4108 38490
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4066 38040 4122 38049
rect 4220 38032 4516 38052
rect 4632 38010 4660 38830
rect 4724 38010 4752 39238
rect 4816 39098 4844 39902
rect 4804 39092 4856 39098
rect 4804 39034 4856 39040
rect 4816 38962 4844 39034
rect 4804 38956 4856 38962
rect 4804 38898 4856 38904
rect 4066 37975 4122 37984
rect 4620 38004 4672 38010
rect 4620 37946 4672 37952
rect 4712 38004 4764 38010
rect 4712 37946 4764 37952
rect 4816 37466 4844 38898
rect 4804 37460 4856 37466
rect 4804 37402 4856 37408
rect 4804 37256 4856 37262
rect 4804 37198 4856 37204
rect 4068 37120 4120 37126
rect 4068 37062 4120 37068
rect 4080 36009 4108 37062
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4816 36854 4844 37198
rect 4804 36848 4856 36854
rect 4804 36790 4856 36796
rect 4804 36372 4856 36378
rect 4804 36314 4856 36320
rect 4066 36000 4122 36009
rect 4066 35935 4122 35944
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4068 35828 4120 35834
rect 4068 35770 4120 35776
rect 4080 35465 4108 35770
rect 4712 35624 4764 35630
rect 4712 35566 4764 35572
rect 4160 35488 4212 35494
rect 4066 35456 4122 35465
rect 4160 35430 4212 35436
rect 4066 35391 4122 35400
rect 4172 35034 4200 35430
rect 4080 35006 4200 35034
rect 3974 34776 4030 34785
rect 3974 34711 4030 34720
rect 3976 33516 4028 33522
rect 3976 33458 4028 33464
rect 3712 33238 3832 33266
rect 3528 31198 3648 31226
rect 3516 31136 3568 31142
rect 3516 31078 3568 31084
rect 3528 30841 3556 31078
rect 3514 30832 3570 30841
rect 3514 30767 3570 30776
rect 3620 30716 3648 31198
rect 3344 29294 3464 29322
rect 3528 30688 3648 30716
rect 3344 27577 3372 29294
rect 3424 29164 3476 29170
rect 3424 29106 3476 29112
rect 3330 27568 3386 27577
rect 3330 27503 3386 27512
rect 3436 26897 3464 29106
rect 3528 28082 3556 30688
rect 3608 30388 3660 30394
rect 3608 30330 3660 30336
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 3422 26888 3478 26897
rect 3620 26874 3648 30330
rect 3422 26823 3478 26832
rect 3528 26846 3648 26874
rect 3424 26784 3476 26790
rect 3424 26726 3476 26732
rect 3238 26344 3294 26353
rect 3238 26279 3294 26288
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3146 21720 3202 21729
rect 3146 21655 3202 21664
rect 2596 20392 2648 20398
rect 2596 20334 2648 20340
rect 2608 18290 2636 20334
rect 3344 19145 3372 24142
rect 3436 23662 3464 26726
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3330 19136 3386 19145
rect 3330 19071 3386 19080
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 2608 17202 2636 18226
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16046 2636 17138
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2608 13938 2636 14894
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2608 12850 2636 13874
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2608 11762 2636 12786
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3344 12073 3372 12242
rect 3330 12064 3386 12073
rect 3330 11999 3386 12008
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2608 10674 2636 11698
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2608 8498 2636 10610
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 3436 5545 3464 22918
rect 3528 17241 3556 26846
rect 3712 26790 3740 33238
rect 3792 33108 3844 33114
rect 3792 33050 3844 33056
rect 3804 32745 3832 33050
rect 3790 32736 3846 32745
rect 3790 32671 3846 32680
rect 3792 32564 3844 32570
rect 3792 32506 3844 32512
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3804 26602 3832 32506
rect 3884 30320 3936 30326
rect 3884 30262 3936 30268
rect 3896 30161 3924 30262
rect 3882 30152 3938 30161
rect 3882 30087 3938 30096
rect 3988 30036 4016 33458
rect 4080 33425 4108 35006
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4528 34060 4580 34066
rect 4528 34002 4580 34008
rect 4540 33946 4568 34002
rect 4540 33918 4660 33946
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4066 33416 4122 33425
rect 4066 33351 4122 33360
rect 4160 33312 4212 33318
rect 4160 33254 4212 33260
rect 4172 32858 4200 33254
rect 4080 32830 4200 32858
rect 4080 32201 4108 32830
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4066 32192 4122 32201
rect 4066 32127 4122 32136
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4066 31512 4122 31521
rect 4220 31504 4516 31524
rect 4066 31447 4122 31456
rect 4080 31414 4108 31447
rect 4068 31408 4120 31414
rect 4068 31350 4120 31356
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 3896 30008 4016 30036
rect 3896 26874 3924 30008
rect 4080 29617 4108 30534
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4436 30048 4488 30054
rect 4436 29990 4488 29996
rect 4448 29850 4476 29990
rect 4436 29844 4488 29850
rect 4436 29786 4488 29792
rect 4066 29608 4122 29617
rect 4066 29543 4122 29552
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 3974 28928 4030 28937
rect 3974 28863 4030 28872
rect 3988 28694 4016 28863
rect 3976 28688 4028 28694
rect 3976 28630 4028 28636
rect 3896 26846 4016 26874
rect 3620 26574 3832 26602
rect 3514 17232 3570 17241
rect 3514 17167 3570 17176
rect 3620 15881 3648 26574
rect 3884 25968 3936 25974
rect 3884 25910 3936 25916
rect 3792 25696 3844 25702
rect 3896 25673 3924 25910
rect 3792 25638 3844 25644
rect 3882 25664 3938 25673
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 3712 18465 3740 23462
rect 3804 23089 3832 25638
rect 3882 25599 3938 25608
rect 3790 23080 3846 23089
rect 3790 23015 3846 23024
rect 3792 22500 3844 22506
rect 3792 22442 3844 22448
rect 3804 21146 3832 22442
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3896 21554 3924 22374
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3698 18456 3754 18465
rect 3698 18391 3754 18400
rect 3606 15872 3662 15881
rect 3606 15807 3662 15816
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3516 9376 3568 9382
rect 3514 9344 3516 9353
rect 3568 9344 3570 9353
rect 3514 9279 3570 9288
rect 3712 7410 3740 13942
rect 3804 8129 3832 21082
rect 3988 20618 4016 26846
rect 4080 24206 4108 29446
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4632 28762 4660 33918
rect 4724 33658 4752 35566
rect 4712 33652 4764 33658
rect 4712 33594 4764 33600
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4724 31278 4752 32166
rect 4712 31272 4764 31278
rect 4712 31214 4764 31220
rect 4724 31142 4752 31214
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4724 30734 4752 31078
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4724 30258 4752 30670
rect 4712 30252 4764 30258
rect 4712 30194 4764 30200
rect 4724 29714 4752 30194
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 4724 29306 4752 29650
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4632 28626 4660 28698
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4252 26852 4304 26858
rect 4252 26794 4304 26800
rect 4264 26518 4292 26794
rect 4528 26784 4580 26790
rect 4528 26726 4580 26732
rect 4540 26518 4568 26726
rect 4252 26512 4304 26518
rect 4252 26454 4304 26460
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4632 26382 4660 28358
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4436 25696 4488 25702
rect 4436 25638 4488 25644
rect 4448 25362 4476 25638
rect 4436 25356 4488 25362
rect 4436 25298 4488 25304
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4080 23769 4108 23802
rect 4066 23760 4122 23769
rect 4066 23695 4122 23704
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 4080 21049 4108 23598
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4172 22098 4200 22510
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4632 21622 4660 21830
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4066 21040 4122 21049
rect 4066 20975 4122 20984
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 3896 20590 4016 20618
rect 3896 19825 3924 20590
rect 3976 20528 4028 20534
rect 3974 20496 3976 20505
rect 4028 20496 4030 20505
rect 3974 20431 4030 20440
rect 4632 20262 4660 21286
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 3882 19816 3938 19825
rect 3882 19751 3938 19760
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4632 18766 4660 20198
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4632 18086 4660 18702
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4066 17912 4122 17921
rect 4172 17898 4200 18022
rect 4122 17870 4200 17898
rect 4066 17847 4122 17856
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 3896 13297 3924 17002
rect 4632 16998 4660 18022
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4066 16552 4122 16561
rect 4172 16538 4200 16934
rect 4632 16658 4660 16934
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4122 16510 4200 16538
rect 4066 16487 4122 16496
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4632 16046 4660 16594
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15450 4200 15846
rect 4080 15422 4200 15450
rect 4080 15201 4108 15422
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4066 15192 4122 15201
rect 4220 15184 4516 15204
rect 4066 15127 4122 15136
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14657 4016 14894
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 3974 14648 4030 14657
rect 3974 14583 4030 14592
rect 4080 13977 4108 14758
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4632 14074 4660 14758
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4066 13968 4122 13977
rect 4066 13903 4122 13912
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3882 13288 3938 13297
rect 3882 13223 3938 13232
rect 3988 12617 4016 13670
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4632 12986 4660 14010
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4160 12640 4212 12646
rect 3974 12608 4030 12617
rect 4160 12582 4212 12588
rect 3974 12543 4030 12552
rect 4172 12186 4200 12582
rect 3988 12158 4200 12186
rect 3988 11393 4016 12158
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4632 11558 4660 12922
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 4172 11098 4200 11494
rect 4632 11218 4660 11494
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4080 11070 4200 11098
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3988 10713 4016 10746
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 4080 10146 4108 11070
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4632 10742 4660 11154
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4632 10606 4660 10678
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 3988 10118 4108 10146
rect 3988 10033 4016 10118
rect 3974 10024 4030 10033
rect 4172 10010 4200 10406
rect 3974 9959 4030 9968
rect 4080 9982 4200 10010
rect 4080 8809 4108 9982
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3790 8120 3846 8129
rect 3790 8055 3846 8064
rect 3988 7449 4016 8230
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4080 7546 4108 7890
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3974 7440 4030 7449
rect 3700 7404 3752 7410
rect 3974 7375 4030 7384
rect 3700 7346 3752 7352
rect 4080 6882 4108 7482
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3896 6854 4108 6882
rect 3896 6458 3924 6854
rect 3976 6792 4028 6798
rect 3974 6760 3976 6769
rect 4028 6760 4030 6769
rect 4172 6746 4200 7142
rect 3974 6695 4030 6704
rect 4080 6718 4200 6746
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2976 4185 3004 5306
rect 2962 4176 3018 4185
rect 3896 4162 3924 6394
rect 4080 6225 4108 6718
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5658 4200 6054
rect 4080 5630 4200 5658
rect 4080 4865 4108 5630
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3896 4134 4016 4162
rect 2962 4111 3018 4120
rect 3988 4078 4016 4134
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3344 2961 3372 3606
rect 3988 2990 4016 4014
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4080 3505 4108 3674
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4724 3194 4752 26318
rect 4816 25906 4844 36314
rect 4896 35692 4948 35698
rect 4896 35634 4948 35640
rect 4908 35154 4936 35634
rect 4896 35148 4948 35154
rect 4896 35090 4948 35096
rect 4908 34542 4936 35090
rect 4896 34536 4948 34542
rect 4896 34478 4948 34484
rect 4908 34202 4936 34478
rect 4896 34196 4948 34202
rect 4896 34138 4948 34144
rect 4896 33992 4948 33998
rect 4896 33934 4948 33940
rect 4908 30394 4936 33934
rect 5000 33862 5028 40054
rect 5080 38208 5132 38214
rect 5080 38150 5132 38156
rect 5092 38010 5120 38150
rect 5080 38004 5132 38010
rect 5080 37946 5132 37952
rect 5092 37806 5120 37946
rect 5080 37800 5132 37806
rect 5080 37742 5132 37748
rect 5632 37800 5684 37806
rect 5632 37742 5684 37748
rect 5092 36582 5120 37742
rect 5644 37466 5672 37742
rect 5724 37732 5776 37738
rect 5724 37674 5776 37680
rect 5632 37460 5684 37466
rect 5632 37402 5684 37408
rect 5736 37330 5764 37674
rect 6000 37392 6052 37398
rect 6000 37334 6052 37340
rect 5724 37324 5776 37330
rect 5724 37266 5776 37272
rect 5736 36922 5764 37266
rect 5724 36916 5776 36922
rect 5724 36858 5776 36864
rect 5540 36848 5592 36854
rect 5540 36790 5592 36796
rect 5080 36576 5132 36582
rect 5080 36518 5132 36524
rect 5264 36236 5316 36242
rect 5264 36178 5316 36184
rect 5276 35698 5304 36178
rect 5264 35692 5316 35698
rect 5264 35634 5316 35640
rect 5552 35290 5580 36790
rect 6012 35766 6040 37334
rect 6920 36644 6972 36650
rect 6920 36586 6972 36592
rect 6000 35760 6052 35766
rect 6000 35702 6052 35708
rect 5540 35284 5592 35290
rect 5540 35226 5592 35232
rect 5552 35154 5580 35226
rect 6932 35154 6960 36586
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 6092 35148 6144 35154
rect 6092 35090 6144 35096
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 5080 35012 5132 35018
rect 5080 34954 5132 34960
rect 4988 33856 5040 33862
rect 4988 33798 5040 33804
rect 4896 30388 4948 30394
rect 4896 30330 4948 30336
rect 4896 29300 4948 29306
rect 4896 29242 4948 29248
rect 4908 27878 4936 29242
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4908 25362 4936 27814
rect 5000 27130 5028 33798
rect 5092 28558 5120 34954
rect 5264 34468 5316 34474
rect 5264 34410 5316 34416
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 4988 26308 5040 26314
rect 4988 26250 5040 26256
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 5000 24750 5028 26250
rect 5184 26246 5212 26386
rect 5172 26240 5224 26246
rect 5170 26208 5172 26217
rect 5224 26208 5226 26217
rect 5170 26143 5226 26152
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4816 23322 4844 24006
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4816 5370 4844 23258
rect 4908 21486 4936 23666
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5092 22710 5120 23122
rect 5080 22704 5132 22710
rect 5080 22646 5132 22652
rect 5092 22098 5120 22646
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 5092 21690 5120 22034
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 5276 20602 5304 34410
rect 6104 34202 6132 35090
rect 6368 34400 6420 34406
rect 6368 34342 6420 34348
rect 6092 34196 6144 34202
rect 6092 34138 6144 34144
rect 6380 29073 6408 34342
rect 6552 32496 6604 32502
rect 6552 32438 6604 32444
rect 6366 29064 6422 29073
rect 6366 28999 6422 29008
rect 6564 26586 6592 32438
rect 7024 31346 7052 40870
rect 7300 35494 7328 41618
rect 7576 40934 7604 43046
rect 7564 40928 7616 40934
rect 7564 40870 7616 40876
rect 7288 35488 7340 35494
rect 7288 35430 7340 35436
rect 7300 34678 7328 35430
rect 7288 34672 7340 34678
rect 7288 34614 7340 34620
rect 7104 34536 7156 34542
rect 7104 34478 7156 34484
rect 7116 34066 7144 34478
rect 7104 34060 7156 34066
rect 7104 34002 7156 34008
rect 7116 33454 7144 34002
rect 7104 33448 7156 33454
rect 7104 33390 7156 33396
rect 7576 33114 7604 40870
rect 7748 40724 7800 40730
rect 7748 40666 7800 40672
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7760 30802 7788 40666
rect 7838 40624 7894 40633
rect 7838 40559 7894 40568
rect 7852 40526 7880 40559
rect 7840 40520 7892 40526
rect 7840 40462 7892 40468
rect 7944 37126 7972 46310
rect 8036 46034 8064 46430
rect 8024 46028 8076 46034
rect 8024 45970 8076 45976
rect 9034 44432 9090 44441
rect 9034 44367 9090 44376
rect 9048 44334 9076 44367
rect 8944 44328 8996 44334
rect 8944 44270 8996 44276
rect 9036 44328 9088 44334
rect 9036 44270 9088 44276
rect 8956 43382 8984 44270
rect 9680 44260 9732 44266
rect 9680 44202 9732 44208
rect 9692 43858 9720 44202
rect 9680 43852 9732 43858
rect 9680 43794 9732 43800
rect 9772 43648 9824 43654
rect 9772 43590 9824 43596
rect 8668 43376 8720 43382
rect 8668 43318 8720 43324
rect 8944 43376 8996 43382
rect 8944 43318 8996 43324
rect 8680 43246 8708 43318
rect 8668 43240 8720 43246
rect 8944 43240 8996 43246
rect 8720 43200 8944 43228
rect 8668 43182 8720 43188
rect 8944 43182 8996 43188
rect 9784 43110 9812 43590
rect 11612 43444 11664 43450
rect 11612 43386 11664 43392
rect 9772 43104 9824 43110
rect 9772 43046 9824 43052
rect 10140 43104 10192 43110
rect 10140 43046 10192 43052
rect 10152 40730 10180 43046
rect 11060 42696 11112 42702
rect 11060 42638 11112 42644
rect 11072 41274 11100 42638
rect 11152 41744 11204 41750
rect 11150 41712 11152 41721
rect 11204 41712 11206 41721
rect 11150 41647 11206 41656
rect 11336 41608 11388 41614
rect 11336 41550 11388 41556
rect 11348 41274 11376 41550
rect 11060 41268 11112 41274
rect 11060 41210 11112 41216
rect 11336 41268 11388 41274
rect 11336 41210 11388 41216
rect 11428 41268 11480 41274
rect 11428 41210 11480 41216
rect 11060 40928 11112 40934
rect 11060 40870 11112 40876
rect 11072 40730 11100 40870
rect 10140 40724 10192 40730
rect 10140 40666 10192 40672
rect 11060 40724 11112 40730
rect 11060 40666 11112 40672
rect 10232 40588 10284 40594
rect 10232 40530 10284 40536
rect 9864 40384 9916 40390
rect 9864 40326 9916 40332
rect 9404 39976 9456 39982
rect 9404 39918 9456 39924
rect 9128 39500 9180 39506
rect 9128 39442 9180 39448
rect 9140 39302 9168 39442
rect 9128 39296 9180 39302
rect 9128 39238 9180 39244
rect 7932 37120 7984 37126
rect 7932 37062 7984 37068
rect 9140 36786 9168 39238
rect 9416 39030 9444 39918
rect 9876 39098 9904 40326
rect 10244 40186 10272 40530
rect 11440 40526 11468 41210
rect 11428 40520 11480 40526
rect 11428 40462 11480 40468
rect 10232 40180 10284 40186
rect 10232 40122 10284 40128
rect 10600 39840 10652 39846
rect 10600 39782 10652 39788
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 9404 39024 9456 39030
rect 9404 38966 9456 38972
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 9692 36242 9720 37198
rect 9876 36922 9904 39034
rect 10232 39024 10284 39030
rect 10232 38966 10284 38972
rect 10244 38894 10272 38966
rect 10232 38888 10284 38894
rect 10232 38830 10284 38836
rect 10244 37806 10272 38830
rect 10612 38418 10640 39782
rect 10600 38412 10652 38418
rect 10600 38354 10652 38360
rect 11060 38344 11112 38350
rect 11060 38286 11112 38292
rect 11072 38010 11100 38286
rect 11060 38004 11112 38010
rect 11060 37946 11112 37952
rect 10968 37868 11020 37874
rect 10968 37810 11020 37816
rect 10232 37800 10284 37806
rect 10232 37742 10284 37748
rect 10508 37732 10560 37738
rect 10508 37674 10560 37680
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 9864 36916 9916 36922
rect 9864 36858 9916 36864
rect 9956 36916 10008 36922
rect 9956 36858 10008 36864
rect 9876 36718 9904 36858
rect 9968 36786 9996 36858
rect 9956 36780 10008 36786
rect 9956 36722 10008 36728
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 9772 36644 9824 36650
rect 9772 36586 9824 36592
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 9784 36106 9812 36586
rect 10336 36106 10364 37266
rect 10520 37262 10548 37674
rect 10980 37466 11008 37810
rect 10968 37460 11020 37466
rect 10968 37402 11020 37408
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 10876 37324 10928 37330
rect 10980 37312 11008 37402
rect 10928 37284 11008 37312
rect 10876 37266 10928 37272
rect 11072 37262 11100 37402
rect 10508 37256 10560 37262
rect 10508 37198 10560 37204
rect 11060 37256 11112 37262
rect 11060 37198 11112 37204
rect 11072 36922 11100 37198
rect 11060 36916 11112 36922
rect 11060 36858 11112 36864
rect 9772 36100 9824 36106
rect 9772 36042 9824 36048
rect 10324 36100 10376 36106
rect 10324 36042 10376 36048
rect 9404 35760 9456 35766
rect 9404 35702 9456 35708
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 9036 34468 9088 34474
rect 9036 34410 9088 34416
rect 8944 33380 8996 33386
rect 8944 33322 8996 33328
rect 8024 33312 8076 33318
rect 8024 33254 8076 33260
rect 8036 32978 8064 33254
rect 8956 33114 8984 33322
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8956 32978 8984 33050
rect 8024 32972 8076 32978
rect 8024 32914 8076 32920
rect 8944 32972 8996 32978
rect 8944 32914 8996 32920
rect 8036 32366 8064 32914
rect 8668 32904 8720 32910
rect 8668 32846 8720 32852
rect 8484 32428 8536 32434
rect 8484 32370 8536 32376
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 7748 30796 7800 30802
rect 7748 30738 7800 30744
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 6656 29782 6684 30534
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 7760 29782 7788 29990
rect 6644 29776 6696 29782
rect 6644 29718 6696 29724
rect 7748 29776 7800 29782
rect 7748 29718 7800 29724
rect 8496 29714 8524 32370
rect 8484 29708 8536 29714
rect 8484 29650 8536 29656
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 8220 27878 8248 28426
rect 8312 28422 8340 28562
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 7288 27532 7340 27538
rect 7288 27474 7340 27480
rect 7300 27130 7328 27474
rect 8220 27402 8248 27814
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 7932 26784 7984 26790
rect 7932 26726 7984 26732
rect 8024 26784 8076 26790
rect 8024 26726 8076 26732
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 6552 26580 6604 26586
rect 6552 26522 6604 26528
rect 5828 26450 5856 26522
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5368 24750 5396 26318
rect 7944 25702 7972 26726
rect 8036 26246 8064 26726
rect 8024 26240 8076 26246
rect 8024 26182 8076 26188
rect 8036 25888 8064 26182
rect 8036 25860 8156 25888
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 6092 25288 6144 25294
rect 6092 25230 6144 25236
rect 5356 24744 5408 24750
rect 5356 24686 5408 24692
rect 5908 24676 5960 24682
rect 5908 24618 5960 24624
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5552 23118 5580 23598
rect 5644 23254 5672 24210
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5644 21486 5672 23190
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5644 20398 5672 21422
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5000 19514 5028 19654
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4908 12850 4936 14214
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 5000 12306 5028 19450
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5644 8090 5672 8910
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 5920 4146 5948 24618
rect 6104 24410 6132 25230
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7208 24886 7236 25094
rect 7196 24880 7248 24886
rect 7196 24822 7248 24828
rect 7208 24750 7236 24822
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6092 24404 6144 24410
rect 6092 24346 6144 24352
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 6104 23186 6132 23462
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6012 19922 6040 20198
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 6196 14074 6224 24550
rect 6932 24274 6960 24550
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 7472 21888 7524 21894
rect 7472 21830 7524 21836
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6288 18834 6316 19722
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6380 14958 6408 15370
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6196 13530 6224 14010
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6564 6798 6592 21830
rect 7484 21146 7512 21830
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6932 19310 6960 19858
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7024 17134 7052 20198
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 18970 7236 19110
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7024 15570 7052 17070
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7300 16658 7328 16934
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7116 16114 7144 16594
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7484 15706 7512 15982
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6840 13870 6868 14010
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 7576 13530 7604 21082
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 17134 7788 17478
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7852 16946 7880 19110
rect 7760 16918 7880 16946
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7024 11694 7052 12242
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 9586 6960 11086
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7116 8498 7144 13126
rect 7300 12442 7328 13398
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7484 11150 7512 12242
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7392 10606 7420 11018
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 9110 7420 10542
rect 7484 9518 7512 11086
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7760 9382 7788 16918
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7852 10674 7880 12922
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7852 9178 7880 9454
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7392 8498 7420 9046
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 8090 7420 8434
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7410 7420 8026
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 3976 2984 4028 2990
rect 3330 2952 3386 2961
rect 3976 2926 4028 2932
rect 3330 2887 3386 2896
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 921 2820 2790
rect 5000 2310 5028 3878
rect 7944 3670 7972 25638
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 8036 21554 8064 22170
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 2872 2304 2924 2310
rect 2870 2272 2872 2281
rect 4988 2304 5040 2310
rect 2924 2272 2926 2281
rect 4988 2246 5040 2252
rect 2870 2207 2926 2216
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 8036 1766 8064 17750
rect 8128 17678 8156 25860
rect 8220 17814 8248 27338
rect 8312 27062 8340 28358
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 8300 26784 8352 26790
rect 8300 26726 8352 26732
rect 8312 26450 8340 26726
rect 8404 26586 8432 27406
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8300 26240 8352 26246
rect 8298 26208 8300 26217
rect 8352 26208 8354 26217
rect 8298 26143 8354 26152
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 8404 20346 8432 22646
rect 8496 22574 8524 22714
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 8576 22432 8628 22438
rect 8576 22374 8628 22380
rect 8588 22098 8616 22374
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8404 20318 8524 20346
rect 8392 20256 8444 20262
rect 8312 20204 8392 20210
rect 8312 20198 8444 20204
rect 8312 20182 8432 20198
rect 8312 19990 8340 20182
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8312 19310 8340 19926
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 12764 8156 17478
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 13734 8248 14350
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8404 13938 8432 14282
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13326 8248 13670
rect 8496 13394 8524 20318
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17066 8616 17478
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 16794 8616 17002
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8680 16250 8708 32846
rect 8760 22500 8812 22506
rect 8760 22442 8812 22448
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8772 13870 8800 22442
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 16250 8984 16526
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 9048 14346 9076 34410
rect 9324 34202 9352 35566
rect 9312 34196 9364 34202
rect 9312 34138 9364 34144
rect 9312 33584 9364 33590
rect 9312 33526 9364 33532
rect 9324 33454 9352 33526
rect 9312 33448 9364 33454
rect 9312 33390 9364 33396
rect 9220 33312 9272 33318
rect 9220 33254 9272 33260
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12918 8248 13262
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8128 12736 8248 12764
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8128 10062 8156 10542
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9586 8156 9998
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 6866 8156 7822
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 8024 1760 8076 1766
rect 8024 1702 8076 1708
rect 3252 1601 3280 1702
rect 3238 1592 3294 1601
rect 3238 1527 3294 1536
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 8220 746 8248 12736
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8404 11898 8432 12650
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8404 10810 8432 11630
rect 8496 11098 8524 13126
rect 9140 12986 9168 19994
rect 9232 18426 9260 33254
rect 9416 32434 9444 35702
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9588 34060 9640 34066
rect 9588 34002 9640 34008
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9600 31142 9628 34002
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9600 30190 9628 31078
rect 9588 30184 9640 30190
rect 9588 30126 9640 30132
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9692 29714 9720 29990
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9692 29510 9720 29650
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 9600 28218 9628 28698
rect 9876 28506 9904 35430
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 9956 32564 10008 32570
rect 9956 32506 10008 32512
rect 9968 32366 9996 32506
rect 10048 32428 10100 32434
rect 10048 32370 10100 32376
rect 9956 32360 10008 32366
rect 9956 32302 10008 32308
rect 9956 30116 10008 30122
rect 9956 30058 10008 30064
rect 9968 29714 9996 30058
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 9876 28478 9996 28506
rect 9864 28416 9916 28422
rect 9864 28358 9916 28364
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9600 27334 9628 28154
rect 9876 28150 9904 28358
rect 9864 28144 9916 28150
rect 9864 28086 9916 28092
rect 9680 27872 9732 27878
rect 9732 27820 9812 27826
rect 9680 27814 9812 27820
rect 9692 27798 9812 27814
rect 9784 27402 9812 27798
rect 9864 27532 9916 27538
rect 9864 27474 9916 27480
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9784 26790 9812 27338
rect 9876 27130 9904 27474
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9876 26926 9904 27066
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9876 26042 9904 26862
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9968 25974 9996 28478
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9324 21690 9352 22714
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 18834 9996 19314
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9692 18086 9720 18702
rect 10060 18306 10088 32370
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 10152 27520 10180 27950
rect 10232 27532 10284 27538
rect 10152 27492 10232 27520
rect 10152 26926 10180 27492
rect 10232 27474 10284 27480
rect 10140 26920 10192 26926
rect 10140 26862 10192 26868
rect 10152 26586 10180 26862
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 9784 18278 10088 18306
rect 9680 18080 9732 18086
rect 9600 18028 9680 18034
rect 9600 18022 9732 18028
rect 9600 18006 9720 18022
rect 9600 16590 9628 18006
rect 9784 17338 9812 18278
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9876 17338 9904 18158
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15570 9812 15846
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 10428 15162 10456 32846
rect 10796 32570 10824 33254
rect 10784 32564 10836 32570
rect 10784 32506 10836 32512
rect 11244 31816 11296 31822
rect 11244 31758 11296 31764
rect 11256 30870 11284 31758
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 11624 30784 11652 43386
rect 12084 39642 12112 46922
rect 13372 46578 13400 46922
rect 13740 46578 13768 47534
rect 14004 46980 14056 46986
rect 14004 46922 14056 46928
rect 14188 46980 14240 46986
rect 14188 46922 14240 46928
rect 14016 46646 14044 46922
rect 14004 46640 14056 46646
rect 14004 46582 14056 46588
rect 13360 46572 13412 46578
rect 13360 46514 13412 46520
rect 13728 46572 13780 46578
rect 13728 46514 13780 46520
rect 13452 46504 13504 46510
rect 13452 46446 13504 46452
rect 13464 45490 13492 46446
rect 13912 46368 13964 46374
rect 13912 46310 13964 46316
rect 13924 46034 13952 46310
rect 14016 46170 14044 46582
rect 14004 46164 14056 46170
rect 14004 46106 14056 46112
rect 14200 46034 14228 46922
rect 13912 46028 13964 46034
rect 13912 45970 13964 45976
rect 14188 46028 14240 46034
rect 14188 45970 14240 45976
rect 13452 45484 13504 45490
rect 13452 45426 13504 45432
rect 13464 44334 13492 45426
rect 13820 45416 13872 45422
rect 13820 45358 13872 45364
rect 13452 44328 13504 44334
rect 13452 44270 13504 44276
rect 12716 43716 12768 43722
rect 12716 43658 12768 43664
rect 12900 43716 12952 43722
rect 12900 43658 12952 43664
rect 12728 43450 12756 43658
rect 12716 43444 12768 43450
rect 12716 43386 12768 43392
rect 12912 43246 12940 43658
rect 12900 43240 12952 43246
rect 12900 43182 12952 43188
rect 13464 41818 13492 44270
rect 13832 43994 13860 45358
rect 14004 44328 14056 44334
rect 14004 44270 14056 44276
rect 13820 43988 13872 43994
rect 13820 43930 13872 43936
rect 14016 43450 14044 44270
rect 14280 43920 14332 43926
rect 14280 43862 14332 43868
rect 14004 43444 14056 43450
rect 14004 43386 14056 43392
rect 13636 43172 13688 43178
rect 13636 43114 13688 43120
rect 13648 42702 13676 43114
rect 14292 42770 14320 43862
rect 13728 42764 13780 42770
rect 13728 42706 13780 42712
rect 14004 42764 14056 42770
rect 14004 42706 14056 42712
rect 14280 42764 14332 42770
rect 14280 42706 14332 42712
rect 13636 42696 13688 42702
rect 13636 42638 13688 42644
rect 13740 42294 13768 42706
rect 13728 42288 13780 42294
rect 13728 42230 13780 42236
rect 13452 41812 13504 41818
rect 13504 41772 13584 41800
rect 13452 41754 13504 41760
rect 12532 41472 12584 41478
rect 12532 41414 12584 41420
rect 12544 40594 12572 41414
rect 12716 41064 12768 41070
rect 12716 41006 12768 41012
rect 13452 41064 13504 41070
rect 13452 41006 13504 41012
rect 12728 40730 12756 41006
rect 13084 40928 13136 40934
rect 13084 40870 13136 40876
rect 12716 40724 12768 40730
rect 12716 40666 12768 40672
rect 13096 40662 13124 40870
rect 13464 40730 13492 41006
rect 13452 40724 13504 40730
rect 13452 40666 13504 40672
rect 13556 40662 13584 41772
rect 13740 41070 13768 42230
rect 14016 41818 14044 42706
rect 14004 41812 14056 41818
rect 14004 41754 14056 41760
rect 14016 41070 14044 41754
rect 13728 41064 13780 41070
rect 13728 41006 13780 41012
rect 14004 41064 14056 41070
rect 14004 41006 14056 41012
rect 13084 40656 13136 40662
rect 13084 40598 13136 40604
rect 13544 40656 13596 40662
rect 13544 40598 13596 40604
rect 12532 40588 12584 40594
rect 12532 40530 12584 40536
rect 12532 40384 12584 40390
rect 12532 40326 12584 40332
rect 12544 40118 12572 40326
rect 12532 40112 12584 40118
rect 12532 40054 12584 40060
rect 12072 39636 12124 39642
rect 12072 39578 12124 39584
rect 13556 39098 13584 40598
rect 13544 39092 13596 39098
rect 13544 39034 13596 39040
rect 13820 39092 13872 39098
rect 13820 39034 13872 39040
rect 12256 38480 12308 38486
rect 12256 38422 12308 38428
rect 12268 38214 12296 38422
rect 13832 38418 13860 39034
rect 13820 38412 13872 38418
rect 13820 38354 13872 38360
rect 12256 38208 12308 38214
rect 12256 38150 12308 38156
rect 12440 38208 12492 38214
rect 12440 38150 12492 38156
rect 12452 37806 12480 38150
rect 12530 37904 12586 37913
rect 12530 37839 12532 37848
rect 12584 37839 12586 37848
rect 12532 37810 12584 37816
rect 12440 37800 12492 37806
rect 12440 37742 12492 37748
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 14292 36718 14320 37062
rect 13544 36712 13596 36718
rect 13544 36654 13596 36660
rect 14280 36712 14332 36718
rect 14280 36654 14332 36660
rect 13556 35630 13584 36654
rect 13636 36576 13688 36582
rect 13636 36518 13688 36524
rect 13648 35698 13676 36518
rect 13636 35692 13688 35698
rect 13636 35634 13688 35640
rect 13544 35624 13596 35630
rect 13544 35566 13596 35572
rect 12716 35556 12768 35562
rect 12716 35498 12768 35504
rect 11704 34196 11756 34202
rect 11704 34138 11756 34144
rect 11716 33998 11744 34138
rect 11704 33992 11756 33998
rect 11704 33934 11756 33940
rect 11716 33046 11744 33934
rect 11704 33040 11756 33046
rect 11704 32982 11756 32988
rect 11716 32026 11744 32982
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 12452 30870 12480 31690
rect 12348 30864 12400 30870
rect 12348 30806 12400 30812
rect 12440 30864 12492 30870
rect 12440 30806 12492 30812
rect 12532 30864 12584 30870
rect 12532 30806 12584 30812
rect 11796 30796 11848 30802
rect 11624 30756 11796 30784
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10704 30054 10732 30330
rect 11164 30190 11192 30670
rect 11716 30598 11744 30756
rect 11796 30738 11848 30744
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 11716 30054 11744 30534
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 11704 30048 11756 30054
rect 11704 29990 11756 29996
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11900 29714 11928 29990
rect 11888 29708 11940 29714
rect 11888 29650 11940 29656
rect 11900 29170 11928 29650
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 12360 29102 12388 30806
rect 12544 30666 12572 30806
rect 12624 30796 12676 30802
rect 12624 30738 12676 30744
rect 12532 30660 12584 30666
rect 12532 30602 12584 30608
rect 12636 30190 12664 30738
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 10692 28620 10744 28626
rect 10692 28562 10744 28568
rect 10704 28082 10732 28562
rect 12728 28422 12756 35498
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13176 34400 13228 34406
rect 13176 34342 13228 34348
rect 13188 34066 13216 34342
rect 13176 34060 13228 34066
rect 13176 34002 13228 34008
rect 12900 33584 12952 33590
rect 12898 33552 12900 33561
rect 12952 33552 12954 33561
rect 12898 33487 12954 33496
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 12912 30938 12940 31078
rect 13004 30938 13032 31622
rect 12900 30932 12952 30938
rect 12900 30874 12952 30880
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 13464 29850 13492 35430
rect 13912 35148 13964 35154
rect 13912 35090 13964 35096
rect 13924 34950 13952 35090
rect 13912 34944 13964 34950
rect 13912 34886 13964 34892
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13832 34202 13860 34478
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 13924 33862 13952 34886
rect 14200 34678 14228 34886
rect 14188 34672 14240 34678
rect 14188 34614 14240 34620
rect 13912 33856 13964 33862
rect 13912 33798 13964 33804
rect 14936 33590 14964 48350
rect 18052 47048 18104 47054
rect 18052 46990 18104 46996
rect 15476 46912 15528 46918
rect 15476 46854 15528 46860
rect 15488 45490 15516 46854
rect 18064 45966 18092 46990
rect 18156 46510 18184 49248
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 22468 47456 22520 47462
rect 22468 47398 22520 47404
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 22480 47258 22508 47398
rect 50300 47356 50596 47376
rect 50356 47354 50380 47356
rect 50436 47354 50460 47356
rect 50516 47354 50540 47356
rect 50378 47302 50380 47354
rect 50442 47302 50454 47354
rect 50516 47302 50518 47354
rect 50356 47300 50380 47302
rect 50436 47300 50460 47302
rect 50516 47300 50540 47302
rect 50300 47280 50596 47300
rect 22284 47252 22336 47258
rect 22284 47194 22336 47200
rect 22468 47252 22520 47258
rect 22468 47194 22520 47200
rect 19064 46912 19116 46918
rect 19064 46854 19116 46860
rect 19076 46510 19104 46854
rect 22296 46714 22324 47194
rect 23296 47184 23348 47190
rect 23296 47126 23348 47132
rect 22284 46708 22336 46714
rect 22284 46650 22336 46656
rect 23308 46510 23336 47126
rect 23388 47116 23440 47122
rect 23388 47058 23440 47064
rect 25412 47116 25464 47122
rect 25412 47058 25464 47064
rect 44364 47116 44416 47122
rect 44364 47058 44416 47064
rect 46664 47116 46716 47122
rect 46664 47058 46716 47064
rect 50160 47116 50212 47122
rect 50160 47058 50212 47064
rect 50528 47116 50580 47122
rect 50528 47058 50580 47064
rect 50896 47116 50948 47122
rect 50896 47058 50948 47064
rect 51908 47116 51960 47122
rect 51908 47058 51960 47064
rect 23400 46986 23428 47058
rect 23388 46980 23440 46986
rect 23388 46922 23440 46928
rect 23940 46980 23992 46986
rect 23940 46922 23992 46928
rect 18144 46504 18196 46510
rect 18144 46446 18196 46452
rect 19064 46504 19116 46510
rect 19064 46446 19116 46452
rect 20720 46504 20772 46510
rect 20720 46446 20772 46452
rect 23296 46504 23348 46510
rect 23296 46446 23348 46452
rect 18144 46368 18196 46374
rect 18144 46310 18196 46316
rect 19156 46368 19208 46374
rect 19156 46310 19208 46316
rect 18052 45960 18104 45966
rect 18052 45902 18104 45908
rect 16764 45892 16816 45898
rect 16764 45834 16816 45840
rect 15660 45552 15712 45558
rect 15660 45494 15712 45500
rect 15476 45484 15528 45490
rect 15476 45426 15528 45432
rect 15292 45076 15344 45082
rect 15292 45018 15344 45024
rect 15304 44470 15332 45018
rect 15488 44470 15516 45426
rect 15292 44464 15344 44470
rect 15292 44406 15344 44412
rect 15476 44464 15528 44470
rect 15476 44406 15528 44412
rect 15304 43450 15332 44406
rect 15672 43994 15700 45494
rect 15660 43988 15712 43994
rect 15660 43930 15712 43936
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 15304 43246 15332 43386
rect 16580 43308 16632 43314
rect 16580 43250 16632 43256
rect 15292 43240 15344 43246
rect 15292 43182 15344 43188
rect 16592 43178 16620 43250
rect 16580 43172 16632 43178
rect 16580 43114 16632 43120
rect 16396 42764 16448 42770
rect 16396 42706 16448 42712
rect 16212 42016 16264 42022
rect 16212 41958 16264 41964
rect 16224 41818 16252 41958
rect 16408 41818 16436 42706
rect 16212 41812 16264 41818
rect 16212 41754 16264 41760
rect 16396 41812 16448 41818
rect 16396 41754 16448 41760
rect 16408 41682 16436 41754
rect 16120 41676 16172 41682
rect 16120 41618 16172 41624
rect 16396 41676 16448 41682
rect 16396 41618 16448 41624
rect 16028 40520 16080 40526
rect 16028 40462 16080 40468
rect 15568 39908 15620 39914
rect 15568 39850 15620 39856
rect 15108 39840 15160 39846
rect 15108 39782 15160 39788
rect 15120 39030 15148 39782
rect 15108 39024 15160 39030
rect 15108 38966 15160 38972
rect 15120 38894 15148 38966
rect 15580 38894 15608 39850
rect 16040 39030 16068 40462
rect 16028 39024 16080 39030
rect 16028 38966 16080 38972
rect 15108 38888 15160 38894
rect 15108 38830 15160 38836
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15108 38752 15160 38758
rect 15108 38694 15160 38700
rect 15120 38214 15148 38694
rect 15108 38208 15160 38214
rect 15108 38150 15160 38156
rect 14924 33584 14976 33590
rect 14924 33526 14976 33532
rect 14936 33454 14964 33526
rect 14924 33448 14976 33454
rect 14924 33390 14976 33396
rect 13452 29844 13504 29850
rect 13452 29786 13504 29792
rect 14936 29102 14964 33390
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 13268 29028 13320 29034
rect 13268 28970 13320 28976
rect 14004 29028 14056 29034
rect 14004 28970 14056 28976
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10692 27464 10744 27470
rect 10692 27406 10744 27412
rect 10704 27130 10732 27406
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10704 27010 10732 27066
rect 10612 26982 10732 27010
rect 10612 26518 10640 26982
rect 10692 26852 10744 26858
rect 10692 26794 10744 26800
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10704 26450 10732 26794
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 11072 25294 11100 28154
rect 12624 27940 12676 27946
rect 12624 27882 12676 27888
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12544 26994 12572 27474
rect 12636 27334 12664 27882
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11624 25498 11652 26250
rect 12728 25974 12756 28358
rect 12716 25968 12768 25974
rect 12636 25916 12716 25922
rect 12636 25910 12768 25916
rect 12636 25894 12756 25910
rect 11612 25492 11664 25498
rect 11612 25434 11664 25440
rect 12164 25424 12216 25430
rect 12164 25366 12216 25372
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11072 21962 11100 25230
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11532 24274 11560 25162
rect 12176 25158 12204 25366
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10520 13530 10548 21286
rect 11072 20874 11100 21898
rect 11164 21486 11192 24006
rect 12176 22098 12204 25094
rect 12636 24750 12664 25894
rect 12728 25845 12756 25894
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12728 24954 12756 25094
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12820 24750 12848 25298
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12636 23322 12664 24686
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12728 23662 12756 24006
rect 12820 23798 12848 24686
rect 12808 23792 12860 23798
rect 12808 23734 12860 23740
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12728 23526 12756 23598
rect 12716 23520 12768 23526
rect 12714 23488 12716 23497
rect 12768 23488 12770 23497
rect 12714 23423 12770 23432
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13188 22166 13216 23054
rect 13176 22160 13228 22166
rect 13176 22102 13228 22108
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12728 21554 12756 21830
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 19922 11468 20198
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10704 19174 10732 19246
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10704 18630 10732 19110
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 11256 18426 11284 19654
rect 12176 18766 12204 19722
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 18834 12480 19654
rect 13004 19446 13032 19858
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12986 9812 13262
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9140 12782 9168 12922
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 8496 11070 8616 11098
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8404 10130 8432 10746
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8496 10062 8524 10950
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8496 9518 8524 9998
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8588 6322 8616 11070
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8864 10810 8892 11018
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 8634 9904 10066
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8772 7546 8800 8366
rect 9784 7546 9812 8434
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8772 6866 8800 7278
rect 9784 7274 9812 7482
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 9968 4690 9996 13126
rect 10612 12442 10640 13874
rect 10796 13870 10824 17274
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12442 11100 12582
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11164 11762 11192 12650
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11256 10742 11284 18362
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 12360 16250 12388 16662
rect 13096 16658 13124 17546
rect 13280 16658 13308 28970
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13912 28620 13964 28626
rect 13912 28562 13964 28568
rect 13832 28150 13860 28562
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13832 27878 13860 28086
rect 13924 28082 13952 28562
rect 14016 28558 14044 28970
rect 14832 28960 14884 28966
rect 14832 28902 14884 28908
rect 14924 28960 14976 28966
rect 14924 28902 14976 28908
rect 14844 28626 14872 28902
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27674 13860 27814
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13634 27568 13690 27577
rect 13924 27538 13952 28018
rect 14016 27946 14044 28494
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 13634 27503 13636 27512
rect 13688 27503 13690 27512
rect 13912 27532 13964 27538
rect 13636 27474 13688 27480
rect 13912 27474 13964 27480
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13740 26926 13768 27338
rect 13924 27334 13952 27474
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 14016 26926 14044 27882
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13556 24750 13584 25094
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13556 24138 13584 24686
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13556 23186 13584 24074
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13924 23662 13952 23734
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13740 23186 13768 23258
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 13832 22778 13860 23530
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 21690 13584 22578
rect 13924 22574 13952 22986
rect 14108 22574 14136 28494
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14200 27538 14228 27610
rect 14188 27532 14240 27538
rect 14188 27474 14240 27480
rect 14292 23662 14320 27950
rect 14476 27946 14504 28018
rect 14464 27940 14516 27946
rect 14464 27882 14516 27888
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14384 27554 14412 27814
rect 14384 27538 14504 27554
rect 14384 27532 14516 27538
rect 14384 27526 14464 27532
rect 14464 27474 14516 27480
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22574 14320 23122
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 14108 21894 14136 22034
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 14108 21418 14136 21830
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14108 21321 14136 21354
rect 14094 21312 14150 21321
rect 14094 21247 14150 21256
rect 14384 20466 14412 27406
rect 14844 26926 14872 28562
rect 14936 28150 14964 28902
rect 15120 28762 15148 38150
rect 15580 37330 15608 38830
rect 15844 38412 15896 38418
rect 15844 38354 15896 38360
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 15856 38214 15884 38354
rect 15844 38208 15896 38214
rect 15844 38150 15896 38156
rect 15856 37942 15884 38150
rect 15844 37936 15896 37942
rect 15844 37878 15896 37884
rect 16040 37874 16068 38354
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 16132 37330 16160 41618
rect 16592 41206 16620 43114
rect 16672 42356 16724 42362
rect 16672 42298 16724 42304
rect 16684 42158 16712 42298
rect 16672 42152 16724 42158
rect 16672 42094 16724 42100
rect 16580 41200 16632 41206
rect 16580 41142 16632 41148
rect 16592 39846 16620 41142
rect 16580 39840 16632 39846
rect 16580 39782 16632 39788
rect 16396 39432 16448 39438
rect 16396 39374 16448 39380
rect 16212 38412 16264 38418
rect 16212 38354 16264 38360
rect 15568 37324 15620 37330
rect 15568 37266 15620 37272
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 15292 36712 15344 36718
rect 15292 36654 15344 36660
rect 15304 36242 15332 36654
rect 16028 36576 16080 36582
rect 16028 36518 16080 36524
rect 15292 36236 15344 36242
rect 15292 36178 15344 36184
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 15212 36038 15240 36110
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15212 35562 15240 35974
rect 16040 35698 16068 36518
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 16132 35630 16160 37266
rect 16224 36242 16252 38354
rect 16408 38282 16436 39374
rect 16396 38276 16448 38282
rect 16396 38218 16448 38224
rect 16684 36854 16712 42094
rect 16776 41274 16804 45834
rect 17224 43988 17276 43994
rect 17224 43930 17276 43936
rect 17132 43784 17184 43790
rect 17132 43726 17184 43732
rect 16764 41268 16816 41274
rect 16764 41210 16816 41216
rect 17144 40050 17172 43726
rect 17236 42838 17264 43930
rect 17776 43104 17828 43110
rect 17776 43046 17828 43052
rect 17868 43104 17920 43110
rect 17868 43046 17920 43052
rect 17224 42832 17276 42838
rect 17224 42774 17276 42780
rect 17408 42084 17460 42090
rect 17408 42026 17460 42032
rect 17420 41138 17448 42026
rect 17408 41132 17460 41138
rect 17408 41074 17460 41080
rect 17132 40044 17184 40050
rect 17132 39986 17184 39992
rect 17316 39976 17368 39982
rect 17316 39918 17368 39924
rect 17328 39846 17356 39918
rect 17316 39840 17368 39846
rect 17316 39782 17368 39788
rect 17132 39092 17184 39098
rect 17132 39034 17184 39040
rect 17144 37330 17172 39034
rect 17328 37670 17356 39782
rect 17316 37664 17368 37670
rect 17316 37606 17368 37612
rect 17132 37324 17184 37330
rect 17132 37266 17184 37272
rect 16396 36848 16448 36854
rect 16672 36848 16724 36854
rect 16448 36796 16528 36802
rect 16396 36790 16528 36796
rect 16672 36790 16724 36796
rect 16408 36774 16528 36790
rect 16500 36768 16528 36774
rect 16580 36780 16632 36786
rect 16500 36740 16580 36768
rect 16580 36722 16632 36728
rect 16684 36650 16712 36790
rect 16672 36644 16724 36650
rect 16672 36586 16724 36592
rect 16684 36378 16712 36586
rect 17144 36378 17172 37266
rect 16672 36372 16724 36378
rect 16672 36314 16724 36320
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 16212 36236 16264 36242
rect 16212 36178 16264 36184
rect 16684 36174 16712 36314
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16684 35714 16712 36110
rect 17512 36038 17540 36178
rect 17500 36032 17552 36038
rect 17500 35974 17552 35980
rect 16684 35686 16804 35714
rect 16120 35624 16172 35630
rect 16120 35566 16172 35572
rect 15200 35556 15252 35562
rect 15200 35498 15252 35504
rect 16672 35556 16724 35562
rect 16672 35498 16724 35504
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16500 35086 16528 35430
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 16684 34678 16712 35498
rect 16776 35494 16804 35686
rect 16764 35488 16816 35494
rect 16764 35430 16816 35436
rect 17316 35284 17368 35290
rect 17316 35226 17368 35232
rect 17224 34944 17276 34950
rect 17224 34886 17276 34892
rect 15752 34672 15804 34678
rect 16672 34672 16724 34678
rect 15752 34614 15804 34620
rect 15764 34542 15792 34614
rect 16132 34598 16620 34626
rect 16672 34614 16724 34620
rect 16132 34542 16160 34598
rect 16592 34542 16620 34598
rect 15752 34536 15804 34542
rect 15752 34478 15804 34484
rect 15844 34536 15896 34542
rect 15844 34478 15896 34484
rect 16120 34536 16172 34542
rect 16120 34478 16172 34484
rect 16212 34536 16264 34542
rect 16212 34478 16264 34484
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 15568 34468 15620 34474
rect 15568 34410 15620 34416
rect 15580 34066 15608 34410
rect 15568 34060 15620 34066
rect 15568 34002 15620 34008
rect 15856 32502 15884 34478
rect 16224 33454 16252 34478
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16684 34134 16712 34342
rect 16672 34128 16724 34134
rect 16672 34070 16724 34076
rect 16488 34060 16540 34066
rect 16488 34002 16540 34008
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16396 33924 16448 33930
rect 16396 33866 16448 33872
rect 16212 33448 16264 33454
rect 16212 33390 16264 33396
rect 16408 33318 16436 33866
rect 16500 33862 16528 34002
rect 16488 33856 16540 33862
rect 16488 33798 16540 33804
rect 16672 33448 16724 33454
rect 16868 33436 16896 34002
rect 17236 33862 17264 34886
rect 17224 33856 17276 33862
rect 17224 33798 17276 33804
rect 17328 33590 17356 35226
rect 17316 33584 17368 33590
rect 17316 33526 17368 33532
rect 17328 33454 17356 33526
rect 16724 33408 16896 33436
rect 17316 33448 17368 33454
rect 16672 33390 16724 33396
rect 17316 33390 17368 33396
rect 16396 33312 16448 33318
rect 16396 33254 16448 33260
rect 16488 33312 16540 33318
rect 16488 33254 16540 33260
rect 15844 32496 15896 32502
rect 15844 32438 15896 32444
rect 15660 32360 15712 32366
rect 15660 32302 15712 32308
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 15396 30666 15424 31758
rect 15672 31278 15700 32302
rect 16120 31952 16172 31958
rect 16120 31894 16172 31900
rect 16132 31346 16160 31894
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16396 31340 16448 31346
rect 16396 31282 16448 31288
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15568 31204 15620 31210
rect 15568 31146 15620 31152
rect 15384 30660 15436 30666
rect 15384 30602 15436 30608
rect 15396 29850 15424 30602
rect 15580 30190 15608 31146
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 15396 28762 15424 29786
rect 15580 29714 15608 29990
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15108 28756 15160 28762
rect 15108 28698 15160 28704
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14936 27878 14964 28086
rect 15120 28082 15240 28098
rect 15120 28076 15252 28082
rect 15120 28070 15200 28076
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 15120 26926 15148 28070
rect 15200 28018 15252 28024
rect 15304 27577 15332 28494
rect 15290 27568 15346 27577
rect 15290 27503 15346 27512
rect 15304 27470 15332 27503
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15672 27402 15700 31214
rect 16132 30802 16160 31282
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15764 27946 15792 28562
rect 16132 27946 16160 29650
rect 16408 28218 16436 31282
rect 16500 31210 16528 33254
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16672 32768 16724 32774
rect 16672 32710 16724 32716
rect 16684 32298 16712 32710
rect 16868 32502 16896 32846
rect 16856 32496 16908 32502
rect 16856 32438 16908 32444
rect 16672 32292 16724 32298
rect 16672 32234 16724 32240
rect 17040 31884 17092 31890
rect 17040 31826 17092 31832
rect 17408 31884 17460 31890
rect 17408 31826 17460 31832
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16488 31204 16540 31210
rect 16488 31146 16540 31152
rect 16592 30802 16620 31758
rect 17052 31210 17080 31826
rect 17420 31686 17448 31826
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17040 31204 17092 31210
rect 17040 31146 17092 31152
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16500 30394 16528 30670
rect 17420 30598 17448 31622
rect 17512 31482 17540 35974
rect 17788 35834 17816 43046
rect 17880 42362 17908 43046
rect 17868 42356 17920 42362
rect 17868 42298 17920 42304
rect 17868 39432 17920 39438
rect 17868 39374 17920 39380
rect 17880 38826 17908 39374
rect 17868 38820 17920 38826
rect 17868 38762 17920 38768
rect 17880 38486 17908 38762
rect 17868 38480 17920 38486
rect 17868 38422 17920 38428
rect 17868 37664 17920 37670
rect 17868 37606 17920 37612
rect 17880 35834 17908 37606
rect 17776 35828 17828 35834
rect 17776 35770 17828 35776
rect 17868 35828 17920 35834
rect 17868 35770 17920 35776
rect 18156 35290 18184 46310
rect 19168 46034 19196 46310
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 20732 46034 20760 46446
rect 21916 46436 21968 46442
rect 21916 46378 21968 46384
rect 21824 46368 21876 46374
rect 21824 46310 21876 46316
rect 19156 46028 19208 46034
rect 19156 45970 19208 45976
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 18972 44328 19024 44334
rect 18972 44270 19024 44276
rect 18984 43382 19012 44270
rect 20904 44260 20956 44266
rect 20904 44202 20956 44208
rect 21088 44260 21140 44266
rect 21088 44202 21140 44208
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 20916 43858 20944 44202
rect 20904 43852 20956 43858
rect 20904 43794 20956 43800
rect 20352 43648 20404 43654
rect 20352 43590 20404 43596
rect 20996 43648 21048 43654
rect 20996 43590 21048 43596
rect 18972 43376 19024 43382
rect 18972 43318 19024 43324
rect 19892 43376 19944 43382
rect 19892 43318 19944 43324
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19904 42294 19932 43318
rect 20364 43246 20392 43590
rect 21008 43382 21036 43590
rect 20996 43376 21048 43382
rect 20996 43318 21048 43324
rect 20260 43240 20312 43246
rect 20260 43182 20312 43188
rect 20352 43240 20404 43246
rect 20352 43182 20404 43188
rect 19892 42288 19944 42294
rect 19892 42230 19944 42236
rect 20272 42226 20300 43182
rect 20812 43172 20864 43178
rect 20812 43114 20864 43120
rect 20824 42362 20852 43114
rect 21100 42566 21128 44202
rect 21836 44198 21864 46310
rect 21928 46034 21956 46378
rect 23388 46164 23440 46170
rect 23388 46106 23440 46112
rect 22652 46096 22704 46102
rect 22652 46038 22704 46044
rect 21916 46028 21968 46034
rect 21916 45970 21968 45976
rect 22192 46028 22244 46034
rect 22192 45970 22244 45976
rect 21928 44266 21956 45970
rect 22204 45830 22232 45970
rect 22192 45824 22244 45830
rect 22192 45766 22244 45772
rect 22664 44334 22692 46038
rect 23400 45422 23428 46106
rect 23952 46034 23980 46922
rect 24032 46912 24084 46918
rect 24032 46854 24084 46860
rect 24044 46510 24072 46854
rect 25424 46714 25452 47058
rect 32588 47048 32640 47054
rect 32588 46990 32640 46996
rect 32864 47048 32916 47054
rect 32864 46990 32916 46996
rect 40592 47048 40644 47054
rect 40592 46990 40644 46996
rect 40684 47048 40736 47054
rect 40684 46990 40736 46996
rect 31024 46912 31076 46918
rect 31024 46854 31076 46860
rect 24952 46708 25004 46714
rect 24952 46650 25004 46656
rect 25412 46708 25464 46714
rect 25412 46650 25464 46656
rect 24032 46504 24084 46510
rect 24032 46446 24084 46452
rect 23940 46028 23992 46034
rect 23940 45970 23992 45976
rect 24492 46028 24544 46034
rect 24492 45970 24544 45976
rect 24676 46028 24728 46034
rect 24676 45970 24728 45976
rect 24504 45898 24532 45970
rect 24492 45892 24544 45898
rect 24492 45834 24544 45840
rect 24688 45830 24716 45970
rect 24964 45966 24992 46650
rect 30840 46572 30892 46578
rect 30840 46514 30892 46520
rect 26700 46504 26752 46510
rect 26700 46446 26752 46452
rect 29184 46504 29236 46510
rect 29184 46446 29236 46452
rect 26712 46170 26740 46446
rect 27068 46368 27120 46374
rect 27068 46310 27120 46316
rect 26700 46164 26752 46170
rect 26700 46106 26752 46112
rect 27080 46034 27108 46310
rect 27068 46028 27120 46034
rect 27068 45970 27120 45976
rect 27804 46028 27856 46034
rect 27804 45970 27856 45976
rect 29092 46028 29144 46034
rect 29092 45970 29144 45976
rect 24952 45960 25004 45966
rect 24952 45902 25004 45908
rect 24676 45824 24728 45830
rect 24676 45766 24728 45772
rect 27160 45824 27212 45830
rect 27160 45766 27212 45772
rect 27172 45626 27200 45766
rect 27160 45620 27212 45626
rect 27160 45562 27212 45568
rect 23388 45416 23440 45422
rect 23388 45358 23440 45364
rect 23400 45082 23428 45358
rect 23388 45076 23440 45082
rect 23388 45018 23440 45024
rect 23848 44940 23900 44946
rect 23848 44882 23900 44888
rect 23860 44742 23888 44882
rect 23848 44736 23900 44742
rect 23848 44678 23900 44684
rect 22652 44328 22704 44334
rect 22652 44270 22704 44276
rect 21916 44260 21968 44266
rect 21916 44202 21968 44208
rect 21824 44192 21876 44198
rect 21876 44140 21956 44146
rect 21824 44134 21956 44140
rect 21836 44118 21956 44134
rect 21928 43654 21956 44118
rect 22192 43784 22244 43790
rect 22192 43726 22244 43732
rect 21916 43648 21968 43654
rect 21916 43590 21968 43596
rect 21088 42560 21140 42566
rect 21088 42502 21140 42508
rect 20812 42356 20864 42362
rect 20812 42298 20864 42304
rect 20260 42220 20312 42226
rect 20260 42162 20312 42168
rect 19156 42152 19208 42158
rect 19208 42100 19288 42106
rect 19156 42094 19288 42100
rect 19168 42078 19288 42094
rect 18694 41712 18750 41721
rect 18694 41647 18750 41656
rect 18420 41268 18472 41274
rect 18420 41210 18472 41216
rect 18432 40526 18460 41210
rect 18708 41138 18736 41647
rect 18696 41132 18748 41138
rect 18696 41074 18748 41080
rect 19260 41070 19288 42078
rect 19340 42016 19392 42022
rect 19340 41958 19392 41964
rect 19248 41064 19300 41070
rect 19248 41006 19300 41012
rect 19352 41018 19380 41958
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19432 41812 19484 41818
rect 19432 41754 19484 41760
rect 19444 41138 19472 41754
rect 19432 41132 19484 41138
rect 19432 41074 19484 41080
rect 19260 40662 19288 41006
rect 19352 41002 19472 41018
rect 19352 40996 19484 41002
rect 19352 40990 19432 40996
rect 19432 40938 19484 40944
rect 19248 40656 19300 40662
rect 19248 40598 19300 40604
rect 19444 40610 19472 40938
rect 21824 40928 21876 40934
rect 21822 40896 21824 40905
rect 21876 40896 21878 40905
rect 19580 40828 19876 40848
rect 21822 40831 21878 40840
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 20350 40760 20406 40769
rect 20350 40695 20406 40704
rect 20364 40662 20392 40695
rect 20352 40656 20404 40662
rect 19444 40594 19564 40610
rect 20352 40598 20404 40604
rect 19444 40588 19576 40594
rect 19444 40582 19524 40588
rect 19524 40530 19576 40536
rect 21928 40526 21956 43590
rect 22204 43450 22232 43726
rect 22664 43450 22692 44270
rect 23388 43648 23440 43654
rect 23388 43590 23440 43596
rect 23664 43648 23716 43654
rect 23664 43590 23716 43596
rect 23400 43450 23428 43590
rect 22192 43444 22244 43450
rect 22192 43386 22244 43392
rect 22652 43444 22704 43450
rect 22652 43386 22704 43392
rect 23388 43444 23440 43450
rect 23388 43386 23440 43392
rect 23676 43246 23704 43590
rect 22468 43240 22520 43246
rect 22468 43182 22520 43188
rect 23664 43240 23716 43246
rect 23664 43182 23716 43188
rect 22480 43110 22508 43182
rect 22468 43104 22520 43110
rect 22468 43046 22520 43052
rect 23756 43104 23808 43110
rect 23756 43046 23808 43052
rect 23768 42838 23796 43046
rect 23756 42832 23808 42838
rect 23756 42774 23808 42780
rect 23756 42016 23808 42022
rect 23756 41958 23808 41964
rect 23768 41138 23796 41958
rect 23756 41132 23808 41138
rect 23756 41074 23808 41080
rect 23768 40934 23796 41074
rect 23756 40928 23808 40934
rect 23756 40870 23808 40876
rect 18420 40520 18472 40526
rect 18420 40462 18472 40468
rect 21916 40520 21968 40526
rect 21916 40462 21968 40468
rect 22376 40520 22428 40526
rect 22376 40462 22428 40468
rect 18432 40050 18460 40462
rect 21928 40390 21956 40462
rect 21088 40384 21140 40390
rect 21088 40326 21140 40332
rect 21916 40384 21968 40390
rect 21916 40326 21968 40332
rect 18420 40044 18472 40050
rect 18420 39986 18472 39992
rect 19340 39840 19392 39846
rect 19340 39782 19392 39788
rect 19352 39624 19380 39782
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19260 39596 19380 39624
rect 19260 39302 19288 39596
rect 21100 39506 21128 40326
rect 22388 39642 22416 40462
rect 23664 40384 23716 40390
rect 23664 40326 23716 40332
rect 23676 39982 23704 40326
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 22744 39908 22796 39914
rect 22744 39850 22796 39856
rect 22756 39642 22784 39850
rect 22376 39636 22428 39642
rect 22376 39578 22428 39584
rect 22744 39636 22796 39642
rect 22744 39578 22796 39584
rect 21088 39500 21140 39506
rect 21088 39442 21140 39448
rect 21364 39500 21416 39506
rect 21364 39442 21416 39448
rect 19248 39296 19300 39302
rect 19248 39238 19300 39244
rect 20720 39296 20772 39302
rect 20720 39238 20772 39244
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 20732 37806 20760 39238
rect 21100 38486 21128 39442
rect 21376 39370 21404 39442
rect 21364 39364 21416 39370
rect 21364 39306 21416 39312
rect 21376 38894 21404 39306
rect 22192 39092 22244 39098
rect 22192 39034 22244 39040
rect 21364 38888 21416 38894
rect 21364 38830 21416 38836
rect 20812 38480 20864 38486
rect 20812 38422 20864 38428
rect 21088 38480 21140 38486
rect 21088 38422 21140 38428
rect 20720 37800 20772 37806
rect 20720 37742 20772 37748
rect 20076 37664 20128 37670
rect 20076 37606 20128 37612
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 19260 36718 19288 36858
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 18420 36372 18472 36378
rect 18420 36314 18472 36320
rect 18144 35284 18196 35290
rect 18144 35226 18196 35232
rect 18432 34066 18460 36314
rect 19892 36236 19944 36242
rect 19892 36178 19944 36184
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 19352 34746 19380 36110
rect 19904 35630 19932 36178
rect 19892 35624 19944 35630
rect 19892 35566 19944 35572
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19904 34542 19932 35566
rect 19892 34536 19944 34542
rect 19892 34478 19944 34484
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 18972 34196 19024 34202
rect 18972 34138 19024 34144
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 17972 33318 18000 33798
rect 18064 33454 18092 33934
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 18328 33448 18380 33454
rect 18328 33390 18380 33396
rect 18340 33318 18368 33390
rect 17960 33312 18012 33318
rect 17960 33254 18012 33260
rect 18328 33312 18380 33318
rect 18328 33254 18380 33260
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17972 31822 18000 32234
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 18236 31748 18288 31754
rect 18236 31690 18288 31696
rect 17500 31476 17552 31482
rect 17500 31418 17552 31424
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 16488 30388 16540 30394
rect 16488 30330 16540 30336
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 15752 27940 15804 27946
rect 15752 27882 15804 27888
rect 16120 27940 16172 27946
rect 16120 27882 16172 27888
rect 16132 27674 16160 27882
rect 16120 27668 16172 27674
rect 16120 27610 16172 27616
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15764 26926 15792 27406
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15752 26920 15804 26926
rect 15752 26862 15804 26868
rect 14844 26790 14872 26862
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 15764 26518 15792 26862
rect 15752 26512 15804 26518
rect 15752 26454 15804 26460
rect 15948 26042 15976 27066
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15948 25838 15976 25978
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15856 25294 15884 25638
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14476 23662 14504 24618
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14554 22808 14610 22817
rect 14554 22743 14610 22752
rect 14568 22574 14596 22743
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14476 20346 14504 20470
rect 14384 20318 14504 20346
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18630 13768 19110
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17134 13400 17614
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 17270 13584 17478
rect 13544 17264 13596 17270
rect 13832 17218 13860 18022
rect 13544 17206 13596 17212
rect 13648 17202 13860 17218
rect 13636 17196 13860 17202
rect 13688 17190 13860 17196
rect 13636 17138 13688 17144
rect 14384 17134 14412 20318
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 18970 14688 20198
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 13360 17128 13412 17134
rect 14188 17128 14240 17134
rect 13360 17070 13412 17076
rect 14186 17096 14188 17105
rect 14372 17128 14424 17134
rect 14240 17096 14242 17105
rect 14372 17070 14424 17076
rect 14186 17031 14242 17040
rect 13450 16688 13506 16697
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13268 16652 13320 16658
rect 14384 16658 14412 17070
rect 13450 16623 13452 16632
rect 13268 16594 13320 16600
rect 13504 16623 13506 16632
rect 14372 16652 14424 16658
rect 13452 16594 13504 16600
rect 14372 16594 14424 16600
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12452 14482 12480 16594
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 12636 14822 12664 15846
rect 13924 15026 13952 15846
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12636 14278 12664 14758
rect 14752 14550 14780 25162
rect 15948 24750 15976 25774
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16224 25362 16252 25638
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 16316 23798 16344 27406
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 14844 23497 14872 23598
rect 14830 23488 14886 23497
rect 14830 23423 14886 23432
rect 15120 22574 15148 23598
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15120 21894 15148 22510
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15120 20534 15148 21830
rect 15212 21350 15240 23666
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15212 20398 15240 20538
rect 15764 20466 15792 21286
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15212 17134 15240 20334
rect 15580 20262 15608 20334
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 15580 20097 15608 20198
rect 15566 20088 15622 20097
rect 16132 20058 16160 20198
rect 15566 20023 15622 20032
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16224 18970 16252 20810
rect 16592 20602 16620 29038
rect 16764 27940 16816 27946
rect 16764 27882 16816 27888
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16592 20330 16620 20538
rect 16776 20330 16804 27882
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16776 19310 16804 20266
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16868 18970 16896 19790
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 17052 18834 17080 19110
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17236 18426 17264 18634
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17328 17338 17356 29514
rect 17512 29034 17540 31418
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17420 25430 17448 26386
rect 17500 26240 17552 26246
rect 17500 26182 17552 26188
rect 17408 25424 17460 25430
rect 17408 25366 17460 25372
rect 17512 25362 17540 26182
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17512 24274 17540 25298
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17512 23186 17540 24210
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 17696 19242 17724 31214
rect 17972 30938 18000 31418
rect 18248 30938 18276 31690
rect 18340 31278 18368 33254
rect 18432 33046 18460 34002
rect 18984 33590 19012 34138
rect 19904 33862 19932 34478
rect 19892 33856 19944 33862
rect 19892 33798 19944 33804
rect 18972 33584 19024 33590
rect 18972 33526 19024 33532
rect 19260 33522 19380 33538
rect 19248 33516 19392 33522
rect 19300 33510 19340 33516
rect 19248 33458 19300 33464
rect 19340 33458 19392 33464
rect 19904 33454 19932 33798
rect 19892 33448 19944 33454
rect 19892 33390 19944 33396
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 18420 33040 18472 33046
rect 18420 32982 18472 32988
rect 18524 32366 18552 33254
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19628 32502 19656 32914
rect 19616 32496 19668 32502
rect 19616 32438 19668 32444
rect 19996 32366 20024 33254
rect 18512 32360 18564 32366
rect 18512 32302 18564 32308
rect 19984 32360 20036 32366
rect 19984 32302 20036 32308
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19996 31890 20024 32302
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19432 31680 19484 31686
rect 19432 31622 19484 31628
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18328 31136 18380 31142
rect 18328 31078 18380 31084
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 18236 30932 18288 30938
rect 18236 30874 18288 30880
rect 17972 29850 18000 30874
rect 18248 29850 18276 30874
rect 17960 29844 18012 29850
rect 17960 29786 18012 29792
rect 18236 29844 18288 29850
rect 18236 29786 18288 29792
rect 18340 29782 18368 31078
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 17868 28620 17920 28626
rect 17868 28562 17920 28568
rect 17880 28218 17908 28562
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17880 28082 17908 28154
rect 17868 28076 17920 28082
rect 17868 28018 17920 28024
rect 17880 27674 17908 28018
rect 18144 27940 18196 27946
rect 18144 27882 18196 27888
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17880 26382 17908 27610
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17880 22778 17908 22918
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17880 22574 17908 22714
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17880 22030 17908 22510
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21894 17908 21966
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17880 20534 17908 21830
rect 17972 21690 18000 21898
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 20058 18000 20334
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 17746 18000 18090
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 14074 12664 14214
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12544 12374 12572 13806
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11440 10674 11468 12242
rect 12636 10810 12664 14010
rect 13004 13938 13032 14350
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 14752 13870 14780 14486
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14844 12782 14872 16934
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15028 13870 15056 14758
rect 15212 14006 15240 17070
rect 18064 14550 18092 24142
rect 18156 23050 18184 27882
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 18340 22386 18368 29718
rect 18418 26208 18474 26217
rect 18418 26143 18474 26152
rect 18432 26042 18460 26143
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18432 24886 18460 25978
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18432 24410 18460 24686
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18156 22358 18368 22386
rect 18156 21026 18184 22358
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18248 21146 18276 21830
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 18156 20998 18276 21026
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 18834 18184 20198
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18248 17746 18276 20998
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18248 17542 18276 17682
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18524 16658 18552 30194
rect 19248 29844 19300 29850
rect 19248 29786 19300 29792
rect 19260 29646 19288 29786
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 18696 29504 18748 29510
rect 18696 29446 18748 29452
rect 18604 27056 18656 27062
rect 18604 26998 18656 27004
rect 18616 25838 18644 26998
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18616 22098 18644 24550
rect 18708 22574 18736 29446
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 19352 28762 19380 29038
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19352 27470 19380 27950
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19352 26518 19380 27406
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19444 26382 19472 31622
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19996 30802 20024 31826
rect 19984 30796 20036 30802
rect 19984 30738 20036 30744
rect 19892 30592 19944 30598
rect 19892 30534 19944 30540
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19904 28914 19932 30534
rect 19996 30190 20024 30738
rect 20088 30326 20116 37606
rect 20824 37330 20852 38422
rect 21732 38344 21784 38350
rect 21732 38286 21784 38292
rect 21744 37942 21772 38286
rect 22204 38010 22232 39034
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 21732 37936 21784 37942
rect 21732 37878 21784 37884
rect 22204 37806 22232 37946
rect 22652 37936 22704 37942
rect 22650 37904 22652 37913
rect 22704 37904 22706 37913
rect 22650 37839 22706 37848
rect 21364 37800 21416 37806
rect 21364 37742 21416 37748
rect 22192 37800 22244 37806
rect 22192 37742 22244 37748
rect 21376 37670 21404 37742
rect 21364 37664 21416 37670
rect 21364 37606 21416 37612
rect 22204 37398 22232 37742
rect 22756 37398 22784 39578
rect 23664 38888 23716 38894
rect 23664 38830 23716 38836
rect 23676 38486 23704 38830
rect 23768 38554 23796 40870
rect 23756 38548 23808 38554
rect 23756 38490 23808 38496
rect 23664 38480 23716 38486
rect 23664 38422 23716 38428
rect 23860 38282 23888 44678
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 43382 24808 44338
rect 27816 44334 27844 45970
rect 27804 44328 27856 44334
rect 27804 44270 27856 44276
rect 27816 43858 27844 44270
rect 28264 44260 28316 44266
rect 28264 44202 28316 44208
rect 29000 44260 29052 44266
rect 29000 44202 29052 44208
rect 28276 43858 28304 44202
rect 27804 43852 27856 43858
rect 27804 43794 27856 43800
rect 28264 43852 28316 43858
rect 28264 43794 28316 43800
rect 28632 43852 28684 43858
rect 28632 43794 28684 43800
rect 28644 43654 28672 43794
rect 29012 43790 29040 44202
rect 29104 44198 29132 45970
rect 29196 45898 29224 46446
rect 30852 46374 30880 46514
rect 31036 46374 31064 46854
rect 31944 46504 31996 46510
rect 31944 46446 31996 46452
rect 32036 46504 32088 46510
rect 32036 46446 32088 46452
rect 30840 46368 30892 46374
rect 30840 46310 30892 46316
rect 31024 46368 31076 46374
rect 31024 46310 31076 46316
rect 29184 45892 29236 45898
rect 29184 45834 29236 45840
rect 29196 45082 29224 45834
rect 30380 45824 30432 45830
rect 30380 45766 30432 45772
rect 30392 45354 30420 45766
rect 30852 45490 30880 46310
rect 30840 45484 30892 45490
rect 30840 45426 30892 45432
rect 30380 45348 30432 45354
rect 30380 45290 30432 45296
rect 30852 45286 30880 45426
rect 31852 45416 31904 45422
rect 31852 45358 31904 45364
rect 30840 45280 30892 45286
rect 30840 45222 30892 45228
rect 29184 45076 29236 45082
rect 29184 45018 29236 45024
rect 29184 44940 29236 44946
rect 29184 44882 29236 44888
rect 29092 44192 29144 44198
rect 29092 44134 29144 44140
rect 29196 43926 29224 44882
rect 29184 43920 29236 43926
rect 29184 43862 29236 43868
rect 29000 43784 29052 43790
rect 29000 43726 29052 43732
rect 28632 43648 28684 43654
rect 28632 43590 28684 43596
rect 28644 43450 28672 43590
rect 28632 43444 28684 43450
rect 28632 43386 28684 43392
rect 24768 43376 24820 43382
rect 24768 43318 24820 43324
rect 24124 43308 24176 43314
rect 24124 43250 24176 43256
rect 24136 41070 24164 43250
rect 26240 43240 26292 43246
rect 26240 43182 26292 43188
rect 25044 43104 25096 43110
rect 25044 43046 25096 43052
rect 24124 41064 24176 41070
rect 24124 41006 24176 41012
rect 24676 41064 24728 41070
rect 24676 41006 24728 41012
rect 24688 40390 24716 41006
rect 24676 40384 24728 40390
rect 24676 40326 24728 40332
rect 24124 39840 24176 39846
rect 24124 39782 24176 39788
rect 24136 39642 24164 39782
rect 24124 39636 24176 39642
rect 24124 39578 24176 39584
rect 23848 38276 23900 38282
rect 23848 38218 23900 38224
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 22192 37392 22244 37398
rect 22744 37392 22796 37398
rect 22244 37340 22416 37346
rect 22192 37334 22416 37340
rect 22744 37334 22796 37340
rect 22204 37330 22416 37334
rect 20812 37324 20864 37330
rect 20812 37266 20864 37272
rect 21456 37324 21508 37330
rect 22204 37324 22428 37330
rect 22204 37318 22376 37324
rect 21456 37266 21508 37272
rect 22376 37266 22428 37272
rect 21468 36718 21496 37266
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 21836 36718 21864 37198
rect 21456 36712 21508 36718
rect 21456 36654 21508 36660
rect 21824 36712 21876 36718
rect 21876 36660 21956 36666
rect 21824 36654 21956 36660
rect 21468 36242 21496 36654
rect 21836 36638 21956 36654
rect 21928 36242 21956 36638
rect 21456 36236 21508 36242
rect 21456 36178 21508 36184
rect 21916 36236 21968 36242
rect 21916 36178 21968 36184
rect 22284 36236 22336 36242
rect 22284 36178 22336 36184
rect 21928 35834 21956 36178
rect 22296 36038 22324 36178
rect 22284 36032 22336 36038
rect 22284 35974 22336 35980
rect 20628 35828 20680 35834
rect 20628 35770 20680 35776
rect 21916 35828 21968 35834
rect 21916 35770 21968 35776
rect 20640 35494 20668 35770
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 20536 35488 20588 35494
rect 20536 35430 20588 35436
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 20548 34950 20576 35430
rect 20536 34944 20588 34950
rect 20536 34886 20588 34892
rect 20548 34542 20576 34886
rect 20536 34536 20588 34542
rect 20536 34478 20588 34484
rect 20640 32842 20668 35430
rect 21100 35290 21128 35634
rect 21364 35624 21416 35630
rect 21364 35566 21416 35572
rect 21376 35290 21404 35566
rect 21088 35284 21140 35290
rect 21088 35226 21140 35232
rect 21364 35284 21416 35290
rect 21364 35226 21416 35232
rect 21100 34678 21128 35226
rect 21376 35154 21404 35226
rect 21364 35148 21416 35154
rect 21364 35090 21416 35096
rect 21088 34672 21140 34678
rect 21088 34614 21140 34620
rect 21100 34542 21128 34614
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21376 34066 21404 35090
rect 21836 34746 21864 35634
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21928 34762 21956 34886
rect 21928 34746 22048 34762
rect 21824 34740 21876 34746
rect 21928 34740 22060 34746
rect 21928 34734 22008 34740
rect 21824 34682 21876 34688
rect 22008 34682 22060 34688
rect 21364 34060 21416 34066
rect 21364 34002 21416 34008
rect 21376 33454 21404 34002
rect 21914 33960 21970 33969
rect 21914 33895 21916 33904
rect 21968 33895 21970 33904
rect 21916 33866 21968 33872
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22756 33561 22784 33594
rect 22742 33552 22798 33561
rect 22742 33487 22798 33496
rect 21364 33448 21416 33454
rect 21364 33390 21416 33396
rect 20628 32836 20680 32842
rect 20628 32778 20680 32784
rect 21376 32502 21404 33390
rect 21548 32972 21600 32978
rect 21548 32914 21600 32920
rect 21560 32502 21588 32914
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21730 32328 21786 32337
rect 21730 32263 21732 32272
rect 21784 32263 21786 32272
rect 21732 32234 21784 32240
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 20076 30320 20128 30326
rect 20076 30262 20128 30268
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 19996 29714 20024 29990
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 20258 29472 20314 29481
rect 20258 29407 20314 29416
rect 19904 28886 20024 28914
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19996 28014 20024 28886
rect 20272 28218 20300 29407
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20444 29028 20496 29034
rect 20732 29016 20760 29106
rect 20496 28988 20760 29016
rect 20444 28970 20496 28976
rect 20260 28212 20312 28218
rect 20260 28154 20312 28160
rect 20272 28082 20300 28154
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19892 27940 19944 27946
rect 19892 27882 19944 27888
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 18800 26042 18828 26318
rect 18788 26036 18840 26042
rect 18788 25978 18840 25984
rect 18972 25832 19024 25838
rect 18972 25774 19024 25780
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18800 24206 18828 24686
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18984 23662 19012 25774
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19076 24886 19104 25298
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19064 24880 19116 24886
rect 19064 24822 19116 24828
rect 19352 23730 19380 25094
rect 19444 24342 19472 25230
rect 19616 25152 19668 25158
rect 19616 25094 19668 25100
rect 19628 24818 19656 25094
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19432 24336 19484 24342
rect 19432 24278 19484 24284
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18788 23520 18840 23526
rect 18786 23488 18788 23497
rect 18840 23488 18842 23497
rect 18786 23423 18842 23432
rect 18984 22658 19012 23598
rect 18984 22630 19104 22658
rect 19076 22574 19104 22630
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18972 22568 19024 22574
rect 18972 22510 19024 22516
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18984 22438 19012 22510
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18616 22003 18644 22034
rect 18984 20777 19012 22374
rect 19076 22234 19104 22510
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 19168 21962 19196 22034
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 18970 20768 19026 20777
rect 18970 20703 19026 20712
rect 18984 18902 19012 20703
rect 19168 19417 19196 21898
rect 19154 19408 19210 19417
rect 19154 19343 19210 19352
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18222 18828 18702
rect 19168 18630 19196 19343
rect 19444 18834 19472 24142
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 19352 17814 19380 18702
rect 19444 18222 19472 18770
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18340 15434 18368 16594
rect 18616 15502 18644 17614
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19444 17202 19472 17546
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19904 16538 19932 27882
rect 20168 27328 20220 27334
rect 19812 16510 19932 16538
rect 20088 27288 20168 27316
rect 19812 15994 19840 16510
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19904 16114 19932 16390
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19812 15966 19932 15994
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 12986 15240 13806
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15764 13190 15792 13670
rect 16684 13462 16712 14350
rect 18064 13530 18092 14486
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12986 15792 13126
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15764 12782 15792 12922
rect 17972 12918 18000 13262
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11762 13768 12174
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11286 12756 11630
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 12636 10266 12664 10746
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12636 8634 12664 10202
rect 13004 10130 13032 10474
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13740 9586 13768 11698
rect 13832 11354 13860 11834
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 15396 11218 15424 12718
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 11762 17540 12174
rect 17972 11830 18000 12854
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 19168 11694 19196 11766
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 17052 11150 17080 11494
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 14752 11014 14780 11086
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10606 14780 10950
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14108 10266 14136 10542
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14016 8634 14044 9454
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11072 7954 11100 8434
rect 12636 8430 12664 8570
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 15212 7546 15240 11018
rect 16132 10674 16160 11018
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 9722 15332 10474
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 17052 9518 17080 11086
rect 18524 11082 18552 11630
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 9586 18552 11018
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17788 9042 17816 9522
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 9042 18092 9386
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 19076 8634 19104 9454
rect 19352 8974 19380 9862
rect 19904 9654 19932 15966
rect 20088 12238 20116 27288
rect 20168 27270 20220 27276
rect 20456 20058 20484 28970
rect 20824 28966 20852 29990
rect 20916 29238 20944 29990
rect 20904 29232 20956 29238
rect 20904 29174 20956 29180
rect 20904 29028 20956 29034
rect 20904 28970 20956 28976
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20824 28014 20852 28902
rect 20916 28762 20944 28970
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 20812 28008 20864 28014
rect 20812 27950 20864 27956
rect 20824 27538 20852 27950
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 21008 25362 21036 32166
rect 21364 31748 21416 31754
rect 21364 31690 21416 31696
rect 21180 28212 21232 28218
rect 21180 28154 21232 28160
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 21192 22030 21220 28154
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21376 21690 21404 31690
rect 22296 30122 22324 32166
rect 23676 31414 23704 37810
rect 23756 37732 23808 37738
rect 23860 37720 23888 38218
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 23808 37692 23888 37720
rect 23756 37674 23808 37680
rect 23768 32842 23796 37674
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 24504 36174 24532 36314
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 24688 33590 24716 38150
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 24780 35562 24808 36518
rect 24768 35556 24820 35562
rect 24768 35498 24820 35504
rect 24676 33584 24728 33590
rect 24676 33526 24728 33532
rect 24688 33386 24716 33526
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 24124 33380 24176 33386
rect 24124 33322 24176 33328
rect 24676 33380 24728 33386
rect 24676 33322 24728 33328
rect 23756 32836 23808 32842
rect 23756 32778 23808 32784
rect 23664 31408 23716 31414
rect 22742 31376 22798 31385
rect 23664 31350 23716 31356
rect 22742 31311 22744 31320
rect 22796 31311 22798 31320
rect 22744 31282 22796 31288
rect 22742 31240 22798 31249
rect 22742 31175 22744 31184
rect 22796 31175 22798 31184
rect 24032 31204 24084 31210
rect 22744 31146 22796 31152
rect 24032 31146 24084 31152
rect 24044 30802 24072 31146
rect 24032 30796 24084 30802
rect 24032 30738 24084 30744
rect 24136 30682 24164 33322
rect 24872 33046 24900 33390
rect 24860 33040 24912 33046
rect 24860 32982 24912 32988
rect 24308 32768 24360 32774
rect 24308 32710 24360 32716
rect 24044 30654 24164 30682
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22284 30116 22336 30122
rect 22284 30058 22336 30064
rect 22480 30054 22508 30194
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 23296 30048 23348 30054
rect 23296 29990 23348 29996
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23018 29336 23074 29345
rect 23018 29271 23020 29280
rect 23072 29271 23074 29280
rect 23112 29300 23164 29306
rect 23020 29242 23072 29248
rect 23112 29242 23164 29248
rect 22836 26512 22888 26518
rect 22836 26454 22888 26460
rect 22376 26444 22428 26450
rect 22376 26386 22428 26392
rect 22388 25498 22416 26386
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22388 25362 22416 25434
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 21548 24880 21600 24886
rect 21548 24822 21600 24828
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21376 20058 21404 21626
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 18034 20208 19654
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20272 18426 20300 18702
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20180 18006 20300 18034
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20180 16794 20208 17818
rect 20272 17542 20300 18006
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20272 12442 20300 17478
rect 20824 17066 20852 17478
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20824 16697 20852 17002
rect 20810 16688 20866 16697
rect 21008 16658 21036 18158
rect 20810 16623 20866 16632
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 21008 15706 21036 16594
rect 21560 16250 21588 24822
rect 21744 21486 21772 25230
rect 22480 24342 22508 25230
rect 22756 24750 22784 26318
rect 22848 25362 22876 26454
rect 23124 25498 23152 29242
rect 23308 28966 23336 29990
rect 23676 29782 23704 29990
rect 23664 29776 23716 29782
rect 23664 29718 23716 29724
rect 24044 29646 24072 30654
rect 24124 30592 24176 30598
rect 24124 30534 24176 30540
rect 24136 29714 24164 30534
rect 24124 29708 24176 29714
rect 24124 29650 24176 29656
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 24214 29200 24270 29209
rect 24214 29135 24270 29144
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23940 28960 23992 28966
rect 23940 28902 23992 28908
rect 23308 26518 23336 28902
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23296 26512 23348 26518
rect 23296 26454 23348 26460
rect 23400 26450 23428 27474
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22468 24336 22520 24342
rect 22468 24278 22520 24284
rect 22480 23322 22508 24278
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22296 20058 22324 20878
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22388 19922 22416 20198
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22020 19174 22048 19858
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22020 18902 22048 19110
rect 22008 18896 22060 18902
rect 22008 18838 22060 18844
rect 22848 18766 22876 25298
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23216 24274 23244 24550
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23492 22574 23520 27406
rect 23676 26926 23704 28494
rect 23952 27130 23980 28902
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23664 26920 23716 26926
rect 23664 26862 23716 26868
rect 24228 26078 24256 29135
rect 23768 26050 24256 26078
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 23676 21078 23704 22170
rect 23664 21072 23716 21078
rect 23492 21032 23664 21060
rect 23492 20398 23520 21032
rect 23664 21014 23716 21020
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23676 20262 23704 20334
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23584 18970 23612 19110
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21652 16794 21680 16934
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21270 16008 21326 16017
rect 21270 15943 21272 15952
rect 21324 15943 21326 15952
rect 21272 15914 21324 15920
rect 21284 15706 21312 15914
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21560 14618 21588 16186
rect 21652 15910 21680 16730
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20640 14074 20668 14418
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20640 12306 20668 14010
rect 21008 13870 21036 14214
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 11898 20116 12174
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 21008 11762 21036 13806
rect 21652 13530 21680 15846
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21652 13326 21680 13466
rect 22296 13394 22324 13670
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 22848 12442 22876 16594
rect 23676 16250 23704 20198
rect 23768 18970 23796 26050
rect 24320 25498 24348 32710
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 24952 31272 25004 31278
rect 25056 31260 25084 43046
rect 26252 42362 26280 43182
rect 27528 43104 27580 43110
rect 27528 43046 27580 43052
rect 27540 42362 27568 43046
rect 26240 42356 26292 42362
rect 26240 42298 26292 42304
rect 27528 42356 27580 42362
rect 27528 42298 27580 42304
rect 29196 42294 29224 43862
rect 29920 42764 29972 42770
rect 29920 42706 29972 42712
rect 29184 42288 29236 42294
rect 28998 42256 29054 42265
rect 27344 42220 27396 42226
rect 29184 42230 29236 42236
rect 28998 42191 29000 42200
rect 27344 42162 27396 42168
rect 29052 42191 29054 42200
rect 29000 42162 29052 42168
rect 25136 42152 25188 42158
rect 25136 42094 25188 42100
rect 25148 41818 25176 42094
rect 26516 42016 26568 42022
rect 26516 41958 26568 41964
rect 25136 41812 25188 41818
rect 25136 41754 25188 41760
rect 26528 41682 26556 41958
rect 27356 41818 27384 42162
rect 29644 42084 29696 42090
rect 29644 42026 29696 42032
rect 29276 42016 29328 42022
rect 29276 41958 29328 41964
rect 27344 41812 27396 41818
rect 27344 41754 27396 41760
rect 26516 41676 26568 41682
rect 26516 41618 26568 41624
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26516 41132 26568 41138
rect 26516 41074 26568 41080
rect 26148 41064 26200 41070
rect 26148 41006 26200 41012
rect 26160 40934 26188 41006
rect 26148 40928 26200 40934
rect 26148 40870 26200 40876
rect 26528 40769 26556 41074
rect 26514 40760 26570 40769
rect 26514 40695 26570 40704
rect 26240 38480 26292 38486
rect 26240 38422 26292 38428
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25516 37874 25544 38150
rect 25504 37868 25556 37874
rect 25504 37810 25556 37816
rect 25596 37868 25648 37874
rect 25596 37810 25648 37816
rect 25504 36848 25556 36854
rect 25608 36836 25636 37810
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 26160 37670 26188 37742
rect 26148 37664 26200 37670
rect 26148 37606 26200 37612
rect 26252 36854 26280 38422
rect 25556 36808 25636 36836
rect 26240 36848 26292 36854
rect 25504 36790 25556 36796
rect 26240 36790 26292 36796
rect 26332 36848 26384 36854
rect 26384 36808 26464 36836
rect 26332 36790 26384 36796
rect 26056 36644 26108 36650
rect 26056 36586 26108 36592
rect 26332 36644 26384 36650
rect 26332 36586 26384 36592
rect 25872 36576 25924 36582
rect 25872 36518 25924 36524
rect 25884 36038 25912 36518
rect 25504 36032 25556 36038
rect 25504 35974 25556 35980
rect 25872 36032 25924 36038
rect 25872 35974 25924 35980
rect 25412 34060 25464 34066
rect 25412 34002 25464 34008
rect 25320 33040 25372 33046
rect 25320 32982 25372 32988
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25240 32434 25268 32846
rect 25228 32428 25280 32434
rect 25228 32370 25280 32376
rect 25004 31232 25084 31260
rect 24952 31214 25004 31220
rect 24688 30258 24716 31214
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 24964 30190 24992 31078
rect 24768 30184 24820 30190
rect 24768 30126 24820 30132
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24584 29572 24636 29578
rect 24584 29514 24636 29520
rect 24596 29238 24624 29514
rect 24780 29510 24808 30126
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 25044 29232 25096 29238
rect 25044 29174 25096 29180
rect 25056 29102 25084 29174
rect 25044 29096 25096 29102
rect 25136 29096 25188 29102
rect 25044 29038 25096 29044
rect 25134 29064 25136 29073
rect 25188 29064 25190 29073
rect 25134 28999 25190 29008
rect 25240 28422 25268 32370
rect 25332 30938 25360 32982
rect 25424 31822 25452 34002
rect 25412 31816 25464 31822
rect 25412 31758 25464 31764
rect 25516 31414 25544 35974
rect 26068 35834 26096 36586
rect 26344 36242 26372 36586
rect 26332 36236 26384 36242
rect 26332 36178 26384 36184
rect 26436 36038 26464 36808
rect 26620 36718 26648 41414
rect 27356 40730 27384 41754
rect 27712 41540 27764 41546
rect 27712 41482 27764 41488
rect 27724 41274 27752 41482
rect 27988 41472 28040 41478
rect 27988 41414 28040 41420
rect 27712 41268 27764 41274
rect 27712 41210 27764 41216
rect 28000 41070 28028 41414
rect 27988 41064 28040 41070
rect 27988 41006 28040 41012
rect 27896 40928 27948 40934
rect 27434 40896 27490 40905
rect 27896 40870 27948 40876
rect 27434 40831 27490 40840
rect 27448 40730 27476 40831
rect 27344 40724 27396 40730
rect 27344 40666 27396 40672
rect 27436 40724 27488 40730
rect 27436 40666 27488 40672
rect 26976 40656 27028 40662
rect 26976 40598 27028 40604
rect 26700 39364 26752 39370
rect 26700 39306 26752 39312
rect 26712 39030 26740 39306
rect 26700 39024 26752 39030
rect 26700 38966 26752 38972
rect 26712 38418 26740 38966
rect 26700 38412 26752 38418
rect 26700 38354 26752 38360
rect 26988 37482 27016 40598
rect 27252 40588 27304 40594
rect 27356 40576 27384 40666
rect 27304 40548 27384 40576
rect 27252 40530 27304 40536
rect 27710 40352 27766 40361
rect 27710 40287 27766 40296
rect 27356 40186 27568 40202
rect 27724 40186 27752 40287
rect 27344 40180 27580 40186
rect 27396 40174 27528 40180
rect 27344 40122 27396 40128
rect 27528 40122 27580 40128
rect 27712 40180 27764 40186
rect 27712 40122 27764 40128
rect 27908 39506 27936 40870
rect 28000 40526 28028 41006
rect 29184 40928 29236 40934
rect 29184 40870 29236 40876
rect 29000 40656 29052 40662
rect 29000 40598 29052 40604
rect 29090 40624 29146 40633
rect 27988 40520 28040 40526
rect 27988 40462 28040 40468
rect 29012 40390 29040 40598
rect 29090 40559 29146 40568
rect 29104 40526 29132 40559
rect 29196 40526 29224 40870
rect 29092 40520 29144 40526
rect 29092 40462 29144 40468
rect 29184 40520 29236 40526
rect 29184 40462 29236 40468
rect 29196 40390 29224 40462
rect 29000 40384 29052 40390
rect 29184 40384 29236 40390
rect 29000 40326 29052 40332
rect 29182 40352 29184 40361
rect 29236 40352 29238 40361
rect 29182 40287 29238 40296
rect 28448 39976 28500 39982
rect 28448 39918 28500 39924
rect 27896 39500 27948 39506
rect 27896 39442 27948 39448
rect 27620 37936 27672 37942
rect 27672 37896 27752 37924
rect 27620 37878 27672 37884
rect 27724 37806 27752 37896
rect 27712 37800 27764 37806
rect 27712 37742 27764 37748
rect 27160 37732 27212 37738
rect 27160 37674 27212 37680
rect 26896 37454 27016 37482
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 26516 36236 26568 36242
rect 26516 36178 26568 36184
rect 26424 36032 26476 36038
rect 26424 35974 26476 35980
rect 26056 35828 26108 35834
rect 26056 35770 26108 35776
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 26240 35556 26292 35562
rect 26240 35498 26292 35504
rect 25608 34610 26004 34626
rect 25596 34604 26016 34610
rect 25648 34598 25964 34604
rect 25596 34546 25648 34552
rect 25964 34546 26016 34552
rect 25688 34536 25740 34542
rect 25686 34504 25688 34513
rect 26148 34536 26200 34542
rect 25740 34504 25742 34513
rect 25686 34439 25742 34448
rect 25792 34484 26148 34490
rect 25792 34478 26200 34484
rect 25792 34462 26188 34478
rect 25792 34406 25820 34462
rect 25780 34400 25832 34406
rect 26252 34388 26280 35498
rect 25780 34342 25832 34348
rect 26068 34360 26280 34388
rect 26068 33998 26096 34360
rect 26344 34066 26372 35566
rect 26528 35222 26556 36178
rect 26700 35828 26752 35834
rect 26700 35770 26752 35776
rect 26608 35624 26660 35630
rect 26608 35566 26660 35572
rect 26516 35216 26568 35222
rect 26516 35158 26568 35164
rect 26620 35154 26648 35566
rect 26608 35148 26660 35154
rect 26608 35090 26660 35096
rect 26712 35086 26740 35770
rect 26700 35080 26752 35086
rect 26700 35022 26752 35028
rect 26804 34513 26832 37198
rect 26896 36310 26924 37454
rect 27172 37330 27200 37674
rect 27160 37324 27212 37330
rect 27160 37266 27212 37272
rect 27908 37262 27936 39442
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 28276 38486 28304 39374
rect 28460 39098 28488 39918
rect 28448 39092 28500 39098
rect 28448 39034 28500 39040
rect 28460 38894 28488 39034
rect 28448 38888 28500 38894
rect 28448 38830 28500 38836
rect 28264 38480 28316 38486
rect 28264 38422 28316 38428
rect 27896 37256 27948 37262
rect 27896 37198 27948 37204
rect 26884 36304 26936 36310
rect 26884 36246 26936 36252
rect 27620 35760 27672 35766
rect 26896 35686 27292 35714
rect 27620 35702 27672 35708
rect 26896 35630 26924 35686
rect 26884 35624 26936 35630
rect 26884 35566 26936 35572
rect 27068 35624 27120 35630
rect 27068 35566 27120 35572
rect 27080 35494 27108 35566
rect 27264 35562 27292 35686
rect 27252 35556 27304 35562
rect 27252 35498 27304 35504
rect 27068 35488 27120 35494
rect 27068 35430 27120 35436
rect 27160 35488 27212 35494
rect 27160 35430 27212 35436
rect 26884 35216 26936 35222
rect 26884 35158 26936 35164
rect 26896 35018 26924 35158
rect 27172 35154 27200 35430
rect 27160 35148 27212 35154
rect 27160 35090 27212 35096
rect 27252 35080 27304 35086
rect 27252 35022 27304 35028
rect 27436 35080 27488 35086
rect 27436 35022 27488 35028
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26790 34504 26846 34513
rect 26790 34439 26846 34448
rect 27068 34128 27120 34134
rect 27066 34096 27068 34105
rect 27120 34096 27122 34105
rect 26332 34060 26384 34066
rect 27264 34082 27292 35022
rect 27448 34746 27476 35022
rect 27632 34746 27660 35702
rect 28080 35488 28132 35494
rect 28080 35430 28132 35436
rect 28092 35154 28120 35430
rect 28080 35148 28132 35154
rect 28080 35090 28132 35096
rect 28092 35018 28120 35090
rect 28080 35012 28132 35018
rect 28080 34954 28132 34960
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 27620 34740 27672 34746
rect 27620 34682 27672 34688
rect 27264 34066 27384 34082
rect 27066 34031 27122 34040
rect 27160 34060 27212 34066
rect 26332 34002 26384 34008
rect 27160 34002 27212 34008
rect 27264 34060 27396 34066
rect 27264 34054 27344 34060
rect 26056 33992 26108 33998
rect 26240 33992 26292 33998
rect 26056 33934 26108 33940
rect 26160 33940 26240 33946
rect 26160 33934 26292 33940
rect 26068 33590 26096 33934
rect 26160 33918 26280 33934
rect 26056 33584 26108 33590
rect 26056 33526 26108 33532
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 25596 32496 25648 32502
rect 25596 32438 25648 32444
rect 25608 32366 25636 32438
rect 26068 32434 26096 33390
rect 26160 32910 26188 33918
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26344 32366 26372 34002
rect 27172 32502 27200 34002
rect 27264 33318 27292 34054
rect 27344 34002 27396 34008
rect 27448 33538 27476 34682
rect 27712 34672 27764 34678
rect 27712 34614 27764 34620
rect 27526 34504 27582 34513
rect 27526 34439 27582 34448
rect 27540 34406 27568 34439
rect 27528 34400 27580 34406
rect 27528 34342 27580 34348
rect 27620 34128 27672 34134
rect 27618 34096 27620 34105
rect 27672 34096 27674 34105
rect 27618 34031 27674 34040
rect 27724 33862 27752 34614
rect 29288 34066 29316 41958
rect 29656 41818 29684 42026
rect 29932 41818 29960 42706
rect 30852 42634 30880 45222
rect 31864 44334 31892 45358
rect 31956 44554 31984 46446
rect 32048 46102 32076 46446
rect 32128 46368 32180 46374
rect 32128 46310 32180 46316
rect 32312 46368 32364 46374
rect 32312 46310 32364 46316
rect 32140 46170 32168 46310
rect 32128 46164 32180 46170
rect 32128 46106 32180 46112
rect 32036 46096 32088 46102
rect 32036 46038 32088 46044
rect 32324 46034 32352 46310
rect 32312 46028 32364 46034
rect 32312 45970 32364 45976
rect 32600 45966 32628 46990
rect 32588 45960 32640 45966
rect 32588 45902 32640 45908
rect 32876 45490 32904 46990
rect 38752 46980 38804 46986
rect 38752 46922 38804 46928
rect 33784 46912 33836 46918
rect 33784 46854 33836 46860
rect 33796 46510 33824 46854
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 38764 46510 38792 46922
rect 40040 46912 40092 46918
rect 40040 46854 40092 46860
rect 33784 46504 33836 46510
rect 33784 46446 33836 46452
rect 34428 46504 34480 46510
rect 34428 46446 34480 46452
rect 38752 46504 38804 46510
rect 38752 46446 38804 46452
rect 33876 46368 33928 46374
rect 33876 46310 33928 46316
rect 32864 45484 32916 45490
rect 32864 45426 32916 45432
rect 33888 45286 33916 46310
rect 34440 46170 34468 46446
rect 34980 46368 35032 46374
rect 34980 46310 35032 46316
rect 38476 46368 38528 46374
rect 38476 46310 38528 46316
rect 34428 46164 34480 46170
rect 34428 46106 34480 46112
rect 34992 45898 35020 46310
rect 38488 46034 38516 46310
rect 38476 46028 38528 46034
rect 38476 45970 38528 45976
rect 35440 45960 35492 45966
rect 35440 45902 35492 45908
rect 34980 45892 35032 45898
rect 34980 45834 35032 45840
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 33876 45280 33928 45286
rect 33876 45222 33928 45228
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 31956 44526 32076 44554
rect 31944 44396 31996 44402
rect 31944 44338 31996 44344
rect 31852 44328 31904 44334
rect 31852 44270 31904 44276
rect 31956 43994 31984 44338
rect 31944 43988 31996 43994
rect 31944 43930 31996 43936
rect 32048 43926 32076 44526
rect 32864 44328 32916 44334
rect 32864 44270 32916 44276
rect 32036 43920 32088 43926
rect 32036 43862 32088 43868
rect 30840 42628 30892 42634
rect 30840 42570 30892 42576
rect 32048 42294 32076 43862
rect 32770 43344 32826 43353
rect 32770 43279 32772 43288
rect 32824 43279 32826 43288
rect 32772 43250 32824 43256
rect 32312 43104 32364 43110
rect 32312 43046 32364 43052
rect 32324 42906 32352 43046
rect 32312 42900 32364 42906
rect 32312 42842 32364 42848
rect 32324 42770 32352 42842
rect 32876 42770 32904 44270
rect 32956 43988 33008 43994
rect 32956 43930 33008 43936
rect 34244 43988 34296 43994
rect 34244 43930 34296 43936
rect 32968 43858 32996 43930
rect 32956 43852 33008 43858
rect 32956 43794 33008 43800
rect 32968 43246 32996 43794
rect 34256 43654 34284 43930
rect 35452 43654 35480 45902
rect 38568 45620 38620 45626
rect 38568 45562 38620 45568
rect 36360 43852 36412 43858
rect 36360 43794 36412 43800
rect 38476 43852 38528 43858
rect 38476 43794 38528 43800
rect 34244 43648 34296 43654
rect 34244 43590 34296 43596
rect 35440 43648 35492 43654
rect 35440 43590 35492 43596
rect 33324 43444 33376 43450
rect 33324 43386 33376 43392
rect 33336 43246 33364 43386
rect 32956 43240 33008 43246
rect 32956 43182 33008 43188
rect 33324 43240 33376 43246
rect 33324 43182 33376 43188
rect 33968 43104 34020 43110
rect 33968 43046 34020 43052
rect 33980 42906 34008 43046
rect 33968 42900 34020 42906
rect 33968 42842 34020 42848
rect 34256 42770 34284 43590
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 35452 43314 35480 43590
rect 35440 43308 35492 43314
rect 35440 43250 35492 43256
rect 32312 42764 32364 42770
rect 32312 42706 32364 42712
rect 32864 42764 32916 42770
rect 32864 42706 32916 42712
rect 34244 42764 34296 42770
rect 34244 42706 34296 42712
rect 32876 42566 32904 42706
rect 32864 42560 32916 42566
rect 32864 42502 32916 42508
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 31208 42288 31260 42294
rect 31208 42230 31260 42236
rect 32036 42288 32088 42294
rect 32128 42288 32180 42294
rect 32036 42230 32088 42236
rect 32126 42256 32128 42265
rect 32180 42256 32182 42265
rect 31220 42158 31248 42230
rect 32126 42191 32182 42200
rect 31208 42152 31260 42158
rect 31208 42094 31260 42100
rect 29644 41812 29696 41818
rect 29644 41754 29696 41760
rect 29920 41812 29972 41818
rect 29920 41754 29972 41760
rect 29368 41676 29420 41682
rect 29368 41618 29420 41624
rect 29380 35766 29408 41618
rect 29656 41070 29684 41754
rect 35452 41750 35480 43250
rect 35716 43240 35768 43246
rect 35716 43182 35768 43188
rect 35728 42702 35756 43182
rect 35716 42696 35768 42702
rect 35716 42638 35768 42644
rect 36268 42152 36320 42158
rect 36268 42094 36320 42100
rect 35440 41744 35492 41750
rect 35440 41686 35492 41692
rect 31760 41676 31812 41682
rect 31760 41618 31812 41624
rect 30746 41576 30802 41585
rect 30746 41511 30748 41520
rect 30800 41511 30802 41520
rect 30748 41482 30800 41488
rect 30564 41268 30616 41274
rect 30564 41210 30616 41216
rect 30576 41070 30604 41210
rect 29644 41064 29696 41070
rect 29644 41006 29696 41012
rect 30564 41064 30616 41070
rect 30564 41006 30616 41012
rect 29460 40588 29512 40594
rect 29460 40530 29512 40536
rect 29472 40186 29500 40530
rect 31772 40526 31800 41618
rect 35072 41608 35124 41614
rect 35070 41576 35072 41585
rect 35124 41576 35126 41585
rect 35070 41511 35126 41520
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 33416 40996 33468 41002
rect 33416 40938 33468 40944
rect 33428 40526 33456 40938
rect 34152 40656 34204 40662
rect 34150 40624 34152 40633
rect 34204 40624 34206 40633
rect 34150 40559 34206 40568
rect 31760 40520 31812 40526
rect 31760 40462 31812 40468
rect 32956 40520 33008 40526
rect 32956 40462 33008 40468
rect 33416 40520 33468 40526
rect 33416 40462 33468 40468
rect 32968 40390 32996 40462
rect 32956 40384 33008 40390
rect 32956 40326 33008 40332
rect 34704 40384 34756 40390
rect 34704 40326 34756 40332
rect 29460 40180 29512 40186
rect 29460 40122 29512 40128
rect 29460 39976 29512 39982
rect 29460 39918 29512 39924
rect 29472 39846 29500 39918
rect 29460 39840 29512 39846
rect 29460 39782 29512 39788
rect 32404 39840 32456 39846
rect 32404 39782 32456 39788
rect 29552 39296 29604 39302
rect 29552 39238 29604 39244
rect 29564 39098 29592 39238
rect 29552 39092 29604 39098
rect 29552 39034 29604 39040
rect 32312 37664 32364 37670
rect 32312 37606 32364 37612
rect 30380 37460 30432 37466
rect 30380 37402 30432 37408
rect 30392 36650 30420 37402
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32232 36650 32260 37062
rect 30380 36644 30432 36650
rect 30380 36586 30432 36592
rect 32220 36644 32272 36650
rect 32220 36586 32272 36592
rect 29368 35760 29420 35766
rect 29368 35702 29420 35708
rect 31942 35728 31998 35737
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 27802 33960 27858 33969
rect 27802 33895 27804 33904
rect 27856 33895 27858 33904
rect 27804 33866 27856 33872
rect 27712 33856 27764 33862
rect 27712 33798 27764 33804
rect 27448 33510 27660 33538
rect 27632 33454 27660 33510
rect 27620 33448 27672 33454
rect 27620 33390 27672 33396
rect 27712 33380 27764 33386
rect 27712 33322 27764 33328
rect 27252 33312 27304 33318
rect 27252 33254 27304 33260
rect 27528 33312 27580 33318
rect 27528 33254 27580 33260
rect 27160 32496 27212 32502
rect 27160 32438 27212 32444
rect 25596 32360 25648 32366
rect 25596 32302 25648 32308
rect 26332 32360 26384 32366
rect 26332 32302 26384 32308
rect 27068 32360 27120 32366
rect 27160 32360 27212 32366
rect 27068 32302 27120 32308
rect 27158 32328 27160 32337
rect 27212 32328 27214 32337
rect 27080 31822 27108 32302
rect 27158 32263 27214 32272
rect 27068 31816 27120 31822
rect 27068 31758 27120 31764
rect 25504 31408 25556 31414
rect 25410 31376 25466 31385
rect 25504 31350 25556 31356
rect 25410 31311 25412 31320
rect 25464 31311 25466 31320
rect 25412 31282 25464 31288
rect 25410 31240 25466 31249
rect 25410 31175 25412 31184
rect 25464 31175 25466 31184
rect 25412 31146 25464 31152
rect 25320 30932 25372 30938
rect 25320 30874 25372 30880
rect 25320 30796 25372 30802
rect 25320 30738 25372 30744
rect 25332 29238 25360 30738
rect 26792 30320 26844 30326
rect 26792 30262 26844 30268
rect 26332 30184 26384 30190
rect 26332 30126 26384 30132
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 25594 29336 25650 29345
rect 25594 29271 25650 29280
rect 25320 29232 25372 29238
rect 25320 29174 25372 29180
rect 25504 29232 25556 29238
rect 25504 29174 25556 29180
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 23940 24268 23992 24274
rect 23940 24210 23992 24216
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23860 20602 23888 22510
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23860 19922 23888 20538
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23952 17882 23980 24210
rect 24044 23254 24072 25230
rect 24136 24750 24164 25298
rect 24320 25294 24348 25434
rect 24308 25288 24360 25294
rect 24308 25230 24360 25236
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24596 24274 24624 27066
rect 24780 26450 24808 28018
rect 24964 27538 24992 28154
rect 25044 28008 25096 28014
rect 25044 27950 25096 27956
rect 25056 27606 25084 27950
rect 25044 27600 25096 27606
rect 25044 27542 25096 27548
rect 25332 27538 25360 29174
rect 25412 29096 25464 29102
rect 25410 29064 25412 29073
rect 25464 29064 25466 29073
rect 25410 28999 25466 29008
rect 24952 27532 25004 27538
rect 24952 27474 25004 27480
rect 25320 27532 25372 27538
rect 25320 27474 25372 27480
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24872 26330 24900 26726
rect 24780 26302 24900 26330
rect 24780 25498 24808 26302
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24688 24342 24716 25094
rect 24780 24954 24808 25298
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24584 24268 24636 24274
rect 24584 24210 24636 24216
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 24032 23248 24084 23254
rect 24032 23190 24084 23196
rect 24044 22574 24072 23190
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 24136 22098 24164 24074
rect 24596 24070 24624 24210
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24216 23520 24268 23526
rect 24216 23462 24268 23468
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24228 21894 24256 23462
rect 24412 23322 24440 23598
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24308 23180 24360 23186
rect 24308 23122 24360 23128
rect 24320 22506 24348 23122
rect 24308 22500 24360 22506
rect 24308 22442 24360 22448
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24228 21350 24256 21830
rect 24872 21554 24900 22374
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24216 21344 24268 21350
rect 24964 21298 24992 24550
rect 25148 24410 25176 25298
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25424 24818 25452 25094
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 25516 24614 25544 29174
rect 25608 29170 25636 29271
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25608 28014 25636 28154
rect 25596 28008 25648 28014
rect 25596 27950 25648 27956
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 25884 27334 25912 27406
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25884 27130 25912 27270
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 26160 27062 26188 29582
rect 26344 29510 26372 30126
rect 26804 29782 26832 30262
rect 27160 30184 27212 30190
rect 27160 30126 27212 30132
rect 27252 30184 27304 30190
rect 27252 30126 27304 30132
rect 27172 29850 27200 30126
rect 27264 30054 27292 30126
rect 27252 30048 27304 30054
rect 27252 29990 27304 29996
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 26792 29776 26844 29782
rect 26792 29718 26844 29724
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26240 28416 26292 28422
rect 26240 28358 26292 28364
rect 26252 27470 26280 28358
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 26252 27334 26280 27406
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 25964 25220 26016 25226
rect 25964 25162 26016 25168
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25424 21894 25452 22986
rect 25976 22574 26004 25162
rect 26160 24750 26188 26998
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 26252 22982 26280 27270
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25424 21457 25452 21830
rect 25976 21690 26004 22510
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 25410 21448 25466 21457
rect 25410 21383 25466 21392
rect 24216 21286 24268 21292
rect 24228 20806 24256 21286
rect 24872 21270 24992 21298
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24780 19258 24808 20742
rect 24872 19514 24900 21270
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24860 19304 24912 19310
rect 24780 19252 24860 19258
rect 24780 19246 24912 19252
rect 24780 19230 24900 19246
rect 24872 18222 24900 19230
rect 24964 18834 24992 19654
rect 25688 19236 25740 19242
rect 25688 19178 25740 19184
rect 25700 18970 25728 19178
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24964 18630 24992 18770
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 25148 18290 25176 18634
rect 26252 18426 26280 19858
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24872 18086 24900 18158
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24872 16794 24900 18022
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24872 16250 24900 16730
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 23676 16046 23704 16186
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 15570 24440 15846
rect 25240 15706 25268 15982
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24964 13870 24992 15506
rect 25412 15428 25464 15434
rect 25412 15370 25464 15376
rect 25424 14074 25452 15370
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24320 12986 24348 13466
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24964 12866 24992 13806
rect 24872 12838 24992 12866
rect 24872 12782 24900 12838
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 10810 20668 11562
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 9926 20484 10406
rect 20916 10266 20944 10542
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21652 10130 21680 11494
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19444 9110 19472 9590
rect 21284 9586 21312 10066
rect 22848 10062 22876 12378
rect 25056 11898 25084 12718
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25884 11762 25912 12582
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 25608 9926 25636 10406
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 22204 8974 22232 9318
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 22204 8430 22232 8910
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 22296 8430 22324 8774
rect 23952 8498 23980 8774
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 25608 8430 25636 9862
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12084 6866 12112 7210
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6866 12572 7142
rect 13924 6934 13952 7278
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12084 4826 12112 6802
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 25608 5302 25636 8366
rect 26344 5370 26372 29446
rect 26436 29209 26464 29446
rect 26422 29200 26478 29209
rect 26422 29135 26478 29144
rect 26700 27532 26752 27538
rect 26700 27474 26752 27480
rect 26712 25498 26740 27474
rect 26792 27328 26844 27334
rect 26792 27270 26844 27276
rect 26804 26994 26832 27270
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26896 26874 26924 29582
rect 26804 26846 26924 26874
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26516 24880 26568 24886
rect 26516 24822 26568 24828
rect 26528 23730 26556 24822
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26528 23186 26556 23666
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26436 20398 26464 20742
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26436 19530 26464 20334
rect 26608 19712 26660 19718
rect 26608 19654 26660 19660
rect 26436 19514 26556 19530
rect 26436 19508 26568 19514
rect 26436 19502 26516 19508
rect 26516 19450 26568 19456
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26528 17202 26556 19314
rect 26620 18834 26648 19654
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26804 18222 26832 26846
rect 26884 24676 26936 24682
rect 26884 24618 26936 24624
rect 26896 24274 26924 24618
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 26896 24070 26924 24210
rect 26884 24064 26936 24070
rect 26882 24032 26884 24041
rect 26936 24032 26938 24041
rect 26882 23967 26938 23976
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27172 18834 27200 20198
rect 27264 19174 27292 29990
rect 27540 28082 27568 33254
rect 27724 33046 27752 33322
rect 29288 33046 29316 34002
rect 27712 33040 27764 33046
rect 27712 32982 27764 32988
rect 29276 33040 29328 33046
rect 29276 32982 29328 32988
rect 29380 32502 29408 35702
rect 31942 35663 31944 35672
rect 31996 35663 31998 35672
rect 31944 35634 31996 35640
rect 32036 35624 32088 35630
rect 32034 35592 32036 35601
rect 32088 35592 32090 35601
rect 32034 35527 32090 35536
rect 31668 35148 31720 35154
rect 31668 35090 31720 35096
rect 31680 35057 31708 35090
rect 31666 35048 31722 35057
rect 31666 34983 31722 34992
rect 32048 33862 32076 35527
rect 32128 34060 32180 34066
rect 32128 34002 32180 34008
rect 31208 33856 31260 33862
rect 31208 33798 31260 33804
rect 32036 33856 32088 33862
rect 32036 33798 32088 33804
rect 30564 33448 30616 33454
rect 30840 33448 30892 33454
rect 30564 33390 30616 33396
rect 30654 33416 30710 33425
rect 30576 32978 30604 33390
rect 30840 33390 30892 33396
rect 30654 33351 30656 33360
rect 30708 33351 30710 33360
rect 30656 33322 30708 33328
rect 30852 33046 30880 33390
rect 30840 33040 30892 33046
rect 30840 32982 30892 32988
rect 30564 32972 30616 32978
rect 30564 32914 30616 32920
rect 31220 32842 31248 33798
rect 32140 33590 32168 34002
rect 32128 33584 32180 33590
rect 32128 33526 32180 33532
rect 32128 33312 32180 33318
rect 32128 33254 32180 33260
rect 32140 33046 32168 33254
rect 31576 33040 31628 33046
rect 31576 32982 31628 32988
rect 32128 33040 32180 33046
rect 32128 32982 32180 32988
rect 31392 32972 31444 32978
rect 31392 32914 31444 32920
rect 31208 32836 31260 32842
rect 31208 32778 31260 32784
rect 31404 32502 31432 32914
rect 29368 32496 29420 32502
rect 29368 32438 29420 32444
rect 31392 32496 31444 32502
rect 31392 32438 31444 32444
rect 31588 32434 31616 32982
rect 31852 32768 31904 32774
rect 31852 32710 31904 32716
rect 31864 32434 31892 32710
rect 31576 32428 31628 32434
rect 31576 32370 31628 32376
rect 31852 32428 31904 32434
rect 31852 32370 31904 32376
rect 31588 32230 31616 32370
rect 31576 32224 31628 32230
rect 31576 32166 31628 32172
rect 29460 31272 29512 31278
rect 29460 31214 29512 31220
rect 29472 31142 29500 31214
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 29460 31136 29512 31142
rect 29460 31078 29512 31084
rect 30656 31136 30708 31142
rect 30656 31078 30708 31084
rect 29012 30258 29040 31078
rect 29092 30728 29144 30734
rect 29092 30670 29144 30676
rect 29276 30728 29328 30734
rect 29276 30670 29328 30676
rect 29104 30258 29132 30670
rect 29288 30326 29316 30670
rect 30668 30666 30696 31078
rect 31588 30938 31616 32166
rect 31024 30932 31076 30938
rect 31024 30874 31076 30880
rect 31576 30932 31628 30938
rect 31576 30874 31628 30880
rect 30656 30660 30708 30666
rect 30656 30602 30708 30608
rect 31036 30394 31064 30874
rect 31024 30388 31076 30394
rect 31024 30330 31076 30336
rect 29276 30320 29328 30326
rect 29276 30262 29328 30268
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29092 30252 29144 30258
rect 29092 30194 29144 30200
rect 27804 30184 27856 30190
rect 27804 30126 27856 30132
rect 29368 30184 29420 30190
rect 29368 30126 29420 30132
rect 29644 30184 29696 30190
rect 29644 30126 29696 30132
rect 27816 29850 27844 30126
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27816 29714 27844 29786
rect 28736 29714 28764 29990
rect 29380 29850 29408 30126
rect 29368 29844 29420 29850
rect 29368 29786 29420 29792
rect 29656 29730 29684 30126
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 30840 30048 30892 30054
rect 30840 29990 30892 29996
rect 29840 29850 29868 29990
rect 29828 29844 29880 29850
rect 29828 29786 29880 29792
rect 30852 29782 30880 29990
rect 27804 29708 27856 29714
rect 27804 29650 27856 29656
rect 28724 29708 28776 29714
rect 28724 29650 28776 29656
rect 29380 29702 29684 29730
rect 30840 29776 30892 29782
rect 30840 29718 30892 29724
rect 28172 29640 28224 29646
rect 29380 29594 29408 29702
rect 28172 29582 28224 29588
rect 28184 29481 28212 29582
rect 29288 29566 29408 29594
rect 29460 29572 29512 29578
rect 29288 29510 29316 29566
rect 29460 29514 29512 29520
rect 29276 29504 29328 29510
rect 28170 29472 28226 29481
rect 29276 29446 29328 29452
rect 28170 29407 28226 29416
rect 29472 29102 29500 29514
rect 29460 29096 29512 29102
rect 29460 29038 29512 29044
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27436 28008 27488 28014
rect 27436 27950 27488 27956
rect 27448 27538 27476 27950
rect 27436 27532 27488 27538
rect 27436 27474 27488 27480
rect 27448 26586 27476 27474
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 28092 26450 28120 26726
rect 28172 26580 28224 26586
rect 28172 26522 28224 26528
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 28184 26382 28212 26522
rect 28172 26376 28224 26382
rect 28172 26318 28224 26324
rect 31574 26098 31630 26107
rect 31574 26033 31630 26042
rect 31588 24954 31616 26033
rect 31666 25554 31722 25563
rect 31666 25489 31722 25498
rect 31576 24948 31628 24954
rect 31576 24890 31628 24896
rect 31680 24886 31708 25489
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 31772 25063 31800 25162
rect 31758 25054 31814 25063
rect 31758 24989 31814 24998
rect 31668 24880 31720 24886
rect 31668 24822 31720 24828
rect 27436 24064 27488 24070
rect 27436 24006 27488 24012
rect 31576 24064 31628 24070
rect 31576 24006 31628 24012
rect 27448 20466 27476 24006
rect 31588 23975 31616 24006
rect 31574 23966 31630 23975
rect 31574 23901 31630 23910
rect 32232 23866 32260 36586
rect 32324 33318 32352 37606
rect 32416 35154 32444 39782
rect 32968 39574 32996 40326
rect 34716 40186 34744 40326
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34704 40180 34756 40186
rect 34704 40122 34756 40128
rect 32956 39568 33008 39574
rect 32956 39510 33008 39516
rect 32772 38276 32824 38282
rect 32772 38218 32824 38224
rect 32784 37126 32812 38218
rect 32968 38214 32996 39510
rect 33324 39432 33376 39438
rect 33324 39374 33376 39380
rect 32956 38208 33008 38214
rect 32956 38150 33008 38156
rect 32968 37670 32996 38150
rect 32956 37664 33008 37670
rect 32956 37606 33008 37612
rect 32864 37460 32916 37466
rect 32916 37420 33088 37448
rect 32864 37402 32916 37408
rect 33060 37330 33088 37420
rect 32956 37324 33008 37330
rect 32956 37266 33008 37272
rect 33048 37324 33100 37330
rect 33048 37266 33100 37272
rect 32968 37194 32996 37266
rect 32956 37188 33008 37194
rect 32956 37130 33008 37136
rect 32772 37120 32824 37126
rect 32772 37062 32824 37068
rect 33336 36922 33364 39374
rect 34612 39296 34664 39302
rect 34612 39238 34664 39244
rect 33416 38344 33468 38350
rect 33416 38286 33468 38292
rect 33428 37398 33456 38286
rect 34624 37806 34652 39238
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34796 38276 34848 38282
rect 34796 38218 34848 38224
rect 34808 37806 34836 38218
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34612 37800 34664 37806
rect 34612 37742 34664 37748
rect 34796 37800 34848 37806
rect 34796 37742 34848 37748
rect 33692 37664 33744 37670
rect 33692 37606 33744 37612
rect 34980 37664 35032 37670
rect 34980 37606 35032 37612
rect 33416 37392 33468 37398
rect 33416 37334 33468 37340
rect 33324 36916 33376 36922
rect 33324 36858 33376 36864
rect 33704 36718 33732 37606
rect 34992 37398 35020 37606
rect 34980 37392 35032 37398
rect 34980 37334 35032 37340
rect 34336 37324 34388 37330
rect 34336 37266 34388 37272
rect 34348 37126 34376 37266
rect 34336 37120 34388 37126
rect 34336 37062 34388 37068
rect 32680 36712 32732 36718
rect 32680 36654 32732 36660
rect 33232 36712 33284 36718
rect 33232 36654 33284 36660
rect 33692 36712 33744 36718
rect 33692 36654 33744 36660
rect 32588 36644 32640 36650
rect 32588 36586 32640 36592
rect 32600 36106 32628 36586
rect 32588 36100 32640 36106
rect 32588 36042 32640 36048
rect 32692 36038 32720 36654
rect 33140 36236 33192 36242
rect 33140 36178 33192 36184
rect 32680 36032 32732 36038
rect 32680 35974 32732 35980
rect 32588 35624 32640 35630
rect 32586 35592 32588 35601
rect 32640 35592 32642 35601
rect 32586 35527 32642 35536
rect 32692 35290 32720 35974
rect 32496 35284 32548 35290
rect 32496 35226 32548 35232
rect 32680 35284 32732 35290
rect 32680 35226 32732 35232
rect 32956 35284 33008 35290
rect 32956 35226 33008 35232
rect 32404 35148 32456 35154
rect 32404 35090 32456 35096
rect 32416 34610 32444 35090
rect 32508 34950 32536 35226
rect 32496 34944 32548 34950
rect 32496 34886 32548 34892
rect 32968 34610 32996 35226
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32956 34604 33008 34610
rect 32956 34546 33008 34552
rect 32864 33856 32916 33862
rect 32864 33798 32916 33804
rect 32876 33522 32904 33798
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 32312 33312 32364 33318
rect 32312 33254 32364 33260
rect 32968 32026 32996 34546
rect 33152 33590 33180 36178
rect 33244 36106 33272 36654
rect 34152 36236 34204 36242
rect 34152 36178 34204 36184
rect 33232 36100 33284 36106
rect 33232 36042 33284 36048
rect 34164 36038 34192 36178
rect 34152 36032 34204 36038
rect 34152 35974 34204 35980
rect 33782 35728 33838 35737
rect 33782 35663 33838 35672
rect 33506 35592 33562 35601
rect 33506 35527 33562 35536
rect 33520 35494 33548 35527
rect 33796 35494 33824 35663
rect 34164 35630 34192 35974
rect 34152 35624 34204 35630
rect 34152 35566 34204 35572
rect 33508 35488 33560 35494
rect 33508 35430 33560 35436
rect 33784 35488 33836 35494
rect 33784 35430 33836 35436
rect 33140 33584 33192 33590
rect 33140 33526 33192 33532
rect 33152 33046 33180 33526
rect 33232 33448 33284 33454
rect 33232 33390 33284 33396
rect 33244 33318 33272 33390
rect 33232 33312 33284 33318
rect 33232 33254 33284 33260
rect 33140 33040 33192 33046
rect 33140 32982 33192 32988
rect 33244 32366 33272 33254
rect 34348 32434 34376 37062
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 36280 35222 36308 42094
rect 36372 38758 36400 43794
rect 37188 43648 37240 43654
rect 37188 43590 37240 43596
rect 37200 43382 37228 43590
rect 38488 43466 38516 43794
rect 38396 43450 38516 43466
rect 38384 43444 38516 43450
rect 38436 43438 38516 43444
rect 38384 43386 38436 43392
rect 37188 43376 37240 43382
rect 37188 43318 37240 43324
rect 37830 43344 37886 43353
rect 37830 43279 37832 43288
rect 37884 43279 37886 43288
rect 37832 43250 37884 43256
rect 38016 41064 38068 41070
rect 38016 41006 38068 41012
rect 38028 40934 38056 41006
rect 38016 40928 38068 40934
rect 38016 40870 38068 40876
rect 38028 39642 38056 40870
rect 38016 39636 38068 39642
rect 38016 39578 38068 39584
rect 36360 38752 36412 38758
rect 36360 38694 36412 38700
rect 36372 37874 36400 38694
rect 37096 38548 37148 38554
rect 37096 38490 37148 38496
rect 36636 37936 36688 37942
rect 36636 37878 36688 37884
rect 36360 37868 36412 37874
rect 36360 37810 36412 37816
rect 36648 36582 36676 37878
rect 37108 36650 37136 38490
rect 38488 38418 38516 43438
rect 38580 41750 38608 45562
rect 38764 44878 38792 46446
rect 38936 46436 38988 46442
rect 38936 46378 38988 46384
rect 38752 44872 38804 44878
rect 38752 44814 38804 44820
rect 38764 44742 38792 44814
rect 38752 44736 38804 44742
rect 38752 44678 38804 44684
rect 38764 43654 38792 44678
rect 38752 43648 38804 43654
rect 38752 43590 38804 43596
rect 38568 41744 38620 41750
rect 38568 41686 38620 41692
rect 38580 41546 38792 41562
rect 38568 41540 38804 41546
rect 38620 41534 38752 41540
rect 38568 41482 38620 41488
rect 38752 41482 38804 41488
rect 38844 41268 38896 41274
rect 38844 41210 38896 41216
rect 38752 41064 38804 41070
rect 38856 41052 38884 41210
rect 38804 41024 38884 41052
rect 38752 41006 38804 41012
rect 38660 40996 38712 41002
rect 38660 40938 38712 40944
rect 38672 40905 38700 40938
rect 38658 40896 38714 40905
rect 38658 40831 38714 40840
rect 38856 40594 38884 41024
rect 38844 40588 38896 40594
rect 38844 40530 38896 40536
rect 38568 40520 38620 40526
rect 38568 40462 38620 40468
rect 38580 40118 38608 40462
rect 38568 40112 38620 40118
rect 38568 40054 38620 40060
rect 38948 39914 38976 46378
rect 39212 46368 39264 46374
rect 39212 46310 39264 46316
rect 39224 46170 39252 46310
rect 39212 46164 39264 46170
rect 39212 46106 39264 46112
rect 39212 44872 39264 44878
rect 39212 44814 39264 44820
rect 39224 44538 39252 44814
rect 39212 44532 39264 44538
rect 39212 44474 39264 44480
rect 39488 43784 39540 43790
rect 39488 43726 39540 43732
rect 39500 43654 39528 43726
rect 39488 43648 39540 43654
rect 39488 43590 39540 43596
rect 39488 43104 39540 43110
rect 39488 43046 39540 43052
rect 39500 42770 39528 43046
rect 39488 42764 39540 42770
rect 39488 42706 39540 42712
rect 39396 41676 39448 41682
rect 39396 41618 39448 41624
rect 39304 41608 39356 41614
rect 39304 41550 39356 41556
rect 39120 40996 39172 41002
rect 39120 40938 39172 40944
rect 38936 39908 38988 39914
rect 38936 39850 38988 39856
rect 39028 39500 39080 39506
rect 39028 39442 39080 39448
rect 38936 39432 38988 39438
rect 38936 39374 38988 39380
rect 38476 38412 38528 38418
rect 38476 38354 38528 38360
rect 38752 38344 38804 38350
rect 38752 38286 38804 38292
rect 38292 38208 38344 38214
rect 38292 38150 38344 38156
rect 37280 37868 37332 37874
rect 37280 37810 37332 37816
rect 37096 36644 37148 36650
rect 37096 36586 37148 36592
rect 36636 36576 36688 36582
rect 36636 36518 36688 36524
rect 37292 36310 37320 37810
rect 38304 37398 38332 38150
rect 38292 37392 38344 37398
rect 38764 37346 38792 38286
rect 38844 38208 38896 38214
rect 38844 38150 38896 38156
rect 38856 37738 38884 38150
rect 38844 37732 38896 37738
rect 38844 37674 38896 37680
rect 38344 37340 38516 37346
rect 38292 37334 38516 37340
rect 38304 37318 38516 37334
rect 38764 37318 38884 37346
rect 38488 37262 38516 37318
rect 38476 37256 38528 37262
rect 38476 37198 38528 37204
rect 38752 37256 38804 37262
rect 38752 37198 38804 37204
rect 38384 37120 38436 37126
rect 38384 37062 38436 37068
rect 38396 36718 38424 37062
rect 37648 36712 37700 36718
rect 37648 36654 37700 36660
rect 38108 36712 38160 36718
rect 38108 36654 38160 36660
rect 38384 36712 38436 36718
rect 38384 36654 38436 36660
rect 37372 36576 37424 36582
rect 37372 36518 37424 36524
rect 37280 36304 37332 36310
rect 37280 36246 37332 36252
rect 37384 35630 37412 36518
rect 37660 36378 37688 36654
rect 37740 36644 37792 36650
rect 37740 36586 37792 36592
rect 37648 36372 37700 36378
rect 37648 36314 37700 36320
rect 37372 35624 37424 35630
rect 37372 35566 37424 35572
rect 36268 35216 36320 35222
rect 36268 35158 36320 35164
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 36280 34660 36308 35158
rect 37188 35012 37240 35018
rect 37188 34954 37240 34960
rect 36188 34632 36308 34660
rect 35532 33992 35584 33998
rect 35532 33934 35584 33940
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35544 33522 35572 33934
rect 35532 33516 35584 33522
rect 35532 33458 35584 33464
rect 35440 33448 35492 33454
rect 35438 33416 35440 33425
rect 35492 33416 35494 33425
rect 35438 33351 35494 33360
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 36188 32570 36216 34632
rect 36268 34400 36320 34406
rect 36268 34342 36320 34348
rect 36452 34400 36504 34406
rect 36452 34342 36504 34348
rect 36280 33590 36308 34342
rect 36464 33930 36492 34342
rect 37200 34134 37228 34954
rect 37384 34950 37412 35566
rect 37462 35048 37518 35057
rect 37660 35018 37688 36314
rect 37752 36242 37780 36586
rect 38120 36242 38148 36654
rect 37740 36236 37792 36242
rect 37740 36178 37792 36184
rect 38108 36236 38160 36242
rect 38396 36224 38424 36654
rect 38108 36178 38160 36184
rect 38212 36196 38424 36224
rect 38212 36122 38240 36196
rect 38120 36094 38240 36122
rect 38292 36100 38344 36106
rect 37462 34983 37518 34992
rect 37648 35012 37700 35018
rect 37476 34950 37504 34983
rect 37648 34954 37700 34960
rect 37372 34944 37424 34950
rect 37372 34886 37424 34892
rect 37464 34944 37516 34950
rect 37464 34886 37516 34892
rect 37280 34740 37332 34746
rect 37280 34682 37332 34688
rect 37292 34542 37320 34682
rect 38120 34542 38148 36094
rect 38292 36042 38344 36048
rect 38304 35834 38332 36042
rect 38384 36032 38436 36038
rect 38384 35974 38436 35980
rect 38396 35834 38424 35974
rect 38292 35828 38344 35834
rect 38292 35770 38344 35776
rect 38384 35828 38436 35834
rect 38384 35770 38436 35776
rect 38488 35222 38516 37198
rect 38764 36922 38792 37198
rect 38752 36916 38804 36922
rect 38752 36858 38804 36864
rect 38856 35766 38884 37318
rect 38948 37126 38976 39374
rect 39040 38962 39068 39442
rect 39028 38956 39080 38962
rect 39028 38898 39080 38904
rect 39040 38418 39068 38898
rect 39028 38412 39080 38418
rect 39028 38354 39080 38360
rect 39132 38282 39160 40938
rect 39316 40934 39344 41550
rect 39408 41070 39436 41618
rect 39396 41064 39448 41070
rect 39396 41006 39448 41012
rect 39304 40928 39356 40934
rect 39304 40870 39356 40876
rect 39408 40633 39436 41006
rect 39394 40624 39450 40633
rect 39394 40559 39396 40568
rect 39448 40559 39450 40568
rect 39396 40530 39448 40536
rect 39500 39506 39528 42706
rect 40052 42022 40080 46854
rect 40604 46714 40632 46990
rect 40592 46708 40644 46714
rect 40592 46650 40644 46656
rect 40696 46510 40724 46990
rect 43444 46912 43496 46918
rect 43444 46854 43496 46860
rect 43456 46578 43484 46854
rect 43444 46572 43496 46578
rect 43444 46514 43496 46520
rect 40684 46504 40736 46510
rect 40684 46446 40736 46452
rect 44376 46102 44404 47058
rect 46480 46912 46532 46918
rect 46480 46854 46532 46860
rect 45008 46640 45060 46646
rect 45008 46582 45060 46588
rect 44456 46436 44508 46442
rect 44456 46378 44508 46384
rect 40776 46096 40828 46102
rect 40776 46038 40828 46044
rect 44364 46096 44416 46102
rect 44364 46038 44416 46044
rect 40132 45892 40184 45898
rect 40132 45834 40184 45840
rect 40144 42226 40172 45834
rect 40500 44736 40552 44742
rect 40500 44678 40552 44684
rect 40512 44334 40540 44678
rect 40500 44328 40552 44334
rect 40500 44270 40552 44276
rect 40132 42220 40184 42226
rect 40132 42162 40184 42168
rect 40144 42106 40172 42162
rect 40144 42078 40264 42106
rect 40040 42016 40092 42022
rect 40040 41958 40092 41964
rect 40052 41682 40080 41958
rect 40040 41676 40092 41682
rect 40040 41618 40092 41624
rect 40236 41562 40264 42078
rect 40236 41534 40632 41562
rect 40236 41274 40264 41534
rect 40500 41472 40552 41478
rect 40500 41414 40552 41420
rect 40224 41268 40276 41274
rect 40224 41210 40276 41216
rect 40408 41132 40460 41138
rect 40408 41074 40460 41080
rect 39580 40928 39632 40934
rect 39580 40870 39632 40876
rect 40224 40928 40276 40934
rect 40224 40870 40276 40876
rect 39592 40594 39620 40870
rect 40236 40662 40264 40870
rect 40224 40656 40276 40662
rect 40222 40624 40224 40633
rect 40276 40624 40278 40633
rect 39580 40588 39632 40594
rect 40222 40559 40278 40568
rect 39580 40530 39632 40536
rect 39488 39500 39540 39506
rect 39488 39442 39540 39448
rect 39592 39302 39620 40530
rect 40420 39982 40448 41074
rect 40512 40390 40540 41414
rect 40604 41138 40632 41534
rect 40592 41132 40644 41138
rect 40592 41074 40644 41080
rect 40592 40996 40644 41002
rect 40592 40938 40644 40944
rect 40604 40882 40632 40938
rect 40604 40854 40724 40882
rect 40696 40662 40724 40854
rect 40788 40662 40816 46038
rect 44468 45422 44496 46378
rect 45020 46034 45048 46582
rect 45376 46572 45428 46578
rect 45376 46514 45428 46520
rect 45388 46034 45416 46514
rect 46112 46436 46164 46442
rect 46112 46378 46164 46384
rect 46124 46170 46152 46378
rect 46112 46164 46164 46170
rect 46112 46106 46164 46112
rect 45008 46028 45060 46034
rect 45008 45970 45060 45976
rect 45376 46028 45428 46034
rect 45376 45970 45428 45976
rect 44548 45552 44600 45558
rect 44548 45494 44600 45500
rect 44456 45416 44508 45422
rect 44456 45358 44508 45364
rect 43812 45280 43864 45286
rect 43812 45222 43864 45228
rect 42248 43648 42300 43654
rect 42248 43590 42300 43596
rect 42260 43382 42288 43590
rect 42248 43376 42300 43382
rect 42248 43318 42300 43324
rect 41236 42016 41288 42022
rect 41236 41958 41288 41964
rect 41248 41614 41276 41958
rect 41236 41608 41288 41614
rect 41236 41550 41288 41556
rect 41248 41070 41276 41550
rect 41604 41472 41656 41478
rect 41604 41414 41656 41420
rect 41236 41064 41288 41070
rect 40880 40990 41092 41018
rect 41236 41006 41288 41012
rect 41420 41064 41472 41070
rect 41420 41006 41472 41012
rect 40684 40656 40736 40662
rect 40684 40598 40736 40604
rect 40776 40656 40828 40662
rect 40776 40598 40828 40604
rect 40696 40508 40724 40598
rect 40880 40508 40908 40990
rect 41064 40934 41092 40990
rect 41052 40928 41104 40934
rect 40958 40896 41014 40905
rect 41052 40870 41104 40876
rect 40958 40831 41014 40840
rect 40972 40662 41000 40831
rect 40960 40656 41012 40662
rect 40960 40598 41012 40604
rect 40590 40488 40646 40497
rect 40696 40480 40908 40508
rect 41432 40474 41460 41006
rect 41616 40730 41644 41414
rect 42064 41268 42116 41274
rect 42064 41210 42116 41216
rect 41696 41132 41748 41138
rect 41696 41074 41748 41080
rect 41512 40724 41564 40730
rect 41512 40666 41564 40672
rect 41604 40724 41656 40730
rect 41604 40666 41656 40672
rect 40590 40423 40592 40432
rect 40644 40423 40646 40432
rect 41064 40446 41460 40474
rect 41524 40474 41552 40666
rect 41616 40633 41644 40666
rect 41602 40624 41658 40633
rect 41602 40559 41658 40568
rect 41524 40446 41644 40474
rect 40592 40394 40644 40400
rect 40500 40384 40552 40390
rect 40500 40326 40552 40332
rect 41064 40202 41092 40446
rect 41616 40390 41644 40446
rect 41512 40384 41564 40390
rect 40512 40174 41092 40202
rect 41248 40344 41512 40372
rect 40512 40118 40540 40174
rect 40500 40112 40552 40118
rect 40500 40054 40552 40060
rect 40684 40044 40736 40050
rect 40960 40044 41012 40050
rect 40736 40004 40960 40032
rect 40684 39986 40736 39992
rect 40960 39986 41012 39992
rect 40316 39976 40368 39982
rect 40316 39918 40368 39924
rect 40408 39976 40460 39982
rect 40408 39918 40460 39924
rect 40328 39681 40356 39918
rect 40868 39840 40920 39846
rect 40868 39782 40920 39788
rect 40314 39672 40370 39681
rect 40314 39607 40370 39616
rect 39948 39500 40000 39506
rect 39948 39442 40000 39448
rect 39580 39296 39632 39302
rect 39580 39238 39632 39244
rect 39960 38350 39988 39442
rect 40040 39296 40092 39302
rect 40040 39238 40092 39244
rect 40684 39296 40736 39302
rect 40684 39238 40736 39244
rect 40052 38350 40080 39238
rect 40696 38962 40724 39238
rect 40408 38956 40460 38962
rect 40408 38898 40460 38904
rect 40684 38956 40736 38962
rect 40684 38898 40736 38904
rect 40420 38554 40448 38898
rect 40224 38548 40276 38554
rect 40224 38490 40276 38496
rect 40408 38548 40460 38554
rect 40408 38490 40460 38496
rect 40236 38418 40264 38490
rect 40224 38412 40276 38418
rect 40224 38354 40276 38360
rect 39948 38344 40000 38350
rect 39948 38286 40000 38292
rect 40040 38344 40092 38350
rect 40040 38286 40092 38292
rect 39120 38276 39172 38282
rect 39120 38218 39172 38224
rect 39856 38276 39908 38282
rect 39856 38218 39908 38224
rect 39868 37874 39896 38218
rect 39960 38162 39988 38286
rect 40880 38282 40908 39782
rect 40960 38548 41012 38554
rect 40960 38490 41012 38496
rect 40868 38276 40920 38282
rect 40868 38218 40920 38224
rect 40040 38208 40092 38214
rect 39960 38156 40040 38162
rect 39960 38150 40092 38156
rect 39960 38134 40080 38150
rect 39856 37868 39908 37874
rect 39856 37810 39908 37816
rect 40972 37330 41000 38490
rect 41248 38418 41276 40344
rect 41512 40326 41564 40332
rect 41604 40384 41656 40390
rect 41604 40326 41656 40332
rect 41708 40050 41736 41074
rect 42076 41002 42104 41210
rect 42064 40996 42116 41002
rect 42064 40938 42116 40944
rect 41696 40044 41748 40050
rect 41696 39986 41748 39992
rect 43824 39506 43852 45222
rect 44468 45014 44496 45358
rect 44560 45082 44588 45494
rect 45388 45286 45416 45970
rect 45928 45960 45980 45966
rect 45928 45902 45980 45908
rect 45940 45830 45968 45902
rect 46492 45830 46520 46854
rect 46676 46034 46704 47058
rect 47308 47048 47360 47054
rect 47308 46990 47360 46996
rect 47492 47048 47544 47054
rect 47492 46990 47544 46996
rect 47320 46918 47348 46990
rect 47400 46980 47452 46986
rect 47400 46922 47452 46928
rect 47308 46912 47360 46918
rect 47308 46854 47360 46860
rect 46940 46436 46992 46442
rect 46940 46378 46992 46384
rect 46952 46170 46980 46378
rect 46940 46164 46992 46170
rect 46940 46106 46992 46112
rect 47320 46102 47348 46854
rect 47412 46714 47440 46922
rect 47400 46708 47452 46714
rect 47400 46650 47452 46656
rect 47412 46442 47440 46650
rect 47504 46510 47532 46990
rect 48688 46912 48740 46918
rect 48688 46854 48740 46860
rect 48700 46510 48728 46854
rect 50172 46510 50200 47058
rect 50540 46578 50568 47058
rect 50908 46714 50936 47058
rect 51356 47048 51408 47054
rect 51356 46990 51408 46996
rect 50896 46708 50948 46714
rect 50896 46650 50948 46656
rect 51368 46578 51396 46990
rect 51724 46912 51776 46918
rect 51724 46854 51776 46860
rect 50528 46572 50580 46578
rect 50528 46514 50580 46520
rect 51356 46572 51408 46578
rect 51356 46514 51408 46520
rect 47492 46504 47544 46510
rect 47492 46446 47544 46452
rect 48688 46504 48740 46510
rect 48688 46446 48740 46452
rect 50160 46504 50212 46510
rect 50160 46446 50212 46452
rect 51172 46504 51224 46510
rect 51448 46504 51500 46510
rect 51172 46446 51224 46452
rect 51368 46452 51448 46458
rect 51368 46446 51500 46452
rect 47400 46436 47452 46442
rect 47400 46378 47452 46384
rect 47308 46096 47360 46102
rect 47308 46038 47360 46044
rect 46664 46028 46716 46034
rect 46664 45970 46716 45976
rect 45928 45824 45980 45830
rect 45928 45766 45980 45772
rect 46480 45824 46532 45830
rect 46480 45766 46532 45772
rect 46112 45416 46164 45422
rect 46112 45358 46164 45364
rect 45376 45280 45428 45286
rect 45376 45222 45428 45228
rect 44548 45076 44600 45082
rect 44548 45018 44600 45024
rect 44732 45076 44784 45082
rect 44732 45018 44784 45024
rect 45468 45076 45520 45082
rect 45468 45018 45520 45024
rect 44456 45008 44508 45014
rect 44456 44950 44508 44956
rect 44560 44946 44588 45018
rect 44364 44940 44416 44946
rect 44364 44882 44416 44888
rect 44548 44940 44600 44946
rect 44548 44882 44600 44888
rect 44376 44470 44404 44882
rect 44364 44464 44416 44470
rect 44364 44406 44416 44412
rect 44376 42770 44404 44406
rect 44560 43858 44588 44882
rect 44548 43852 44600 43858
rect 44548 43794 44600 43800
rect 44548 43648 44600 43654
rect 44548 43590 44600 43596
rect 44560 42838 44588 43590
rect 44744 42906 44772 45018
rect 45480 44946 45508 45018
rect 45468 44940 45520 44946
rect 45468 44882 45520 44888
rect 45468 44464 45520 44470
rect 45468 44406 45520 44412
rect 45284 43852 45336 43858
rect 45284 43794 45336 43800
rect 45100 43784 45152 43790
rect 45100 43726 45152 43732
rect 45112 43654 45140 43726
rect 45100 43648 45152 43654
rect 45100 43590 45152 43596
rect 44824 43308 44876 43314
rect 44824 43250 44876 43256
rect 44836 43178 44864 43250
rect 44824 43172 44876 43178
rect 44824 43114 44876 43120
rect 44836 42906 44864 43114
rect 44732 42900 44784 42906
rect 44732 42842 44784 42848
rect 44824 42900 44876 42906
rect 44824 42842 44876 42848
rect 45296 42838 45324 43794
rect 44548 42832 44600 42838
rect 44548 42774 44600 42780
rect 45284 42832 45336 42838
rect 45284 42774 45336 42780
rect 45480 42786 45508 44406
rect 45560 44192 45612 44198
rect 45560 44134 45612 44140
rect 45572 43994 45600 44134
rect 45560 43988 45612 43994
rect 45560 43930 45612 43936
rect 45836 43988 45888 43994
rect 45836 43930 45888 43936
rect 45848 43858 45876 43930
rect 45836 43852 45888 43858
rect 45836 43794 45888 43800
rect 44364 42764 44416 42770
rect 44364 42706 44416 42712
rect 44560 42634 44588 42774
rect 45480 42770 45600 42786
rect 45480 42764 45612 42770
rect 45480 42758 45560 42764
rect 45560 42706 45612 42712
rect 44548 42628 44600 42634
rect 44548 42570 44600 42576
rect 46124 42140 46152 45358
rect 46492 44810 46520 45766
rect 46676 45626 46704 45970
rect 47320 45830 47348 46038
rect 48700 45966 48728 46446
rect 50300 46268 50596 46288
rect 50356 46266 50380 46268
rect 50436 46266 50460 46268
rect 50516 46266 50540 46268
rect 50378 46214 50380 46266
rect 50442 46214 50454 46266
rect 50516 46214 50518 46266
rect 50356 46212 50380 46214
rect 50436 46212 50460 46214
rect 50516 46212 50540 46214
rect 50300 46192 50596 46212
rect 51184 46034 51212 46446
rect 51368 46430 51488 46446
rect 51368 46374 51396 46430
rect 51356 46368 51408 46374
rect 51356 46310 51408 46316
rect 51172 46028 51224 46034
rect 51172 45970 51224 45976
rect 48688 45960 48740 45966
rect 48688 45902 48740 45908
rect 47308 45824 47360 45830
rect 47308 45766 47360 45772
rect 46664 45620 46716 45626
rect 46664 45562 46716 45568
rect 47320 45082 47348 45766
rect 47676 45552 47728 45558
rect 47676 45494 47728 45500
rect 47308 45076 47360 45082
rect 47308 45018 47360 45024
rect 46848 44940 46900 44946
rect 46848 44882 46900 44888
rect 46572 44872 46624 44878
rect 46572 44814 46624 44820
rect 46480 44804 46532 44810
rect 46480 44746 46532 44752
rect 46584 43994 46612 44814
rect 46860 44334 46888 44882
rect 47124 44804 47176 44810
rect 47124 44746 47176 44752
rect 46848 44328 46900 44334
rect 46848 44270 46900 44276
rect 47136 44198 47164 44746
rect 47688 44470 47716 45494
rect 50300 45180 50596 45200
rect 50356 45178 50380 45180
rect 50436 45178 50460 45180
rect 50516 45178 50540 45180
rect 50378 45126 50380 45178
rect 50442 45126 50454 45178
rect 50516 45126 50518 45178
rect 50356 45124 50380 45126
rect 50436 45124 50460 45126
rect 50516 45124 50540 45126
rect 50300 45104 50596 45124
rect 47676 44464 47728 44470
rect 47676 44406 47728 44412
rect 51264 44328 51316 44334
rect 51264 44270 51316 44276
rect 47124 44192 47176 44198
rect 47124 44134 47176 44140
rect 50712 44192 50764 44198
rect 50712 44134 50764 44140
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 46572 43988 46624 43994
rect 46572 43930 46624 43936
rect 46584 42906 46612 43930
rect 46756 43648 46808 43654
rect 46756 43590 46808 43596
rect 46572 42900 46624 42906
rect 46572 42842 46624 42848
rect 46584 42770 46612 42842
rect 46768 42770 46796 43590
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 46572 42764 46624 42770
rect 46572 42706 46624 42712
rect 46756 42764 46808 42770
rect 46756 42706 46808 42712
rect 46296 42152 46348 42158
rect 46124 42112 46296 42140
rect 46124 41682 46152 42112
rect 46296 42094 46348 42100
rect 49516 42084 49568 42090
rect 49516 42026 49568 42032
rect 46756 42016 46808 42022
rect 47676 42016 47728 42022
rect 46808 41976 46888 42004
rect 46756 41958 46808 41964
rect 46112 41676 46164 41682
rect 46112 41618 46164 41624
rect 46756 41676 46808 41682
rect 46756 41618 46808 41624
rect 45468 41472 45520 41478
rect 45468 41414 45520 41420
rect 45480 41206 45508 41414
rect 46768 41206 46796 41618
rect 45468 41200 45520 41206
rect 45468 41142 45520 41148
rect 46756 41200 46808 41206
rect 46756 41142 46808 41148
rect 44652 40594 44864 40610
rect 44456 40588 44508 40594
rect 44652 40588 44876 40594
rect 44652 40582 44824 40588
rect 44652 40576 44680 40582
rect 44508 40548 44680 40576
rect 44456 40530 44508 40536
rect 44824 40530 44876 40536
rect 46572 40588 46624 40594
rect 46572 40530 46624 40536
rect 44638 40488 44694 40497
rect 44364 40452 44416 40458
rect 44638 40423 44640 40432
rect 44364 40394 44416 40400
rect 44692 40423 44694 40432
rect 44640 40394 44692 40400
rect 44180 40384 44232 40390
rect 44180 40326 44232 40332
rect 44192 39506 44220 40326
rect 44272 39908 44324 39914
rect 44272 39850 44324 39856
rect 44284 39642 44312 39850
rect 44376 39642 44404 40394
rect 44456 40044 44508 40050
rect 44456 39986 44508 39992
rect 44272 39636 44324 39642
rect 44272 39578 44324 39584
rect 44364 39636 44416 39642
rect 44364 39578 44416 39584
rect 44468 39506 44496 39986
rect 44836 39574 44864 40530
rect 44916 40520 44968 40526
rect 45744 40520 45796 40526
rect 44916 40462 44968 40468
rect 45572 40468 45744 40474
rect 45572 40462 45796 40468
rect 44928 40050 44956 40462
rect 45572 40446 45784 40462
rect 45572 40390 45600 40446
rect 46584 40390 46612 40530
rect 45560 40384 45612 40390
rect 45560 40326 45612 40332
rect 45744 40384 45796 40390
rect 45744 40326 45796 40332
rect 46020 40384 46072 40390
rect 46020 40326 46072 40332
rect 46572 40384 46624 40390
rect 46572 40326 46624 40332
rect 44916 40044 44968 40050
rect 44916 39986 44968 39992
rect 44824 39568 44876 39574
rect 44824 39510 44876 39516
rect 43812 39500 43864 39506
rect 43812 39442 43864 39448
rect 44180 39500 44232 39506
rect 44180 39442 44232 39448
rect 44456 39500 44508 39506
rect 44456 39442 44508 39448
rect 44916 39500 44968 39506
rect 44916 39442 44968 39448
rect 42616 39296 42668 39302
rect 42616 39238 42668 39244
rect 42156 39024 42208 39030
rect 42154 38992 42156 39001
rect 42208 38992 42210 39001
rect 42154 38927 42210 38936
rect 41236 38412 41288 38418
rect 41236 38354 41288 38360
rect 41236 38208 41288 38214
rect 41236 38150 41288 38156
rect 40960 37324 41012 37330
rect 40960 37266 41012 37272
rect 38936 37120 38988 37126
rect 38936 37062 38988 37068
rect 38844 35760 38896 35766
rect 38844 35702 38896 35708
rect 38476 35216 38528 35222
rect 38476 35158 38528 35164
rect 38488 35086 38516 35158
rect 38476 35080 38528 35086
rect 38476 35022 38528 35028
rect 38752 35080 38804 35086
rect 38752 35022 38804 35028
rect 38292 34604 38344 34610
rect 38292 34546 38344 34552
rect 37280 34536 37332 34542
rect 37280 34478 37332 34484
rect 37372 34536 37424 34542
rect 37372 34478 37424 34484
rect 38108 34536 38160 34542
rect 38108 34478 38160 34484
rect 38200 34536 38252 34542
rect 38200 34478 38252 34484
rect 37384 34406 37412 34478
rect 38212 34406 38240 34478
rect 37372 34400 37424 34406
rect 37372 34342 37424 34348
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 37188 34128 37240 34134
rect 37188 34070 37240 34076
rect 36452 33924 36504 33930
rect 36452 33866 36504 33872
rect 36268 33584 36320 33590
rect 36268 33526 36320 33532
rect 37384 33454 37412 34342
rect 38304 33454 38332 34546
rect 38764 34134 38792 35022
rect 38856 34746 38884 35702
rect 41248 35698 41276 38150
rect 42156 37256 42208 37262
rect 42156 37198 42208 37204
rect 42168 36718 42196 37198
rect 42156 36712 42208 36718
rect 42156 36654 42208 36660
rect 41236 35692 41288 35698
rect 41236 35634 41288 35640
rect 42432 35556 42484 35562
rect 42432 35498 42484 35504
rect 39764 35488 39816 35494
rect 39764 35430 39816 35436
rect 39580 35216 39632 35222
rect 39580 35158 39632 35164
rect 39672 35216 39724 35222
rect 39672 35158 39724 35164
rect 39592 35018 39620 35158
rect 39580 35012 39632 35018
rect 39580 34954 39632 34960
rect 39684 34746 39712 35158
rect 38844 34740 38896 34746
rect 38844 34682 38896 34688
rect 39672 34740 39724 34746
rect 39672 34682 39724 34688
rect 39210 34640 39266 34649
rect 39210 34575 39266 34584
rect 39224 34542 39252 34575
rect 39684 34542 39712 34682
rect 39776 34542 39804 35430
rect 42444 35154 42472 35498
rect 42628 35222 42656 39238
rect 44928 39030 44956 39442
rect 44916 39024 44968 39030
rect 44916 38966 44968 38972
rect 44732 38888 44784 38894
rect 44732 38830 44784 38836
rect 44546 37496 44602 37505
rect 44546 37431 44602 37440
rect 44560 37330 44588 37431
rect 44548 37324 44600 37330
rect 44548 37266 44600 37272
rect 44744 37126 44772 38830
rect 44822 37496 44878 37505
rect 44822 37431 44878 37440
rect 44836 37330 44864 37431
rect 44824 37324 44876 37330
rect 44824 37266 44876 37272
rect 44916 37256 44968 37262
rect 44916 37198 44968 37204
rect 45192 37256 45244 37262
rect 45192 37198 45244 37204
rect 44732 37120 44784 37126
rect 44732 37062 44784 37068
rect 43720 36644 43772 36650
rect 43720 36586 43772 36592
rect 43732 35630 43760 36586
rect 43720 35624 43772 35630
rect 43720 35566 43772 35572
rect 43536 35556 43588 35562
rect 43536 35498 43588 35504
rect 43260 35488 43312 35494
rect 43260 35430 43312 35436
rect 42616 35216 42668 35222
rect 42616 35158 42668 35164
rect 42432 35148 42484 35154
rect 42432 35090 42484 35096
rect 42984 35148 43036 35154
rect 42984 35090 43036 35096
rect 41604 34672 41656 34678
rect 41604 34614 41656 34620
rect 39212 34536 39264 34542
rect 39212 34478 39264 34484
rect 39672 34536 39724 34542
rect 39672 34478 39724 34484
rect 39764 34536 39816 34542
rect 39764 34478 39816 34484
rect 41512 34536 41564 34542
rect 41512 34478 41564 34484
rect 39396 34400 39448 34406
rect 39396 34342 39448 34348
rect 39488 34400 39540 34406
rect 39488 34342 39540 34348
rect 38752 34128 38804 34134
rect 38752 34070 38804 34076
rect 39408 34066 39436 34342
rect 38844 34060 38896 34066
rect 38844 34002 38896 34008
rect 39396 34060 39448 34066
rect 39396 34002 39448 34008
rect 38750 33688 38806 33697
rect 38750 33623 38806 33632
rect 38764 33590 38792 33623
rect 38752 33584 38804 33590
rect 38658 33552 38714 33561
rect 38752 33526 38804 33532
rect 38658 33487 38660 33496
rect 38712 33487 38714 33496
rect 38660 33458 38712 33464
rect 37372 33448 37424 33454
rect 37372 33390 37424 33396
rect 38292 33448 38344 33454
rect 38658 33416 38714 33425
rect 38292 33390 38344 33396
rect 38304 33318 38332 33390
rect 38580 33386 38658 33402
rect 38568 33380 38658 33386
rect 38620 33374 38658 33380
rect 38856 33386 38884 34002
rect 39500 33697 39528 34342
rect 39486 33688 39542 33697
rect 39486 33623 39542 33632
rect 38658 33351 38714 33360
rect 38844 33380 38896 33386
rect 38568 33322 38620 33328
rect 38844 33322 38896 33328
rect 38292 33312 38344 33318
rect 38292 33254 38344 33260
rect 37924 32972 37976 32978
rect 37924 32914 37976 32920
rect 37188 32836 37240 32842
rect 37188 32778 37240 32784
rect 37200 32570 37228 32778
rect 37936 32774 37964 32914
rect 37924 32768 37976 32774
rect 37924 32710 37976 32716
rect 36176 32564 36228 32570
rect 36176 32506 36228 32512
rect 37188 32564 37240 32570
rect 37188 32506 37240 32512
rect 34336 32428 34388 32434
rect 34336 32370 34388 32376
rect 36188 32366 36216 32506
rect 33232 32360 33284 32366
rect 33232 32302 33284 32308
rect 36176 32360 36228 32366
rect 36176 32302 36228 32308
rect 35072 32224 35124 32230
rect 35072 32166 35124 32172
rect 36544 32224 36596 32230
rect 36544 32166 36596 32172
rect 36636 32224 36688 32230
rect 36636 32166 36688 32172
rect 32956 32020 33008 32026
rect 32956 31962 33008 31968
rect 35084 31890 35112 32166
rect 35072 31884 35124 31890
rect 35124 31844 35296 31872
rect 35072 31826 35124 31832
rect 34796 31748 34848 31754
rect 34796 31690 34848 31696
rect 34808 30870 34836 31690
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35268 31414 35296 31844
rect 35256 31408 35308 31414
rect 35256 31350 35308 31356
rect 35164 31340 35216 31346
rect 35164 31282 35216 31288
rect 35624 31340 35676 31346
rect 35624 31282 35676 31288
rect 35176 30938 35204 31282
rect 35164 30932 35216 30938
rect 35164 30874 35216 30880
rect 34796 30864 34848 30870
rect 34796 30806 34848 30812
rect 35636 30802 35664 31282
rect 35900 31272 35952 31278
rect 35900 31214 35952 31220
rect 35624 30796 35676 30802
rect 35624 30738 35676 30744
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 35716 30184 35768 30190
rect 35912 30138 35940 31214
rect 36360 30796 36412 30802
rect 36360 30738 36412 30744
rect 36372 30598 36400 30738
rect 36360 30592 36412 30598
rect 36360 30534 36412 30540
rect 35768 30132 35940 30138
rect 35716 30126 35940 30132
rect 35728 30110 35940 30126
rect 35912 29510 35940 30110
rect 36556 29850 36584 32166
rect 36648 32026 36676 32166
rect 36636 32020 36688 32026
rect 36636 31962 36688 31968
rect 36728 31272 36780 31278
rect 36728 31214 36780 31220
rect 36740 30870 36768 31214
rect 36728 30864 36780 30870
rect 36728 30806 36780 30812
rect 37200 30802 37228 32506
rect 37936 32366 37964 32710
rect 40960 32428 41012 32434
rect 40960 32370 41012 32376
rect 37924 32360 37976 32366
rect 37924 32302 37976 32308
rect 40972 32026 41000 32370
rect 41236 32292 41288 32298
rect 41236 32234 41288 32240
rect 40960 32020 41012 32026
rect 40960 31962 41012 31968
rect 40972 31822 41000 31962
rect 41248 31890 41276 32234
rect 41524 31958 41552 34478
rect 41616 32502 41644 34614
rect 42892 34536 42944 34542
rect 42892 34478 42944 34484
rect 42904 33862 42932 34478
rect 42892 33856 42944 33862
rect 42892 33798 42944 33804
rect 41880 33448 41932 33454
rect 41880 33390 41932 33396
rect 41788 32768 41840 32774
rect 41892 32756 41920 33390
rect 42340 33312 42392 33318
rect 42340 33254 42392 33260
rect 41972 32972 42024 32978
rect 41972 32914 42024 32920
rect 41984 32774 42012 32914
rect 42352 32842 42380 33254
rect 42340 32836 42392 32842
rect 42340 32778 42392 32784
rect 41840 32728 41920 32756
rect 41788 32710 41840 32716
rect 41604 32496 41656 32502
rect 41604 32438 41656 32444
rect 41616 32366 41644 32438
rect 41604 32360 41656 32366
rect 41604 32302 41656 32308
rect 41512 31952 41564 31958
rect 41512 31894 41564 31900
rect 41892 31890 41920 32728
rect 41972 32768 42024 32774
rect 41972 32710 42024 32716
rect 41984 32230 42012 32710
rect 42352 32366 42380 32778
rect 42432 32768 42484 32774
rect 42432 32710 42484 32716
rect 42444 32502 42472 32710
rect 42996 32502 43024 35090
rect 43272 34950 43300 35430
rect 43260 34944 43312 34950
rect 43260 34886 43312 34892
rect 43272 34542 43300 34886
rect 43548 34649 43576 35498
rect 44364 35488 44416 35494
rect 44364 35430 44416 35436
rect 43812 35216 43864 35222
rect 43732 35176 43812 35204
rect 43534 34640 43590 34649
rect 43534 34575 43590 34584
rect 43732 34542 43760 35176
rect 43812 35158 43864 35164
rect 43812 34944 43864 34950
rect 43812 34886 43864 34892
rect 43824 34542 43852 34886
rect 44376 34762 44404 35430
rect 44008 34734 44404 34762
rect 44008 34542 44036 34734
rect 44376 34678 44404 34734
rect 44272 34672 44324 34678
rect 44272 34614 44324 34620
rect 44364 34672 44416 34678
rect 44364 34614 44416 34620
rect 43260 34536 43312 34542
rect 43260 34478 43312 34484
rect 43720 34536 43772 34542
rect 43720 34478 43772 34484
rect 43812 34536 43864 34542
rect 43812 34478 43864 34484
rect 43996 34536 44048 34542
rect 43996 34478 44048 34484
rect 43732 33561 43760 34478
rect 44284 34066 44312 34614
rect 44272 34060 44324 34066
rect 44272 34002 44324 34008
rect 43812 33992 43864 33998
rect 43812 33934 43864 33940
rect 43718 33552 43774 33561
rect 43718 33487 43774 33496
rect 43824 32910 43852 33934
rect 43444 32904 43496 32910
rect 43444 32846 43496 32852
rect 43812 32904 43864 32910
rect 43812 32846 43864 32852
rect 44088 32904 44140 32910
rect 44088 32846 44140 32852
rect 42432 32496 42484 32502
rect 42432 32438 42484 32444
rect 42984 32496 43036 32502
rect 42984 32438 43036 32444
rect 42996 32366 43024 32438
rect 42340 32360 42392 32366
rect 42340 32302 42392 32308
rect 42984 32360 43036 32366
rect 42984 32302 43036 32308
rect 42708 32292 42760 32298
rect 42708 32234 42760 32240
rect 41972 32224 42024 32230
rect 41972 32166 42024 32172
rect 41236 31884 41288 31890
rect 41236 31826 41288 31832
rect 41880 31884 41932 31890
rect 41880 31826 41932 31832
rect 40960 31816 41012 31822
rect 40960 31758 41012 31764
rect 41892 31754 41920 31826
rect 41880 31748 41932 31754
rect 41880 31690 41932 31696
rect 41984 31414 42012 32166
rect 42720 32026 42748 32234
rect 42800 32224 42852 32230
rect 42800 32166 42852 32172
rect 42812 32026 42840 32166
rect 42708 32020 42760 32026
rect 42708 31962 42760 31968
rect 42800 32020 42852 32026
rect 42800 31962 42852 31968
rect 42720 31822 42748 31962
rect 42708 31816 42760 31822
rect 42708 31758 42760 31764
rect 43352 31816 43404 31822
rect 43456 31804 43484 32846
rect 44100 32570 44128 32846
rect 44088 32564 44140 32570
rect 44088 32506 44140 32512
rect 44364 32360 44416 32366
rect 44364 32302 44416 32308
rect 44376 32026 44404 32302
rect 44548 32224 44600 32230
rect 44548 32166 44600 32172
rect 44364 32020 44416 32026
rect 44364 31962 44416 31968
rect 44560 31958 44588 32166
rect 44548 31952 44600 31958
rect 44548 31894 44600 31900
rect 43404 31776 43484 31804
rect 43352 31758 43404 31764
rect 41972 31408 42024 31414
rect 41972 31350 42024 31356
rect 41236 31340 41288 31346
rect 41236 31282 41288 31288
rect 41788 31340 41840 31346
rect 41788 31282 41840 31288
rect 43260 31340 43312 31346
rect 43260 31282 43312 31288
rect 40776 31272 40828 31278
rect 40776 31214 40828 31220
rect 38108 31204 38160 31210
rect 38108 31146 38160 31152
rect 37924 31136 37976 31142
rect 37924 31078 37976 31084
rect 37188 30796 37240 30802
rect 37188 30738 37240 30744
rect 37556 30728 37608 30734
rect 37556 30670 37608 30676
rect 37936 30682 37964 31078
rect 38016 30728 38068 30734
rect 37936 30676 38016 30682
rect 37936 30670 38068 30676
rect 37464 30592 37516 30598
rect 37464 30534 37516 30540
rect 37476 30394 37504 30534
rect 37464 30388 37516 30394
rect 37464 30330 37516 30336
rect 37568 30326 37596 30670
rect 37936 30654 38056 30670
rect 37556 30320 37608 30326
rect 37556 30262 37608 30268
rect 37936 30190 37964 30654
rect 38120 30274 38148 31146
rect 40788 30818 40816 31214
rect 40788 30802 41000 30818
rect 38660 30796 38712 30802
rect 38660 30738 38712 30744
rect 40788 30796 41012 30802
rect 40788 30790 40960 30796
rect 38292 30660 38344 30666
rect 38292 30602 38344 30608
rect 38028 30246 38148 30274
rect 38028 30190 38056 30246
rect 37280 30184 37332 30190
rect 37280 30126 37332 30132
rect 37464 30184 37516 30190
rect 37464 30126 37516 30132
rect 37924 30184 37976 30190
rect 37924 30126 37976 30132
rect 38016 30184 38068 30190
rect 38016 30126 38068 30132
rect 37004 30048 37056 30054
rect 37004 29990 37056 29996
rect 36544 29844 36596 29850
rect 36544 29786 36596 29792
rect 37016 29714 37044 29990
rect 37292 29714 37320 30126
rect 37476 29850 37504 30126
rect 37924 30048 37976 30054
rect 38028 30002 38056 30126
rect 37976 29996 38056 30002
rect 37924 29990 38056 29996
rect 37936 29974 38056 29990
rect 37464 29844 37516 29850
rect 37464 29786 37516 29792
rect 37004 29708 37056 29714
rect 37004 29650 37056 29656
rect 37280 29708 37332 29714
rect 37280 29650 37332 29656
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35452 27606 35480 29106
rect 37936 28490 37964 29974
rect 38304 29714 38332 30602
rect 38672 30598 38700 30738
rect 40788 30734 40816 30790
rect 40960 30738 41012 30744
rect 40776 30728 40828 30734
rect 40776 30670 40828 30676
rect 40500 30660 40552 30666
rect 40500 30602 40552 30608
rect 38660 30592 38712 30598
rect 38660 30534 38712 30540
rect 38292 29708 38344 29714
rect 38292 29650 38344 29656
rect 40512 29578 40540 30602
rect 40972 29850 41000 30738
rect 40960 29844 41012 29850
rect 40960 29786 41012 29792
rect 40972 29714 41000 29786
rect 41248 29714 41276 31282
rect 41800 30870 41828 31282
rect 42064 31136 42116 31142
rect 42064 31078 42116 31084
rect 42432 31136 42484 31142
rect 42432 31078 42484 31084
rect 41604 30864 41656 30870
rect 41604 30806 41656 30812
rect 41788 30864 41840 30870
rect 41788 30806 41840 30812
rect 41616 30666 41644 30806
rect 41696 30796 41748 30802
rect 41696 30738 41748 30744
rect 41880 30796 41932 30802
rect 41880 30738 41932 30744
rect 41708 30705 41736 30738
rect 41694 30696 41750 30705
rect 41604 30660 41656 30666
rect 41694 30631 41750 30640
rect 41604 30602 41656 30608
rect 41604 30184 41656 30190
rect 41604 30126 41656 30132
rect 40960 29708 41012 29714
rect 40960 29650 41012 29656
rect 41236 29708 41288 29714
rect 41236 29650 41288 29656
rect 40500 29572 40552 29578
rect 40500 29514 40552 29520
rect 41616 29510 41644 30126
rect 41788 29844 41840 29850
rect 41788 29786 41840 29792
rect 41800 29714 41828 29786
rect 41788 29708 41840 29714
rect 41788 29650 41840 29656
rect 41604 29504 41656 29510
rect 41604 29446 41656 29452
rect 37924 28484 37976 28490
rect 37924 28426 37976 28432
rect 35440 27600 35492 27606
rect 35440 27542 35492 27548
rect 41892 27130 41920 30738
rect 42076 29850 42104 31078
rect 42444 30802 42472 31078
rect 42432 30796 42484 30802
rect 42432 30738 42484 30744
rect 43168 30796 43220 30802
rect 43168 30738 43220 30744
rect 43180 30326 43208 30738
rect 43272 30598 43300 31282
rect 43456 31226 43484 31776
rect 43364 31198 43484 31226
rect 43260 30592 43312 30598
rect 43260 30534 43312 30540
rect 43168 30320 43220 30326
rect 43168 30262 43220 30268
rect 43364 30190 43392 31198
rect 43536 30796 43588 30802
rect 43536 30738 43588 30744
rect 43548 30598 43576 30738
rect 43628 30728 43680 30734
rect 43628 30670 43680 30676
rect 43444 30592 43496 30598
rect 43444 30534 43496 30540
rect 43536 30592 43588 30598
rect 43536 30534 43588 30540
rect 42248 30184 42300 30190
rect 42248 30126 42300 30132
rect 43352 30184 43404 30190
rect 43352 30126 43404 30132
rect 42260 29850 42288 30126
rect 42064 29844 42116 29850
rect 42064 29786 42116 29792
rect 42248 29844 42300 29850
rect 42248 29786 42300 29792
rect 42800 29844 42852 29850
rect 42800 29786 42852 29792
rect 42076 29730 42104 29786
rect 42076 29702 42288 29730
rect 42812 29714 42840 29786
rect 42260 29646 42288 29702
rect 42800 29708 42852 29714
rect 42800 29650 42852 29656
rect 42248 29640 42300 29646
rect 42248 29582 42300 29588
rect 42812 29170 42840 29650
rect 43364 29510 43392 30126
rect 43456 29850 43484 30534
rect 43640 30190 43668 30670
rect 44744 30190 44772 37062
rect 44928 36174 44956 37198
rect 44916 36168 44968 36174
rect 44916 36110 44968 36116
rect 45204 35698 45232 37198
rect 45192 35692 45244 35698
rect 45192 35634 45244 35640
rect 45572 35222 45600 40326
rect 45756 40118 45784 40326
rect 45744 40112 45796 40118
rect 45744 40054 45796 40060
rect 46032 40050 46060 40326
rect 46020 40044 46072 40050
rect 46020 39986 46072 39992
rect 46032 39642 46060 39986
rect 46020 39636 46072 39642
rect 46020 39578 46072 39584
rect 46584 39438 46612 40326
rect 46860 39982 46888 41976
rect 47676 41958 47728 41964
rect 47688 41750 47716 41958
rect 47676 41744 47728 41750
rect 47676 41686 47728 41692
rect 47400 41676 47452 41682
rect 47400 41618 47452 41624
rect 48780 41676 48832 41682
rect 48780 41618 48832 41624
rect 47412 41070 47440 41618
rect 47400 41064 47452 41070
rect 47400 41006 47452 41012
rect 48228 40996 48280 41002
rect 48228 40938 48280 40944
rect 48136 40928 48188 40934
rect 48136 40870 48188 40876
rect 48148 40118 48176 40870
rect 48136 40112 48188 40118
rect 48136 40054 48188 40060
rect 46848 39976 46900 39982
rect 46848 39918 46900 39924
rect 46860 39846 46888 39918
rect 48240 39914 48268 40938
rect 48792 40934 48820 41618
rect 48780 40928 48832 40934
rect 48780 40870 48832 40876
rect 48872 40520 48924 40526
rect 48872 40462 48924 40468
rect 48780 40112 48832 40118
rect 48780 40054 48832 40060
rect 48228 39908 48280 39914
rect 48228 39850 48280 39856
rect 46848 39840 46900 39846
rect 46848 39782 46900 39788
rect 46940 39840 46992 39846
rect 46940 39782 46992 39788
rect 46572 39432 46624 39438
rect 46572 39374 46624 39380
rect 46112 39024 46164 39030
rect 46164 38972 46428 38978
rect 46112 38966 46428 38972
rect 46124 38962 46428 38966
rect 46124 38956 46440 38962
rect 46124 38950 46388 38956
rect 46388 38898 46440 38904
rect 46584 38894 46612 39374
rect 46572 38888 46624 38894
rect 46572 38830 46624 38836
rect 46860 38758 46888 39782
rect 46952 39642 46980 39782
rect 47582 39672 47638 39681
rect 46940 39636 46992 39642
rect 47582 39607 47638 39616
rect 48044 39636 48096 39642
rect 46940 39578 46992 39584
rect 47596 39506 47624 39607
rect 48044 39578 48096 39584
rect 47032 39500 47084 39506
rect 47032 39442 47084 39448
rect 47400 39500 47452 39506
rect 47400 39442 47452 39448
rect 47584 39500 47636 39506
rect 47584 39442 47636 39448
rect 47044 38894 47072 39442
rect 47306 39400 47362 39409
rect 47306 39335 47362 39344
rect 47320 39302 47348 39335
rect 47412 39302 47440 39442
rect 47308 39296 47360 39302
rect 47308 39238 47360 39244
rect 47400 39296 47452 39302
rect 47400 39238 47452 39244
rect 47860 39296 47912 39302
rect 47860 39238 47912 39244
rect 47032 38888 47084 38894
rect 47032 38830 47084 38836
rect 47124 38888 47176 38894
rect 47124 38830 47176 38836
rect 47136 38758 47164 38830
rect 46848 38752 46900 38758
rect 46848 38694 46900 38700
rect 47124 38752 47176 38758
rect 47124 38694 47176 38700
rect 46020 38344 46072 38350
rect 46020 38286 46072 38292
rect 46032 37738 46060 38286
rect 46572 37800 46624 37806
rect 46572 37742 46624 37748
rect 46020 37732 46072 37738
rect 46020 37674 46072 37680
rect 46204 37664 46256 37670
rect 46204 37606 46256 37612
rect 46216 35630 46244 37606
rect 46584 37398 46612 37742
rect 46662 37496 46718 37505
rect 46662 37431 46718 37440
rect 46676 37398 46704 37431
rect 46572 37392 46624 37398
rect 46572 37334 46624 37340
rect 46664 37392 46716 37398
rect 47136 37380 47164 38694
rect 46664 37334 46716 37340
rect 47044 37352 47164 37380
rect 46756 37120 46808 37126
rect 46756 37062 46808 37068
rect 46768 36718 46796 37062
rect 46756 36712 46808 36718
rect 46756 36654 46808 36660
rect 47044 36106 47072 37352
rect 47872 36922 47900 39238
rect 48056 38962 48084 39578
rect 48792 39574 48820 40054
rect 48884 39574 48912 40462
rect 49528 40390 49556 42026
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 49608 41608 49660 41614
rect 49608 41550 49660 41556
rect 49620 41274 49648 41550
rect 49608 41268 49660 41274
rect 49608 41210 49660 41216
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 49516 40384 49568 40390
rect 49516 40326 49568 40332
rect 49056 39908 49108 39914
rect 49056 39850 49108 39856
rect 48136 39568 48188 39574
rect 48136 39510 48188 39516
rect 48780 39568 48832 39574
rect 48780 39510 48832 39516
rect 48872 39568 48924 39574
rect 48872 39510 48924 39516
rect 48148 39438 48176 39510
rect 48136 39432 48188 39438
rect 49068 39409 49096 39850
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50300 39664 50596 39684
rect 48136 39374 48188 39380
rect 49054 39400 49110 39409
rect 48148 38962 48176 39374
rect 49054 39335 49110 39344
rect 48044 38956 48096 38962
rect 48044 38898 48096 38904
rect 48136 38956 48188 38962
rect 48136 38898 48188 38904
rect 49240 38820 49292 38826
rect 49240 38762 49292 38768
rect 49252 38418 49280 38762
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 49240 38412 49292 38418
rect 49240 38354 49292 38360
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 50724 36922 50752 44134
rect 51276 43858 51304 44270
rect 51264 43852 51316 43858
rect 51264 43794 51316 43800
rect 51264 42900 51316 42906
rect 51264 42842 51316 42848
rect 51276 42702 51304 42842
rect 51264 42696 51316 42702
rect 51264 42638 51316 42644
rect 51172 42560 51224 42566
rect 51092 42520 51172 42548
rect 51092 39982 51120 42520
rect 51172 42502 51224 42508
rect 51172 42016 51224 42022
rect 51172 41958 51224 41964
rect 51264 42016 51316 42022
rect 51264 41958 51316 41964
rect 51080 39976 51132 39982
rect 51080 39918 51132 39924
rect 51184 39001 51212 41958
rect 51276 41818 51304 41958
rect 51264 41812 51316 41818
rect 51264 41754 51316 41760
rect 51170 38992 51226 39001
rect 51170 38927 51226 38936
rect 50988 37392 51040 37398
rect 50986 37360 50988 37369
rect 51040 37360 51042 37369
rect 50986 37295 51042 37304
rect 47860 36916 47912 36922
rect 47860 36858 47912 36864
rect 50712 36916 50764 36922
rect 50712 36858 50764 36864
rect 47872 36310 47900 36858
rect 48136 36848 48188 36854
rect 48136 36790 48188 36796
rect 48148 36310 48176 36790
rect 48504 36576 48556 36582
rect 48504 36518 48556 36524
rect 47860 36304 47912 36310
rect 47860 36246 47912 36252
rect 48136 36304 48188 36310
rect 48136 36246 48188 36252
rect 47032 36100 47084 36106
rect 47032 36042 47084 36048
rect 46756 36032 46808 36038
rect 46756 35974 46808 35980
rect 46768 35698 46796 35974
rect 47044 35766 47072 36042
rect 48516 36038 48544 36518
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 48504 36032 48556 36038
rect 48504 35974 48556 35980
rect 47032 35760 47084 35766
rect 47032 35702 47084 35708
rect 46756 35692 46808 35698
rect 46756 35634 46808 35640
rect 46204 35624 46256 35630
rect 46204 35566 46256 35572
rect 45560 35216 45612 35222
rect 45560 35158 45612 35164
rect 45572 33998 45600 35158
rect 46940 34604 46992 34610
rect 46940 34546 46992 34552
rect 45560 33992 45612 33998
rect 45560 33934 45612 33940
rect 46848 33856 46900 33862
rect 46848 33798 46900 33804
rect 46860 33454 46888 33798
rect 46952 33658 46980 34546
rect 46940 33652 46992 33658
rect 46940 33594 46992 33600
rect 46848 33448 46900 33454
rect 46848 33390 46900 33396
rect 48044 32360 48096 32366
rect 48044 32302 48096 32308
rect 45008 31136 45060 31142
rect 45008 31078 45060 31084
rect 46940 31136 46992 31142
rect 46940 31078 46992 31084
rect 43628 30184 43680 30190
rect 43628 30126 43680 30132
rect 44732 30184 44784 30190
rect 44732 30126 44784 30132
rect 45020 30122 45048 31078
rect 46952 30666 46980 31078
rect 46940 30660 46992 30666
rect 46940 30602 46992 30608
rect 47492 30660 47544 30666
rect 47492 30602 47544 30608
rect 47216 30592 47268 30598
rect 47216 30534 47268 30540
rect 47228 30190 47256 30534
rect 45468 30184 45520 30190
rect 45468 30126 45520 30132
rect 46940 30184 46992 30190
rect 46940 30126 46992 30132
rect 47216 30184 47268 30190
rect 47216 30126 47268 30132
rect 47308 30184 47360 30190
rect 47308 30126 47360 30132
rect 45008 30116 45060 30122
rect 45008 30058 45060 30064
rect 43444 29844 43496 29850
rect 43444 29786 43496 29792
rect 45284 29776 45336 29782
rect 45282 29744 45284 29753
rect 45336 29744 45338 29753
rect 45480 29730 45508 30126
rect 46848 30116 46900 30122
rect 46848 30058 46900 30064
rect 46860 29782 46888 30058
rect 46952 30002 46980 30126
rect 47320 30002 47348 30126
rect 46952 29974 47348 30002
rect 47504 29850 47532 30602
rect 47492 29844 47544 29850
rect 47492 29786 47544 29792
rect 46848 29776 46900 29782
rect 45480 29702 45600 29730
rect 46848 29718 46900 29724
rect 47030 29744 47086 29753
rect 45282 29679 45338 29688
rect 45572 29646 45600 29702
rect 47030 29679 47032 29688
rect 47084 29679 47086 29688
rect 47032 29650 47084 29656
rect 44180 29640 44232 29646
rect 44178 29608 44180 29617
rect 45376 29640 45428 29646
rect 44232 29608 44234 29617
rect 45376 29582 45428 29588
rect 45560 29640 45612 29646
rect 45560 29582 45612 29588
rect 44178 29543 44234 29552
rect 45388 29510 45416 29582
rect 43352 29504 43404 29510
rect 43352 29446 43404 29452
rect 45376 29504 45428 29510
rect 45376 29446 45428 29452
rect 46204 29504 46256 29510
rect 46204 29446 46256 29452
rect 45388 29170 45416 29446
rect 46216 29306 46244 29446
rect 47044 29306 47072 29650
rect 48056 29578 48084 32302
rect 48516 32230 48544 35974
rect 49700 35556 49752 35562
rect 49700 35498 49752 35504
rect 49148 34740 49200 34746
rect 49148 34682 49200 34688
rect 49160 33046 49188 34682
rect 49712 34542 49740 35498
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 49700 34536 49752 34542
rect 49700 34478 49752 34484
rect 49240 33924 49292 33930
rect 49240 33866 49292 33872
rect 49252 33658 49280 33866
rect 49240 33652 49292 33658
rect 49240 33594 49292 33600
rect 49252 33522 49280 33594
rect 49240 33516 49292 33522
rect 49240 33458 49292 33464
rect 49148 33040 49200 33046
rect 49148 32982 49200 32988
rect 49712 32978 49740 34478
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 50724 34066 50752 36858
rect 51368 36854 51396 46310
rect 51736 46050 51764 46854
rect 51644 46034 51764 46050
rect 51920 46322 51948 47058
rect 52368 46912 52420 46918
rect 52368 46854 52420 46860
rect 52000 46368 52052 46374
rect 51920 46316 52000 46322
rect 51920 46310 52052 46316
rect 51920 46294 52040 46310
rect 51632 46028 51776 46034
rect 51684 46022 51724 46028
rect 51632 45970 51684 45976
rect 51724 45970 51776 45976
rect 51920 45422 51948 46294
rect 51908 45416 51960 45422
rect 51908 45358 51960 45364
rect 52380 45370 52408 46854
rect 52644 45824 52696 45830
rect 52644 45766 52696 45772
rect 52460 45416 52512 45422
rect 52380 45364 52460 45370
rect 52380 45358 52512 45364
rect 52380 45342 52500 45358
rect 51908 45280 51960 45286
rect 51908 45222 51960 45228
rect 51724 44804 51776 44810
rect 51724 44746 51776 44752
rect 51736 44402 51764 44746
rect 51724 44396 51776 44402
rect 51724 44338 51776 44344
rect 51920 44334 51948 45222
rect 52656 44878 52684 45766
rect 54496 45626 54524 49248
rect 73068 48340 73120 48346
rect 73068 48282 73120 48288
rect 65660 47900 65956 47920
rect 65716 47898 65740 47900
rect 65796 47898 65820 47900
rect 65876 47898 65900 47900
rect 65738 47846 65740 47898
rect 65802 47846 65814 47898
rect 65876 47846 65878 47898
rect 65716 47844 65740 47846
rect 65796 47844 65820 47846
rect 65876 47844 65900 47846
rect 65660 47824 65956 47844
rect 56692 47116 56744 47122
rect 56692 47058 56744 47064
rect 56784 47116 56836 47122
rect 56784 47058 56836 47064
rect 62948 47116 63000 47122
rect 62948 47058 63000 47064
rect 56704 46578 56732 47058
rect 56692 46572 56744 46578
rect 56692 46514 56744 46520
rect 54852 46504 54904 46510
rect 54852 46446 54904 46452
rect 54864 46102 54892 46446
rect 56600 46368 56652 46374
rect 56600 46310 56652 46316
rect 54852 46096 54904 46102
rect 54852 46038 54904 46044
rect 55956 46028 56008 46034
rect 55956 45970 56008 45976
rect 54484 45620 54536 45626
rect 54484 45562 54536 45568
rect 55128 45620 55180 45626
rect 55128 45562 55180 45568
rect 54944 45348 54996 45354
rect 54944 45290 54996 45296
rect 52644 44872 52696 44878
rect 52644 44814 52696 44820
rect 52460 44736 52512 44742
rect 52460 44678 52512 44684
rect 52552 44736 52604 44742
rect 52552 44678 52604 44684
rect 54576 44736 54628 44742
rect 54576 44678 54628 44684
rect 51908 44328 51960 44334
rect 51908 44270 51960 44276
rect 52472 43926 52500 44678
rect 52460 43920 52512 43926
rect 52460 43862 52512 43868
rect 51908 43852 51960 43858
rect 51908 43794 51960 43800
rect 51448 43240 51500 43246
rect 51448 43182 51500 43188
rect 51460 43110 51488 43182
rect 51448 43104 51500 43110
rect 51448 43046 51500 43052
rect 51460 42090 51488 43046
rect 51816 42900 51868 42906
rect 51816 42842 51868 42848
rect 51724 42764 51776 42770
rect 51724 42706 51776 42712
rect 51736 42634 51764 42706
rect 51724 42628 51776 42634
rect 51724 42570 51776 42576
rect 51448 42084 51500 42090
rect 51448 42026 51500 42032
rect 51828 41478 51856 42842
rect 51816 41472 51868 41478
rect 51816 41414 51868 41420
rect 51828 39506 51856 41414
rect 51816 39500 51868 39506
rect 51816 39442 51868 39448
rect 51724 39432 51776 39438
rect 51724 39374 51776 39380
rect 51736 39302 51764 39374
rect 51724 39296 51776 39302
rect 51724 39238 51776 39244
rect 51448 38820 51500 38826
rect 51448 38762 51500 38768
rect 51460 37942 51488 38762
rect 51736 38010 51764 39238
rect 51816 38548 51868 38554
rect 51816 38490 51868 38496
rect 51724 38004 51776 38010
rect 51724 37946 51776 37952
rect 51448 37936 51500 37942
rect 51448 37878 51500 37884
rect 51828 37330 51856 38490
rect 51816 37324 51868 37330
rect 51816 37266 51868 37272
rect 51356 36848 51408 36854
rect 51356 36790 51408 36796
rect 51724 36848 51776 36854
rect 51724 36790 51776 36796
rect 50804 36780 50856 36786
rect 50804 36722 50856 36728
rect 50160 34060 50212 34066
rect 50160 34002 50212 34008
rect 50712 34060 50764 34066
rect 50712 34002 50764 34008
rect 49700 32972 49752 32978
rect 49700 32914 49752 32920
rect 50172 32910 50200 34002
rect 50816 33658 50844 36722
rect 51368 36242 51396 36790
rect 51736 36718 51764 36790
rect 51724 36712 51776 36718
rect 51724 36654 51776 36660
rect 51356 36236 51408 36242
rect 51356 36178 51408 36184
rect 50988 36168 51040 36174
rect 50988 36110 51040 36116
rect 51000 34134 51028 36110
rect 51920 35766 51948 43794
rect 52460 43716 52512 43722
rect 52460 43658 52512 43664
rect 52000 43240 52052 43246
rect 52000 43182 52052 43188
rect 52012 42906 52040 43182
rect 52000 42900 52052 42906
rect 52000 42842 52052 42848
rect 52184 42764 52236 42770
rect 52184 42706 52236 42712
rect 52196 42634 52224 42706
rect 52184 42628 52236 42634
rect 52184 42570 52236 42576
rect 52276 42560 52328 42566
rect 52276 42502 52328 42508
rect 52472 42514 52500 43658
rect 52564 42634 52592 44678
rect 52828 44464 52880 44470
rect 52828 44406 52880 44412
rect 52840 43926 52868 44406
rect 53288 44192 53340 44198
rect 53288 44134 53340 44140
rect 52828 43920 52880 43926
rect 52828 43862 52880 43868
rect 53300 43722 53328 44134
rect 54116 43988 54168 43994
rect 54116 43930 54168 43936
rect 53288 43716 53340 43722
rect 53288 43658 53340 43664
rect 52920 43648 52972 43654
rect 52920 43590 52972 43596
rect 52932 43450 52960 43590
rect 52920 43444 52972 43450
rect 52920 43386 52972 43392
rect 53196 43444 53248 43450
rect 53196 43386 53248 43392
rect 53012 43308 53064 43314
rect 53012 43250 53064 43256
rect 53024 42906 53052 43250
rect 53208 43246 53236 43386
rect 53196 43240 53248 43246
rect 53196 43182 53248 43188
rect 53208 42906 53236 43182
rect 53012 42900 53064 42906
rect 53012 42842 53064 42848
rect 53196 42900 53248 42906
rect 53196 42842 53248 42848
rect 52552 42628 52604 42634
rect 52552 42570 52604 42576
rect 52288 42158 52316 42502
rect 52472 42486 52684 42514
rect 52276 42152 52328 42158
rect 52276 42094 52328 42100
rect 52288 41682 52316 42094
rect 52276 41676 52328 41682
rect 52276 41618 52328 41624
rect 52552 41676 52604 41682
rect 52552 41618 52604 41624
rect 52564 41478 52592 41618
rect 52552 41472 52604 41478
rect 52552 41414 52604 41420
rect 52460 40588 52512 40594
rect 52460 40530 52512 40536
rect 52472 40050 52500 40530
rect 52460 40044 52512 40050
rect 52460 39986 52512 39992
rect 52276 39500 52328 39506
rect 52276 39442 52328 39448
rect 52288 39302 52316 39442
rect 52276 39296 52328 39302
rect 52276 39238 52328 39244
rect 52288 38894 52316 39238
rect 52276 38888 52328 38894
rect 52276 38830 52328 38836
rect 52656 38418 52684 42486
rect 53024 42362 53052 42842
rect 53012 42356 53064 42362
rect 53012 42298 53064 42304
rect 53472 42356 53524 42362
rect 53472 42298 53524 42304
rect 53024 42226 53052 42298
rect 53012 42220 53064 42226
rect 53012 42162 53064 42168
rect 53012 42084 53064 42090
rect 53012 42026 53064 42032
rect 52748 40718 52960 40746
rect 52748 40662 52776 40718
rect 52736 40656 52788 40662
rect 52736 40598 52788 40604
rect 52828 40656 52880 40662
rect 52828 40598 52880 40604
rect 52840 40526 52868 40598
rect 52932 40594 52960 40718
rect 52920 40588 52972 40594
rect 52920 40530 52972 40536
rect 53024 40526 53052 42026
rect 53484 41818 53512 42298
rect 53472 41812 53524 41818
rect 53392 41772 53472 41800
rect 53392 41682 53420 41772
rect 53472 41754 53524 41760
rect 53380 41676 53432 41682
rect 53380 41618 53432 41624
rect 53472 41608 53524 41614
rect 53472 41550 53524 41556
rect 53484 41138 53512 41550
rect 53196 41132 53248 41138
rect 53196 41074 53248 41080
rect 53472 41132 53524 41138
rect 53472 41074 53524 41080
rect 52828 40520 52880 40526
rect 52828 40462 52880 40468
rect 53012 40520 53064 40526
rect 53012 40462 53064 40468
rect 53104 40520 53156 40526
rect 53104 40462 53156 40468
rect 53116 40118 53144 40462
rect 53104 40112 53156 40118
rect 53104 40054 53156 40060
rect 52828 39500 52880 39506
rect 52828 39442 52880 39448
rect 52840 39302 52868 39442
rect 52828 39296 52880 39302
rect 52828 39238 52880 39244
rect 53104 39092 53156 39098
rect 53104 39034 53156 39040
rect 53116 38826 53144 39034
rect 53104 38820 53156 38826
rect 53104 38762 53156 38768
rect 52736 38752 52788 38758
rect 52736 38694 52788 38700
rect 52644 38412 52696 38418
rect 52644 38354 52696 38360
rect 52368 38344 52420 38350
rect 52368 38286 52420 38292
rect 52380 37942 52408 38286
rect 52748 38282 52776 38694
rect 53104 38344 53156 38350
rect 53104 38286 53156 38292
rect 52736 38276 52788 38282
rect 52736 38218 52788 38224
rect 52368 37936 52420 37942
rect 52368 37878 52420 37884
rect 52000 37800 52052 37806
rect 52000 37742 52052 37748
rect 52368 37800 52420 37806
rect 52368 37742 52420 37748
rect 52552 37800 52604 37806
rect 52552 37742 52604 37748
rect 52012 37670 52040 37742
rect 52000 37664 52052 37670
rect 52000 37606 52052 37612
rect 52012 37330 52040 37606
rect 52000 37324 52052 37330
rect 52000 37266 52052 37272
rect 52380 36582 52408 37742
rect 52564 37330 52592 37742
rect 53116 37398 53144 38286
rect 53104 37392 53156 37398
rect 53104 37334 53156 37340
rect 52552 37324 52604 37330
rect 52552 37266 52604 37272
rect 53104 37256 53156 37262
rect 53104 37198 53156 37204
rect 53116 36582 53144 37198
rect 52368 36576 52420 36582
rect 52368 36518 52420 36524
rect 53104 36576 53156 36582
rect 53104 36518 53156 36524
rect 53208 36530 53236 41074
rect 53932 40384 53984 40390
rect 53932 40326 53984 40332
rect 53944 39982 53972 40326
rect 54128 40118 54156 43930
rect 54484 40928 54536 40934
rect 54484 40870 54536 40876
rect 54300 40452 54352 40458
rect 54300 40394 54352 40400
rect 54116 40112 54168 40118
rect 54116 40054 54168 40060
rect 53380 39976 53432 39982
rect 53380 39918 53432 39924
rect 53932 39976 53984 39982
rect 54208 39976 54260 39982
rect 53932 39918 53984 39924
rect 54206 39944 54208 39953
rect 54260 39944 54262 39953
rect 53288 39296 53340 39302
rect 53288 39238 53340 39244
rect 53300 39098 53328 39238
rect 53288 39092 53340 39098
rect 53288 39034 53340 39040
rect 53392 39030 53420 39918
rect 54206 39879 54262 39888
rect 53656 39432 53708 39438
rect 53656 39374 53708 39380
rect 53380 39024 53432 39030
rect 53380 38966 53432 38972
rect 53668 38894 53696 39374
rect 54208 39364 54260 39370
rect 54208 39306 54260 39312
rect 54220 38894 54248 39306
rect 53656 38888 53708 38894
rect 53656 38830 53708 38836
rect 54208 38888 54260 38894
rect 54208 38830 54260 38836
rect 53380 37868 53432 37874
rect 53380 37810 53432 37816
rect 53392 37398 53420 37810
rect 53564 37800 53616 37806
rect 53564 37742 53616 37748
rect 53576 37670 53604 37742
rect 53564 37664 53616 37670
rect 53564 37606 53616 37612
rect 53576 37398 53604 37606
rect 53380 37392 53432 37398
rect 53380 37334 53432 37340
rect 53564 37392 53616 37398
rect 53564 37334 53616 37340
rect 52380 36310 52408 36518
rect 52368 36304 52420 36310
rect 52368 36246 52420 36252
rect 51172 35760 51224 35766
rect 51172 35702 51224 35708
rect 51908 35760 51960 35766
rect 51908 35702 51960 35708
rect 50988 34128 51040 34134
rect 50988 34070 51040 34076
rect 50804 33652 50856 33658
rect 50804 33594 50856 33600
rect 50988 33652 51040 33658
rect 50988 33594 51040 33600
rect 50300 33212 50596 33232
rect 50356 33210 50380 33212
rect 50436 33210 50460 33212
rect 50516 33210 50540 33212
rect 50378 33158 50380 33210
rect 50442 33158 50454 33210
rect 50516 33158 50518 33210
rect 50356 33156 50380 33158
rect 50436 33156 50460 33158
rect 50516 33156 50540 33158
rect 50300 33136 50596 33156
rect 51000 32910 51028 33594
rect 51184 33454 51212 35702
rect 53116 35630 53144 36518
rect 53208 36502 53328 36530
rect 53104 35624 53156 35630
rect 53104 35566 53156 35572
rect 52552 35148 52604 35154
rect 52552 35090 52604 35096
rect 51448 34740 51500 34746
rect 51448 34682 51500 34688
rect 51172 33448 51224 33454
rect 51172 33390 51224 33396
rect 51184 32978 51212 33390
rect 51460 33386 51488 34682
rect 52564 34678 52592 35090
rect 52552 34672 52604 34678
rect 52552 34614 52604 34620
rect 52828 34536 52880 34542
rect 52828 34478 52880 34484
rect 52840 33454 52868 34478
rect 52828 33448 52880 33454
rect 51814 33416 51870 33425
rect 51448 33380 51500 33386
rect 52828 33390 52880 33396
rect 53012 33448 53064 33454
rect 53012 33390 53064 33396
rect 51814 33351 51816 33360
rect 51448 33322 51500 33328
rect 51868 33351 51870 33360
rect 51816 33322 51868 33328
rect 51460 33046 51488 33322
rect 53024 33318 53052 33390
rect 53012 33312 53064 33318
rect 53012 33254 53064 33260
rect 51448 33040 51500 33046
rect 51448 32982 51500 32988
rect 51172 32972 51224 32978
rect 51172 32914 51224 32920
rect 50160 32904 50212 32910
rect 50160 32846 50212 32852
rect 50988 32904 51040 32910
rect 50988 32846 51040 32852
rect 48504 32224 48556 32230
rect 48504 32166 48556 32172
rect 48320 31816 48372 31822
rect 48320 31758 48372 31764
rect 48134 30696 48190 30705
rect 48134 30631 48190 30640
rect 48148 29578 48176 30631
rect 48332 30054 48360 31758
rect 48516 30734 48544 32166
rect 50300 32124 50596 32144
rect 50356 32122 50380 32124
rect 50436 32122 50460 32124
rect 50516 32122 50540 32124
rect 50378 32070 50380 32122
rect 50442 32070 50454 32122
rect 50516 32070 50518 32122
rect 50356 32068 50380 32070
rect 50436 32068 50460 32070
rect 50516 32068 50540 32070
rect 50300 32048 50596 32068
rect 52368 32020 52420 32026
rect 52368 31962 52420 31968
rect 50160 31680 50212 31686
rect 50160 31622 50212 31628
rect 49240 31204 49292 31210
rect 49240 31146 49292 31152
rect 49252 30802 49280 31146
rect 49240 30796 49292 30802
rect 49240 30738 49292 30744
rect 48504 30728 48556 30734
rect 48504 30670 48556 30676
rect 50172 30598 50200 31622
rect 52380 31278 52408 31962
rect 53196 31884 53248 31890
rect 53196 31826 53248 31832
rect 53208 31686 53236 31826
rect 53196 31680 53248 31686
rect 53196 31622 53248 31628
rect 52368 31272 52420 31278
rect 52368 31214 52420 31220
rect 53300 31142 53328 36502
rect 53380 32904 53432 32910
rect 53380 32846 53432 32852
rect 53392 31890 53420 32846
rect 53484 32694 53696 32722
rect 53484 32366 53512 32694
rect 53668 32570 53696 32694
rect 53564 32564 53616 32570
rect 53564 32506 53616 32512
rect 53656 32564 53708 32570
rect 53656 32506 53708 32512
rect 53472 32360 53524 32366
rect 53472 32302 53524 32308
rect 53380 31884 53432 31890
rect 53380 31826 53432 31832
rect 53288 31136 53340 31142
rect 53288 31078 53340 31084
rect 50300 31036 50596 31056
rect 50356 31034 50380 31036
rect 50436 31034 50460 31036
rect 50516 31034 50540 31036
rect 50378 30982 50380 31034
rect 50442 30982 50454 31034
rect 50516 30982 50518 31034
rect 50356 30980 50380 30982
rect 50436 30980 50460 30982
rect 50516 30980 50540 30982
rect 50300 30960 50596 30980
rect 48780 30592 48832 30598
rect 48780 30534 48832 30540
rect 50160 30592 50212 30598
rect 50160 30534 50212 30540
rect 48792 30326 48820 30534
rect 48780 30320 48832 30326
rect 48780 30262 48832 30268
rect 48792 30190 48820 30262
rect 48780 30184 48832 30190
rect 48780 30126 48832 30132
rect 48320 30048 48372 30054
rect 48320 29990 48372 29996
rect 48044 29572 48096 29578
rect 48044 29514 48096 29520
rect 48136 29572 48188 29578
rect 48136 29514 48188 29520
rect 46204 29300 46256 29306
rect 46204 29242 46256 29248
rect 47032 29300 47084 29306
rect 47032 29242 47084 29248
rect 42800 29164 42852 29170
rect 42800 29106 42852 29112
rect 45376 29164 45428 29170
rect 45376 29106 45428 29112
rect 48332 28150 48360 29990
rect 48962 29608 49018 29617
rect 48962 29543 49018 29552
rect 48976 29510 49004 29543
rect 48872 29504 48924 29510
rect 48870 29472 48872 29481
rect 48964 29504 49016 29510
rect 48924 29472 48926 29481
rect 48964 29446 49016 29452
rect 48870 29407 48926 29416
rect 48320 28144 48372 28150
rect 48320 28086 48372 28092
rect 50172 27402 50200 30534
rect 52656 30258 53328 30274
rect 52644 30252 53328 30258
rect 52696 30246 53328 30252
rect 52644 30194 52696 30200
rect 53300 30190 53328 30246
rect 53012 30184 53064 30190
rect 53012 30126 53064 30132
rect 53288 30184 53340 30190
rect 53288 30126 53340 30132
rect 52000 30048 52052 30054
rect 52000 29990 52052 29996
rect 50300 29948 50596 29968
rect 50356 29946 50380 29948
rect 50436 29946 50460 29948
rect 50516 29946 50540 29948
rect 50378 29894 50380 29946
rect 50442 29894 50454 29946
rect 50516 29894 50518 29946
rect 50356 29892 50380 29894
rect 50436 29892 50460 29894
rect 50516 29892 50540 29894
rect 50300 29872 50596 29892
rect 50988 29708 51040 29714
rect 50988 29650 51040 29656
rect 51000 29034 51028 29650
rect 52012 29646 52040 29990
rect 53024 29850 53052 30126
rect 52644 29844 52696 29850
rect 52644 29786 52696 29792
rect 53012 29844 53064 29850
rect 53012 29786 53064 29792
rect 52000 29640 52052 29646
rect 52000 29582 52052 29588
rect 52012 29238 52040 29582
rect 52656 29238 52684 29786
rect 52748 29714 53144 29730
rect 52736 29708 53156 29714
rect 52788 29702 53104 29708
rect 52736 29650 52788 29656
rect 53104 29650 53156 29656
rect 53196 29640 53248 29646
rect 53196 29582 53248 29588
rect 53208 29481 53236 29582
rect 53576 29510 53604 32506
rect 53668 31822 53696 32506
rect 54312 32434 54340 40394
rect 54392 40112 54444 40118
rect 54392 40054 54444 40060
rect 54404 39914 54432 40054
rect 54392 39908 54444 39914
rect 54392 39850 54444 39856
rect 54496 39574 54524 40870
rect 54392 39568 54444 39574
rect 54392 39510 54444 39516
rect 54484 39568 54536 39574
rect 54484 39510 54536 39516
rect 54404 38758 54432 39510
rect 54588 39370 54616 44678
rect 54668 44260 54720 44266
rect 54668 44202 54720 44208
rect 54680 43858 54708 44202
rect 54668 43852 54720 43858
rect 54668 43794 54720 43800
rect 54956 43790 54984 45290
rect 54944 43784 54996 43790
rect 54944 43726 54996 43732
rect 54852 40112 54904 40118
rect 54852 40054 54904 40060
rect 54668 40044 54720 40050
rect 54668 39986 54720 39992
rect 54576 39364 54628 39370
rect 54576 39306 54628 39312
rect 54680 39098 54708 39986
rect 54864 39953 54892 40054
rect 54850 39944 54906 39953
rect 54850 39879 54906 39888
rect 54864 39506 54892 39879
rect 54852 39500 54904 39506
rect 54852 39442 54904 39448
rect 54944 39432 54996 39438
rect 54944 39374 54996 39380
rect 54668 39092 54720 39098
rect 54668 39034 54720 39040
rect 54576 38956 54628 38962
rect 54576 38898 54628 38904
rect 54392 38752 54444 38758
rect 54392 38694 54444 38700
rect 54588 38010 54616 38898
rect 54956 38554 54984 39374
rect 54944 38548 54996 38554
rect 54944 38490 54996 38496
rect 55036 38548 55088 38554
rect 55036 38490 55088 38496
rect 54576 38004 54628 38010
rect 54576 37946 54628 37952
rect 55048 37806 55076 38490
rect 55036 37800 55088 37806
rect 55036 37742 55088 37748
rect 54576 34400 54628 34406
rect 54576 34342 54628 34348
rect 54588 33998 54616 34342
rect 54576 33992 54628 33998
rect 54576 33934 54628 33940
rect 54588 33658 54616 33934
rect 54576 33652 54628 33658
rect 54576 33594 54628 33600
rect 54588 33454 54616 33594
rect 54576 33448 54628 33454
rect 54576 33390 54628 33396
rect 54300 32428 54352 32434
rect 54300 32370 54352 32376
rect 54852 32428 54904 32434
rect 54852 32370 54904 32376
rect 53748 32360 53800 32366
rect 53748 32302 53800 32308
rect 53760 32026 53788 32302
rect 54864 32026 54892 32370
rect 55036 32360 55088 32366
rect 55036 32302 55088 32308
rect 55048 32230 55076 32302
rect 55036 32224 55088 32230
rect 55036 32166 55088 32172
rect 55048 32026 55076 32166
rect 53748 32020 53800 32026
rect 53748 31962 53800 31968
rect 54852 32020 54904 32026
rect 54852 31962 54904 31968
rect 55036 32020 55088 32026
rect 55036 31962 55088 31968
rect 53656 31816 53708 31822
rect 53656 31758 53708 31764
rect 53668 31278 53696 31758
rect 54944 31748 54996 31754
rect 54944 31690 54996 31696
rect 54116 31680 54168 31686
rect 54116 31622 54168 31628
rect 54128 31278 54156 31622
rect 54956 31346 54984 31690
rect 54944 31340 54996 31346
rect 54944 31282 54996 31288
rect 55048 31278 55076 31962
rect 53656 31272 53708 31278
rect 53656 31214 53708 31220
rect 53840 31272 53892 31278
rect 54116 31272 54168 31278
rect 53892 31232 54064 31260
rect 53840 31214 53892 31220
rect 54036 30802 54064 31232
rect 54116 31214 54168 31220
rect 55036 31272 55088 31278
rect 55036 31214 55088 31220
rect 54024 30796 54076 30802
rect 54024 30738 54076 30744
rect 54036 30394 54064 30738
rect 54128 30734 54156 31214
rect 54116 30728 54168 30734
rect 54116 30670 54168 30676
rect 54668 30592 54720 30598
rect 54668 30534 54720 30540
rect 54024 30388 54076 30394
rect 54024 30330 54076 30336
rect 54680 29646 54708 30534
rect 54668 29640 54720 29646
rect 54668 29582 54720 29588
rect 53564 29504 53616 29510
rect 53194 29472 53250 29481
rect 53564 29446 53616 29452
rect 53194 29407 53250 29416
rect 52000 29232 52052 29238
rect 52000 29174 52052 29180
rect 52644 29232 52696 29238
rect 52644 29174 52696 29180
rect 50988 29028 51040 29034
rect 50988 28970 51040 28976
rect 53576 28966 53604 29446
rect 53840 29164 53892 29170
rect 53840 29106 53892 29112
rect 53564 28960 53616 28966
rect 53564 28902 53616 28908
rect 50160 27396 50212 27402
rect 50160 27338 50212 27344
rect 41880 27124 41932 27130
rect 41880 27066 41932 27072
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 31574 22834 31630 22843
rect 31574 22769 31630 22778
rect 31588 22234 31616 22769
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 28998 21720 29054 21729
rect 28998 21655 29054 21664
rect 29012 20806 29040 21655
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 28998 20632 29054 20641
rect 28998 20567 29054 20576
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 29012 19922 29040 20567
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28906 19544 28962 19553
rect 28906 19479 28962 19488
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27724 18970 27752 19246
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 27264 18630 27292 18770
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 27264 17066 27292 18566
rect 28920 17746 28948 19479
rect 28080 17740 28132 17746
rect 28080 17682 28132 17688
rect 28908 17740 28960 17746
rect 28908 17682 28960 17688
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27356 17134 27384 17478
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16658 26832 16934
rect 28092 16794 28120 17682
rect 28906 17368 28962 17377
rect 28906 17303 28962 17312
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 28920 16250 28948 17303
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 26528 15570 26556 16186
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 26792 13728 26844 13734
rect 26792 13670 26844 13676
rect 26804 13394 26832 13670
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 27816 13190 27844 13806
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 31760 13184 31812 13190
rect 31760 13126 31812 13132
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26436 10674 26464 11494
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26792 10464 26844 10470
rect 26792 10406 26844 10412
rect 26804 10130 26832 10406
rect 27632 10266 27660 13126
rect 31772 13095 31800 13126
rect 31758 13086 31814 13095
rect 31758 13021 31814 13030
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 25596 5296 25648 5302
rect 25596 5238 25648 5244
rect 29920 5092 29972 5098
rect 29920 5034 29972 5040
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 29932 4865 29960 5034
rect 29918 4856 29974 4865
rect 12072 4820 12124 4826
rect 29918 4791 29974 4800
rect 12072 4762 12124 4768
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 3738 11100 4422
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 53852 898 53880 29106
rect 55140 26246 55168 45562
rect 55864 45348 55916 45354
rect 55864 45290 55916 45296
rect 55876 44946 55904 45290
rect 55968 45286 55996 45970
rect 56612 45422 56640 46310
rect 56796 46102 56824 47058
rect 57244 47048 57296 47054
rect 57244 46990 57296 46996
rect 61476 47048 61528 47054
rect 61476 46990 61528 46996
rect 57256 46578 57284 46990
rect 59544 46980 59596 46986
rect 59544 46922 59596 46928
rect 57244 46572 57296 46578
rect 57244 46514 57296 46520
rect 57336 46504 57388 46510
rect 57336 46446 57388 46452
rect 57428 46504 57480 46510
rect 57428 46446 57480 46452
rect 56784 46096 56836 46102
rect 56784 46038 56836 46044
rect 56600 45416 56652 45422
rect 56600 45358 56652 45364
rect 56612 45286 56640 45358
rect 55956 45280 56008 45286
rect 55956 45222 56008 45228
rect 56600 45280 56652 45286
rect 56600 45222 56652 45228
rect 55864 44940 55916 44946
rect 55864 44882 55916 44888
rect 57348 44878 57376 46446
rect 57440 46170 57468 46446
rect 59176 46368 59228 46374
rect 59176 46310 59228 46316
rect 57428 46164 57480 46170
rect 57428 46106 57480 46112
rect 58532 45416 58584 45422
rect 58532 45358 58584 45364
rect 57520 45280 57572 45286
rect 57520 45222 57572 45228
rect 57704 45280 57756 45286
rect 57704 45222 57756 45228
rect 57336 44872 57388 44878
rect 57336 44814 57388 44820
rect 57244 44804 57296 44810
rect 57244 44746 57296 44752
rect 56784 44532 56836 44538
rect 56784 44474 56836 44480
rect 56600 43376 56652 43382
rect 56600 43318 56652 43324
rect 55864 41268 55916 41274
rect 55864 41210 55916 41216
rect 55876 40730 55904 41210
rect 55864 40724 55916 40730
rect 55864 40666 55916 40672
rect 56508 39840 56560 39846
rect 56508 39782 56560 39788
rect 55220 39568 55272 39574
rect 55220 39510 55272 39516
rect 55232 39438 55260 39510
rect 55220 39432 55272 39438
rect 55220 39374 55272 39380
rect 55312 38208 55364 38214
rect 55312 38150 55364 38156
rect 55324 37369 55352 38150
rect 56520 37738 56548 39782
rect 56508 37732 56560 37738
rect 56508 37674 56560 37680
rect 55310 37360 55366 37369
rect 55310 37295 55366 37304
rect 55220 35216 55272 35222
rect 55218 35184 55220 35193
rect 55272 35184 55274 35193
rect 55218 35119 55274 35128
rect 55324 29578 55352 37295
rect 56612 35562 56640 43318
rect 56600 35556 56652 35562
rect 56600 35498 56652 35504
rect 56598 35320 56654 35329
rect 56598 35255 56600 35264
rect 56652 35255 56654 35264
rect 56600 35226 56652 35232
rect 56048 34400 56100 34406
rect 56048 34342 56100 34348
rect 56060 34066 56088 34342
rect 56796 34134 56824 44474
rect 57256 44402 57284 44746
rect 57244 44396 57296 44402
rect 57244 44338 57296 44344
rect 56968 36168 57020 36174
rect 56968 36110 57020 36116
rect 56876 35556 56928 35562
rect 56876 35498 56928 35504
rect 56784 34128 56836 34134
rect 56784 34070 56836 34076
rect 55496 34060 55548 34066
rect 55496 34002 55548 34008
rect 56048 34060 56100 34066
rect 56048 34002 56100 34008
rect 55508 33590 55536 34002
rect 56692 33992 56744 33998
rect 56692 33934 56744 33940
rect 55496 33584 55548 33590
rect 55496 33526 55548 33532
rect 55864 32972 55916 32978
rect 55864 32914 55916 32920
rect 55876 32298 55904 32914
rect 56704 32910 56732 33934
rect 56888 33658 56916 35498
rect 56980 35329 57008 36110
rect 57060 35692 57112 35698
rect 57060 35634 57112 35640
rect 56966 35320 57022 35329
rect 56966 35255 57022 35264
rect 56968 35148 57020 35154
rect 56968 35090 57020 35096
rect 56980 34746 57008 35090
rect 57072 34746 57100 35634
rect 56968 34740 57020 34746
rect 56968 34682 57020 34688
rect 57060 34740 57112 34746
rect 57060 34682 57112 34688
rect 57532 34066 57560 45222
rect 57716 44946 57744 45222
rect 57704 44940 57756 44946
rect 57704 44882 57756 44888
rect 58544 44538 58572 45358
rect 59188 44878 59216 46310
rect 59176 44872 59228 44878
rect 59176 44814 59228 44820
rect 59084 44736 59136 44742
rect 59084 44678 59136 44684
rect 58532 44532 58584 44538
rect 58532 44474 58584 44480
rect 59096 43926 59124 44678
rect 59176 44328 59228 44334
rect 59176 44270 59228 44276
rect 59452 44328 59504 44334
rect 59452 44270 59504 44276
rect 59084 43920 59136 43926
rect 59084 43862 59136 43868
rect 59096 43450 59124 43862
rect 59084 43444 59136 43450
rect 59084 43386 59136 43392
rect 58714 43344 58770 43353
rect 58714 43279 58716 43288
rect 58768 43279 58770 43288
rect 58716 43250 58768 43256
rect 59188 43110 59216 44270
rect 59464 43994 59492 44270
rect 59452 43988 59504 43994
rect 59452 43930 59504 43936
rect 59556 43602 59584 46922
rect 61488 46102 61516 46990
rect 62960 46918 62988 47058
rect 62120 46912 62172 46918
rect 62120 46854 62172 46860
rect 62948 46912 63000 46918
rect 62948 46854 63000 46860
rect 62132 46714 62160 46854
rect 62120 46708 62172 46714
rect 62120 46650 62172 46656
rect 62132 46510 62160 46650
rect 62120 46504 62172 46510
rect 62120 46446 62172 46452
rect 62028 46368 62080 46374
rect 62028 46310 62080 46316
rect 61476 46096 61528 46102
rect 61476 46038 61528 46044
rect 62040 45898 62068 46310
rect 62304 45960 62356 45966
rect 62304 45902 62356 45908
rect 62028 45892 62080 45898
rect 62028 45834 62080 45840
rect 60924 45076 60976 45082
rect 60924 45018 60976 45024
rect 60372 44940 60424 44946
rect 60372 44882 60424 44888
rect 60188 44260 60240 44266
rect 60188 44202 60240 44208
rect 60200 43858 60228 44202
rect 60384 43994 60412 44882
rect 60740 44872 60792 44878
rect 60740 44814 60792 44820
rect 60464 44736 60516 44742
rect 60464 44678 60516 44684
rect 60476 44538 60504 44678
rect 60752 44538 60780 44814
rect 60936 44538 60964 45018
rect 61568 45008 61620 45014
rect 61568 44950 61620 44956
rect 60464 44532 60516 44538
rect 60464 44474 60516 44480
rect 60740 44532 60792 44538
rect 60740 44474 60792 44480
rect 60924 44532 60976 44538
rect 60924 44474 60976 44480
rect 60740 44396 60792 44402
rect 60740 44338 60792 44344
rect 60372 43988 60424 43994
rect 60372 43930 60424 43936
rect 60464 43988 60516 43994
rect 60464 43930 60516 43936
rect 60188 43852 60240 43858
rect 60188 43794 60240 43800
rect 60004 43716 60056 43722
rect 60004 43658 60056 43664
rect 59464 43574 59584 43602
rect 59464 43246 59492 43574
rect 59544 43444 59596 43450
rect 59544 43386 59596 43392
rect 59452 43240 59504 43246
rect 59452 43182 59504 43188
rect 59176 43104 59228 43110
rect 59176 43046 59228 43052
rect 59464 42770 59492 43182
rect 58900 42764 58952 42770
rect 58900 42706 58952 42712
rect 59452 42764 59504 42770
rect 59452 42706 59504 42712
rect 58808 42560 58860 42566
rect 58808 42502 58860 42508
rect 58164 42288 58216 42294
rect 58164 42230 58216 42236
rect 58176 41682 58204 42230
rect 58820 42226 58848 42502
rect 58912 42362 58940 42706
rect 58900 42356 58952 42362
rect 58900 42298 58952 42304
rect 59268 42288 59320 42294
rect 59268 42230 59320 42236
rect 58808 42220 58860 42226
rect 58808 42162 58860 42168
rect 59280 42158 59308 42230
rect 59268 42152 59320 42158
rect 59268 42094 59320 42100
rect 58440 42016 58492 42022
rect 58440 41958 58492 41964
rect 58164 41676 58216 41682
rect 58164 41618 58216 41624
rect 58452 40730 58480 41958
rect 59176 41200 59228 41206
rect 59174 41168 59176 41177
rect 59228 41168 59230 41177
rect 59280 41138 59308 42094
rect 59556 41138 59584 43386
rect 60016 43178 60044 43658
rect 60200 43382 60228 43794
rect 60476 43738 60504 43930
rect 60752 43926 60780 44338
rect 60740 43920 60792 43926
rect 60740 43862 60792 43868
rect 60556 43852 60608 43858
rect 60556 43794 60608 43800
rect 60292 43710 60504 43738
rect 60292 43654 60320 43710
rect 60280 43648 60332 43654
rect 60280 43590 60332 43596
rect 60464 43648 60516 43654
rect 60464 43590 60516 43596
rect 60188 43376 60240 43382
rect 60188 43318 60240 43324
rect 60476 43314 60504 43590
rect 60464 43308 60516 43314
rect 60464 43250 60516 43256
rect 60096 43240 60148 43246
rect 60096 43182 60148 43188
rect 60004 43172 60056 43178
rect 60004 43114 60056 43120
rect 59636 43104 59688 43110
rect 59636 43046 59688 43052
rect 59648 42090 59676 43046
rect 60108 42634 60136 43182
rect 60568 43178 60596 43794
rect 60188 43172 60240 43178
rect 60188 43114 60240 43120
rect 60556 43172 60608 43178
rect 60556 43114 60608 43120
rect 60200 42770 60228 43114
rect 60648 43104 60700 43110
rect 60648 43046 60700 43052
rect 60188 42764 60240 42770
rect 60188 42706 60240 42712
rect 60096 42628 60148 42634
rect 60096 42570 60148 42576
rect 59636 42084 59688 42090
rect 59636 42026 59688 42032
rect 59728 42016 59780 42022
rect 59728 41958 59780 41964
rect 59174 41103 59230 41112
rect 59268 41132 59320 41138
rect 59268 41074 59320 41080
rect 59544 41132 59596 41138
rect 59544 41074 59596 41080
rect 58900 41064 58952 41070
rect 58900 41006 58952 41012
rect 58716 40928 58768 40934
rect 58716 40870 58768 40876
rect 58440 40724 58492 40730
rect 58440 40666 58492 40672
rect 58452 40594 58480 40666
rect 58072 40588 58124 40594
rect 58072 40530 58124 40536
rect 58440 40588 58492 40594
rect 58440 40530 58492 40536
rect 57796 40180 57848 40186
rect 57796 40122 57848 40128
rect 57808 39982 57836 40122
rect 58084 39982 58112 40530
rect 57796 39976 57848 39982
rect 57796 39918 57848 39924
rect 58072 39976 58124 39982
rect 58072 39918 58124 39924
rect 57808 39846 57836 39918
rect 57796 39840 57848 39846
rect 57796 39782 57848 39788
rect 57888 39296 57940 39302
rect 57888 39238 57940 39244
rect 57900 38418 57928 39238
rect 58084 39030 58112 39918
rect 58452 39642 58480 40530
rect 58728 40390 58756 40870
rect 58912 40730 58940 41006
rect 58900 40724 58952 40730
rect 58900 40666 58952 40672
rect 58808 40656 58860 40662
rect 58808 40598 58860 40604
rect 58716 40384 58768 40390
rect 58716 40326 58768 40332
rect 58820 40186 58848 40598
rect 59740 40594 59768 41958
rect 59176 40588 59228 40594
rect 59176 40530 59228 40536
rect 59728 40588 59780 40594
rect 59728 40530 59780 40536
rect 58808 40180 58860 40186
rect 58808 40122 58860 40128
rect 58820 39982 58848 40122
rect 59188 39982 59216 40530
rect 59544 40112 59596 40118
rect 59544 40054 59596 40060
rect 58808 39976 58860 39982
rect 58808 39918 58860 39924
rect 59176 39976 59228 39982
rect 59176 39918 59228 39924
rect 58440 39636 58492 39642
rect 58440 39578 58492 39584
rect 59188 39030 59216 39918
rect 59556 39914 59584 40054
rect 60556 39976 60608 39982
rect 60556 39918 60608 39924
rect 59544 39908 59596 39914
rect 59544 39850 59596 39856
rect 59452 39840 59504 39846
rect 59452 39782 59504 39788
rect 60004 39840 60056 39846
rect 60004 39782 60056 39788
rect 59464 39030 59492 39782
rect 58072 39024 58124 39030
rect 58072 38966 58124 38972
rect 59176 39024 59228 39030
rect 59176 38966 59228 38972
rect 59452 39024 59504 39030
rect 59452 38966 59504 38972
rect 59084 38888 59136 38894
rect 59452 38888 59504 38894
rect 59136 38848 59452 38876
rect 59084 38830 59136 38836
rect 59452 38830 59504 38836
rect 59728 38820 59780 38826
rect 59728 38762 59780 38768
rect 57888 38412 57940 38418
rect 57888 38354 57940 38360
rect 59740 38350 59768 38762
rect 60016 38758 60044 39782
rect 60372 39636 60424 39642
rect 60372 39578 60424 39584
rect 60096 39364 60148 39370
rect 60096 39306 60148 39312
rect 60108 38758 60136 39306
rect 60384 39302 60412 39578
rect 60568 39438 60596 39918
rect 60556 39432 60608 39438
rect 60556 39374 60608 39380
rect 60280 39296 60332 39302
rect 60280 39238 60332 39244
rect 60372 39296 60424 39302
rect 60372 39238 60424 39244
rect 60004 38752 60056 38758
rect 60004 38694 60056 38700
rect 60096 38752 60148 38758
rect 60096 38694 60148 38700
rect 60292 38418 60320 39238
rect 60280 38412 60332 38418
rect 60280 38354 60332 38360
rect 58716 38344 58768 38350
rect 58716 38286 58768 38292
rect 59728 38344 59780 38350
rect 59728 38286 59780 38292
rect 58728 38010 58756 38286
rect 60660 38196 60688 43046
rect 60752 42566 60780 43862
rect 61580 43246 61608 44950
rect 61752 44940 61804 44946
rect 61752 44882 61804 44888
rect 61568 43240 61620 43246
rect 61568 43182 61620 43188
rect 60740 42560 60792 42566
rect 60740 42502 60792 42508
rect 60752 41818 60780 42502
rect 61108 42288 61160 42294
rect 61108 42230 61160 42236
rect 60740 41812 60792 41818
rect 60740 41754 60792 41760
rect 60832 41676 60884 41682
rect 60832 41618 60884 41624
rect 60844 41206 60872 41618
rect 61120 41206 61148 42230
rect 60832 41200 60884 41206
rect 60832 41142 60884 41148
rect 61108 41200 61160 41206
rect 61108 41142 61160 41148
rect 61580 40662 61608 43182
rect 61568 40656 61620 40662
rect 61568 40598 61620 40604
rect 61016 40384 61068 40390
rect 61016 40326 61068 40332
rect 60832 39908 60884 39914
rect 60832 39850 60884 39856
rect 60844 39642 60872 39850
rect 60832 39636 60884 39642
rect 60832 39578 60884 39584
rect 60740 39568 60792 39574
rect 60740 39510 60792 39516
rect 60752 39001 60780 39510
rect 60832 39500 60884 39506
rect 60832 39442 60884 39448
rect 60844 39137 60872 39442
rect 60830 39128 60886 39137
rect 60830 39063 60886 39072
rect 60738 38992 60794 39001
rect 60738 38927 60794 38936
rect 60740 38344 60792 38350
rect 60740 38286 60792 38292
rect 60752 38196 60780 38286
rect 60660 38168 60780 38196
rect 60832 38208 60884 38214
rect 60832 38150 60884 38156
rect 60844 38010 60872 38150
rect 58716 38004 58768 38010
rect 58716 37946 58768 37952
rect 58900 38004 58952 38010
rect 58900 37946 58952 37952
rect 60832 38004 60884 38010
rect 60832 37946 60884 37952
rect 58624 37936 58676 37942
rect 58912 37890 58940 37946
rect 58676 37884 58940 37890
rect 58624 37878 58940 37884
rect 58636 37862 58940 37878
rect 61028 37806 61056 40326
rect 61580 39506 61608 40598
rect 61764 40390 61792 44882
rect 62040 44878 62068 45834
rect 62316 45082 62344 45902
rect 62304 45076 62356 45082
rect 62304 45018 62356 45024
rect 62028 44872 62080 44878
rect 62028 44814 62080 44820
rect 62960 44810 62988 46854
rect 65660 46812 65956 46832
rect 65716 46810 65740 46812
rect 65796 46810 65820 46812
rect 65876 46810 65900 46812
rect 65738 46758 65740 46810
rect 65802 46758 65814 46810
rect 65876 46758 65878 46810
rect 65716 46756 65740 46758
rect 65796 46756 65820 46758
rect 65876 46756 65900 46758
rect 65660 46736 65956 46756
rect 63224 46028 63276 46034
rect 63224 45970 63276 45976
rect 63236 44878 63264 45970
rect 65660 45724 65956 45744
rect 65716 45722 65740 45724
rect 65796 45722 65820 45724
rect 65876 45722 65900 45724
rect 65738 45670 65740 45722
rect 65802 45670 65814 45722
rect 65876 45670 65878 45722
rect 65716 45668 65740 45670
rect 65796 45668 65820 45670
rect 65876 45668 65900 45670
rect 65660 45648 65956 45668
rect 65064 45552 65116 45558
rect 65064 45494 65116 45500
rect 63224 44872 63276 44878
rect 63224 44814 63276 44820
rect 64328 44872 64380 44878
rect 64328 44814 64380 44820
rect 62948 44804 63000 44810
rect 62948 44746 63000 44752
rect 63236 43722 63264 44814
rect 63224 43716 63276 43722
rect 63224 43658 63276 43664
rect 64340 42362 64368 44814
rect 65076 44334 65104 45494
rect 65248 45348 65300 45354
rect 65248 45290 65300 45296
rect 65260 44538 65288 45290
rect 65524 45008 65576 45014
rect 65524 44950 65576 44956
rect 65248 44532 65300 44538
rect 65248 44474 65300 44480
rect 65536 44334 65564 44950
rect 66904 44872 66956 44878
rect 66904 44814 66956 44820
rect 65660 44636 65956 44656
rect 65716 44634 65740 44636
rect 65796 44634 65820 44636
rect 65876 44634 65900 44636
rect 65738 44582 65740 44634
rect 65802 44582 65814 44634
rect 65876 44582 65878 44634
rect 65716 44580 65740 44582
rect 65796 44580 65820 44582
rect 65876 44580 65900 44582
rect 65660 44560 65956 44580
rect 65984 44532 66036 44538
rect 65984 44474 66036 44480
rect 65996 44402 66024 44474
rect 66076 44464 66128 44470
rect 66168 44464 66220 44470
rect 66128 44412 66168 44418
rect 66076 44406 66220 44412
rect 65984 44396 66036 44402
rect 66088 44390 66208 44406
rect 65984 44338 66036 44344
rect 65064 44328 65116 44334
rect 65064 44270 65116 44276
rect 65524 44328 65576 44334
rect 65524 44270 65576 44276
rect 65996 43926 66024 44338
rect 66168 44192 66220 44198
rect 66220 44140 66300 44146
rect 66168 44134 66300 44140
rect 66180 44118 66300 44134
rect 65984 43920 66036 43926
rect 65984 43862 66036 43868
rect 66272 43858 66300 44118
rect 66916 43926 66944 44814
rect 68560 44736 68612 44742
rect 68560 44678 68612 44684
rect 68572 44334 68600 44678
rect 71320 44532 71372 44538
rect 71320 44474 71372 44480
rect 66996 44328 67048 44334
rect 66996 44270 67048 44276
rect 68560 44328 68612 44334
rect 68560 44270 68612 44276
rect 66904 43920 66956 43926
rect 66904 43862 66956 43868
rect 67008 43858 67036 44270
rect 71332 44198 71360 44474
rect 71412 44464 71464 44470
rect 71412 44406 71464 44412
rect 68744 44192 68796 44198
rect 68744 44134 68796 44140
rect 71320 44192 71372 44198
rect 71320 44134 71372 44140
rect 66260 43852 66312 43858
rect 66260 43794 66312 43800
rect 66996 43852 67048 43858
rect 66996 43794 67048 43800
rect 65660 43548 65956 43568
rect 65716 43546 65740 43548
rect 65796 43546 65820 43548
rect 65876 43546 65900 43548
rect 65738 43494 65740 43546
rect 65802 43494 65814 43546
rect 65876 43494 65878 43546
rect 65716 43492 65740 43494
rect 65796 43492 65820 43494
rect 65876 43492 65900 43494
rect 65660 43472 65956 43492
rect 66904 43240 66956 43246
rect 66904 43182 66956 43188
rect 66720 43172 66772 43178
rect 66720 43114 66772 43120
rect 66352 43104 66404 43110
rect 66352 43046 66404 43052
rect 66364 42838 66392 43046
rect 66352 42832 66404 42838
rect 66352 42774 66404 42780
rect 66628 42560 66680 42566
rect 66628 42502 66680 42508
rect 65660 42460 65956 42480
rect 65716 42458 65740 42460
rect 65796 42458 65820 42460
rect 65876 42458 65900 42460
rect 65738 42406 65740 42458
rect 65802 42406 65814 42458
rect 65876 42406 65878 42458
rect 65716 42404 65740 42406
rect 65796 42404 65820 42406
rect 65876 42404 65900 42406
rect 65660 42384 65956 42404
rect 64328 42356 64380 42362
rect 64328 42298 64380 42304
rect 64340 41206 64368 42298
rect 66640 42226 66668 42502
rect 66732 42226 66760 43114
rect 66812 42560 66864 42566
rect 66812 42502 66864 42508
rect 66628 42220 66680 42226
rect 66628 42162 66680 42168
rect 66720 42220 66772 42226
rect 66720 42162 66772 42168
rect 66076 42084 66128 42090
rect 66076 42026 66128 42032
rect 65984 42016 66036 42022
rect 65984 41958 66036 41964
rect 65660 41372 65956 41392
rect 65716 41370 65740 41372
rect 65796 41370 65820 41372
rect 65876 41370 65900 41372
rect 65738 41318 65740 41370
rect 65802 41318 65814 41370
rect 65876 41318 65878 41370
rect 65716 41316 65740 41318
rect 65796 41316 65820 41318
rect 65876 41316 65900 41318
rect 65660 41296 65956 41316
rect 64328 41200 64380 41206
rect 64328 41142 64380 41148
rect 65996 41070 66024 41958
rect 65340 41064 65392 41070
rect 65340 41006 65392 41012
rect 65984 41064 66036 41070
rect 65984 41006 66036 41012
rect 65352 40526 65380 41006
rect 65432 40724 65484 40730
rect 65432 40666 65484 40672
rect 65340 40520 65392 40526
rect 65340 40462 65392 40468
rect 63132 40452 63184 40458
rect 63132 40394 63184 40400
rect 61752 40384 61804 40390
rect 61752 40326 61804 40332
rect 61200 39500 61252 39506
rect 61200 39442 61252 39448
rect 61568 39500 61620 39506
rect 61568 39442 61620 39448
rect 61936 39500 61988 39506
rect 61936 39442 61988 39448
rect 61212 39302 61240 39442
rect 61200 39296 61252 39302
rect 61200 39238 61252 39244
rect 61476 39024 61528 39030
rect 61476 38966 61528 38972
rect 61488 38876 61516 38966
rect 61948 38894 61976 39442
rect 61660 38888 61712 38894
rect 61488 38848 61660 38876
rect 61660 38830 61712 38836
rect 61936 38888 61988 38894
rect 61936 38830 61988 38836
rect 61384 38752 61436 38758
rect 61384 38694 61436 38700
rect 61016 37800 61068 37806
rect 61016 37742 61068 37748
rect 60188 37664 60240 37670
rect 60188 37606 60240 37612
rect 60924 37664 60976 37670
rect 60924 37606 60976 37612
rect 59728 37392 59780 37398
rect 59728 37334 59780 37340
rect 58440 36712 58492 36718
rect 58440 36654 58492 36660
rect 57704 36236 57756 36242
rect 57704 36178 57756 36184
rect 57716 34542 57744 36178
rect 58072 36032 58124 36038
rect 58072 35974 58124 35980
rect 58084 35698 58112 35974
rect 58072 35692 58124 35698
rect 58072 35634 58124 35640
rect 58452 35290 58480 36654
rect 59452 35488 59504 35494
rect 59452 35430 59504 35436
rect 58440 35284 58492 35290
rect 58440 35226 58492 35232
rect 59464 34610 59492 35430
rect 59740 34610 59768 37334
rect 60200 37330 60228 37606
rect 60188 37324 60240 37330
rect 60188 37266 60240 37272
rect 60936 36922 60964 37606
rect 59912 36916 59964 36922
rect 59912 36858 59964 36864
rect 60924 36916 60976 36922
rect 60924 36858 60976 36864
rect 59924 36582 59952 36858
rect 59912 36576 59964 36582
rect 59912 36518 59964 36524
rect 60936 35494 60964 36858
rect 60924 35488 60976 35494
rect 60924 35430 60976 35436
rect 60936 34678 60964 35430
rect 60924 34672 60976 34678
rect 60924 34614 60976 34620
rect 59452 34604 59504 34610
rect 59452 34546 59504 34552
rect 59728 34604 59780 34610
rect 59912 34604 59964 34610
rect 59728 34546 59780 34552
rect 59832 34564 59912 34592
rect 57704 34536 57756 34542
rect 59832 34490 59860 34564
rect 59912 34546 59964 34552
rect 57704 34478 57756 34484
rect 59556 34474 59860 34490
rect 59544 34468 59860 34474
rect 59596 34462 59860 34468
rect 59544 34410 59596 34416
rect 57520 34060 57572 34066
rect 57520 34002 57572 34008
rect 57704 34060 57756 34066
rect 57704 34002 57756 34008
rect 57532 33658 57560 34002
rect 57716 33862 57744 34002
rect 58440 33924 58492 33930
rect 58440 33866 58492 33872
rect 57704 33856 57756 33862
rect 57704 33798 57756 33804
rect 56876 33652 56928 33658
rect 56876 33594 56928 33600
rect 57520 33652 57572 33658
rect 57520 33594 57572 33600
rect 57532 33454 57560 33594
rect 58452 33590 58480 33866
rect 58532 33856 58584 33862
rect 58532 33798 58584 33804
rect 58624 33856 58676 33862
rect 58624 33798 58676 33804
rect 58440 33584 58492 33590
rect 58440 33526 58492 33532
rect 57520 33448 57572 33454
rect 58256 33448 58308 33454
rect 58176 33408 58256 33436
rect 58176 33402 58204 33408
rect 57520 33390 57572 33396
rect 58084 33386 58204 33402
rect 58256 33390 58308 33396
rect 57060 33380 57112 33386
rect 57060 33322 57112 33328
rect 58072 33380 58204 33386
rect 58124 33374 58204 33380
rect 58072 33322 58124 33328
rect 56692 32904 56744 32910
rect 56692 32846 56744 32852
rect 57072 32434 57100 33322
rect 58544 33318 58572 33798
rect 58636 33658 58664 33798
rect 58624 33652 58676 33658
rect 58624 33594 58676 33600
rect 58532 33312 58584 33318
rect 58532 33254 58584 33260
rect 57060 32428 57112 32434
rect 57060 32370 57112 32376
rect 55864 32292 55916 32298
rect 55864 32234 55916 32240
rect 56232 31952 56284 31958
rect 56232 31894 56284 31900
rect 55404 31680 55456 31686
rect 55404 31622 55456 31628
rect 55416 31414 55444 31622
rect 55404 31408 55456 31414
rect 55404 31350 55456 31356
rect 56244 30802 56272 31894
rect 59268 31272 59320 31278
rect 59268 31214 59320 31220
rect 57336 31204 57388 31210
rect 57336 31146 57388 31152
rect 57348 30938 57376 31146
rect 58440 31136 58492 31142
rect 58440 31078 58492 31084
rect 57336 30932 57388 30938
rect 57336 30874 57388 30880
rect 56232 30796 56284 30802
rect 56232 30738 56284 30744
rect 56600 30728 56652 30734
rect 56600 30670 56652 30676
rect 56612 30054 56640 30670
rect 57796 30660 57848 30666
rect 57796 30602 57848 30608
rect 57808 30190 57836 30602
rect 56784 30184 56836 30190
rect 56784 30126 56836 30132
rect 57796 30184 57848 30190
rect 57796 30126 57848 30132
rect 56600 30048 56652 30054
rect 56600 29990 56652 29996
rect 56796 29714 56824 30126
rect 58452 29714 58480 31078
rect 59176 30932 59228 30938
rect 59176 30874 59228 30880
rect 58716 30796 58768 30802
rect 58716 30738 58768 30744
rect 58728 30258 58756 30738
rect 59188 30682 59216 30874
rect 59096 30654 59216 30682
rect 59096 30598 59124 30654
rect 59084 30592 59136 30598
rect 59084 30534 59136 30540
rect 59176 30592 59228 30598
rect 59176 30534 59228 30540
rect 59188 30258 59216 30534
rect 58716 30252 58768 30258
rect 58716 30194 58768 30200
rect 59176 30252 59228 30258
rect 59176 30194 59228 30200
rect 55496 29708 55548 29714
rect 55496 29650 55548 29656
rect 56784 29708 56836 29714
rect 56784 29650 56836 29656
rect 57888 29708 57940 29714
rect 57888 29650 57940 29656
rect 58440 29708 58492 29714
rect 58440 29650 58492 29656
rect 55312 29572 55364 29578
rect 55312 29514 55364 29520
rect 55508 29306 55536 29650
rect 56796 29306 56824 29650
rect 55496 29300 55548 29306
rect 55496 29242 55548 29248
rect 56784 29300 56836 29306
rect 56784 29242 56836 29248
rect 57796 29028 57848 29034
rect 57796 28970 57848 28976
rect 56692 26308 56744 26314
rect 56692 26250 56744 26256
rect 55128 26240 55180 26246
rect 56600 26240 56652 26246
rect 55128 26182 55180 26188
rect 56598 26208 56600 26217
rect 56652 26208 56654 26217
rect 56598 26143 56654 26152
rect 56704 25673 56732 26250
rect 56690 25664 56746 25673
rect 56690 25599 56746 25608
rect 57808 21865 57836 28970
rect 57900 26518 57928 29650
rect 58728 29510 58756 30194
rect 59084 29572 59136 29578
rect 59084 29514 59136 29520
rect 58716 29504 58768 29510
rect 58716 29446 58768 29452
rect 58992 29504 59044 29510
rect 58992 29446 59044 29452
rect 57888 26512 57940 26518
rect 57888 26454 57940 26460
rect 59004 22893 59032 29446
rect 59096 25069 59124 29514
rect 59176 29504 59228 29510
rect 59176 29446 59228 29452
rect 59188 29073 59216 29446
rect 59280 29170 59308 31214
rect 59452 30184 59504 30190
rect 59452 30126 59504 30132
rect 59360 30048 59412 30054
rect 59360 29990 59412 29996
rect 59268 29164 59320 29170
rect 59268 29106 59320 29112
rect 59174 29064 59230 29073
rect 59174 28999 59230 29008
rect 59082 25060 59138 25069
rect 59082 24995 59138 25004
rect 58990 22884 59046 22893
rect 58990 22819 59046 22828
rect 57794 21856 57850 21865
rect 57794 21791 57850 21800
rect 59280 20717 59308 29106
rect 59372 25613 59400 29990
rect 59358 25604 59414 25613
rect 59358 25539 59414 25548
rect 59358 23916 59414 23925
rect 59464 23902 59492 30126
rect 59556 29578 59584 34410
rect 60936 33998 60964 34614
rect 60924 33992 60976 33998
rect 60924 33934 60976 33940
rect 61292 33992 61344 33998
rect 61292 33934 61344 33940
rect 61108 33448 61160 33454
rect 61108 33390 61160 33396
rect 60280 32224 60332 32230
rect 60280 32166 60332 32172
rect 60292 31210 60320 32166
rect 60464 31272 60516 31278
rect 60464 31214 60516 31220
rect 60832 31272 60884 31278
rect 60832 31214 60884 31220
rect 60280 31204 60332 31210
rect 60280 31146 60332 31152
rect 60476 31142 60504 31214
rect 60844 31142 60872 31214
rect 60464 31136 60516 31142
rect 60464 31078 60516 31084
rect 60832 31136 60884 31142
rect 60832 31078 60884 31084
rect 60372 30592 60424 30598
rect 60372 30534 60424 30540
rect 60384 30190 60412 30534
rect 60476 30394 60504 31078
rect 60924 30728 60976 30734
rect 60924 30670 60976 30676
rect 60936 30394 60964 30670
rect 60464 30388 60516 30394
rect 60464 30330 60516 30336
rect 60924 30388 60976 30394
rect 60924 30330 60976 30336
rect 60372 30184 60424 30190
rect 60476 30172 60504 30330
rect 61120 30326 61148 33390
rect 61108 30320 61160 30326
rect 61108 30262 61160 30268
rect 60476 30144 60688 30172
rect 60372 30126 60424 30132
rect 60660 30138 60688 30144
rect 60660 30122 60872 30138
rect 60188 30116 60240 30122
rect 60660 30116 60884 30122
rect 60660 30110 60832 30116
rect 60188 30058 60240 30064
rect 60832 30058 60884 30064
rect 60004 30048 60056 30054
rect 60004 29990 60056 29996
rect 59636 29640 59688 29646
rect 59636 29582 59688 29588
rect 59544 29572 59596 29578
rect 59544 29514 59596 29520
rect 59414 23874 59492 23902
rect 59358 23851 59414 23860
rect 59358 21448 59414 21457
rect 59358 21383 59414 21392
rect 59372 20806 59400 21383
rect 59360 20800 59412 20806
rect 59360 20742 59412 20748
rect 59266 20708 59322 20717
rect 59266 20643 59322 20652
rect 59372 19629 59400 20742
rect 59358 19620 59414 19629
rect 59358 19555 59414 19564
rect 59360 17403 59412 17406
rect 59358 17400 59414 17403
rect 59358 17394 59360 17400
rect 59412 17394 59414 17400
rect 59358 17329 59414 17338
rect 59556 4729 59584 29514
rect 59648 17406 59676 29582
rect 59728 29504 59780 29510
rect 59728 29446 59780 29452
rect 59912 29504 59964 29510
rect 59912 29446 59964 29452
rect 59740 29034 59768 29446
rect 59728 29028 59780 29034
rect 59728 28970 59780 28976
rect 59924 20806 59952 29446
rect 60016 29238 60044 29990
rect 60200 29646 60228 30058
rect 60648 30048 60700 30054
rect 60646 30016 60648 30025
rect 60700 30016 60702 30025
rect 60646 29951 60702 29960
rect 60556 29844 60608 29850
rect 60556 29786 60608 29792
rect 60568 29714 60596 29786
rect 61304 29782 61332 33934
rect 61396 33454 61424 38694
rect 62212 38412 62264 38418
rect 62212 38354 62264 38360
rect 62224 38214 62252 38354
rect 62212 38208 62264 38214
rect 62212 38150 62264 38156
rect 63144 37670 63172 40394
rect 65156 39908 65208 39914
rect 65156 39850 65208 39856
rect 63590 39128 63646 39137
rect 63590 39063 63646 39072
rect 63316 37800 63368 37806
rect 63316 37742 63368 37748
rect 63328 37670 63356 37742
rect 63132 37664 63184 37670
rect 63132 37606 63184 37612
rect 63316 37664 63368 37670
rect 63316 37606 63368 37612
rect 63328 37466 63356 37606
rect 63316 37460 63368 37466
rect 63316 37402 63368 37408
rect 63132 37392 63184 37398
rect 63132 37334 63184 37340
rect 62028 36780 62080 36786
rect 62028 36722 62080 36728
rect 62040 36242 62068 36722
rect 63144 36650 63172 37334
rect 63224 37120 63276 37126
rect 63224 37062 63276 37068
rect 63132 36644 63184 36650
rect 63132 36586 63184 36592
rect 62028 36236 62080 36242
rect 62028 36178 62080 36184
rect 62040 35698 62068 36178
rect 62764 36032 62816 36038
rect 62764 35974 62816 35980
rect 62776 35834 62804 35974
rect 62764 35828 62816 35834
rect 62764 35770 62816 35776
rect 62028 35692 62080 35698
rect 62028 35634 62080 35640
rect 63144 35630 63172 36586
rect 63132 35624 63184 35630
rect 63132 35566 63184 35572
rect 63236 35494 63264 37062
rect 63224 35488 63276 35494
rect 63224 35430 63276 35436
rect 63236 35154 63264 35430
rect 63224 35148 63276 35154
rect 63224 35090 63276 35096
rect 63040 34740 63092 34746
rect 63040 34682 63092 34688
rect 62580 34672 62632 34678
rect 62580 34614 62632 34620
rect 62396 34536 62448 34542
rect 62396 34478 62448 34484
rect 62408 34406 62436 34478
rect 62396 34400 62448 34406
rect 62396 34342 62448 34348
rect 61660 33584 61712 33590
rect 61660 33526 61712 33532
rect 61384 33448 61436 33454
rect 61384 33390 61436 33396
rect 61566 33008 61622 33017
rect 61566 32943 61568 32952
rect 61620 32943 61622 32952
rect 61568 32914 61620 32920
rect 61672 32502 61700 33526
rect 62028 33108 62080 33114
rect 62028 33050 62080 33056
rect 62040 32978 62068 33050
rect 62408 32978 62436 34342
rect 62592 33522 62620 34614
rect 63052 34542 63080 34682
rect 63040 34536 63092 34542
rect 63040 34478 63092 34484
rect 62580 33516 62632 33522
rect 62580 33458 62632 33464
rect 63052 32978 63080 34478
rect 63132 34128 63184 34134
rect 63132 34070 63184 34076
rect 63144 33386 63172 34070
rect 63132 33380 63184 33386
rect 63132 33322 63184 33328
rect 61844 32972 61896 32978
rect 61844 32914 61896 32920
rect 62028 32972 62080 32978
rect 62028 32914 62080 32920
rect 62396 32972 62448 32978
rect 62396 32914 62448 32920
rect 63040 32972 63092 32978
rect 63040 32914 63092 32920
rect 61660 32496 61712 32502
rect 61660 32438 61712 32444
rect 61856 32366 61884 32914
rect 61844 32360 61896 32366
rect 61844 32302 61896 32308
rect 62040 32298 62068 32914
rect 63224 32768 63276 32774
rect 63224 32710 63276 32716
rect 63500 32768 63552 32774
rect 63500 32710 63552 32716
rect 62304 32564 62356 32570
rect 62304 32506 62356 32512
rect 62028 32292 62080 32298
rect 62028 32234 62080 32240
rect 62120 32224 62172 32230
rect 62120 32166 62172 32172
rect 62132 31482 62160 32166
rect 62316 32026 62344 32506
rect 62396 32224 62448 32230
rect 62396 32166 62448 32172
rect 62408 32026 62436 32166
rect 62304 32020 62356 32026
rect 62304 31962 62356 31968
rect 62396 32020 62448 32026
rect 62396 31962 62448 31968
rect 63236 31482 63264 32710
rect 63512 32366 63540 32710
rect 63500 32360 63552 32366
rect 63500 32302 63552 32308
rect 61936 31476 61988 31482
rect 61936 31418 61988 31424
rect 62120 31476 62172 31482
rect 62120 31418 62172 31424
rect 63224 31476 63276 31482
rect 63224 31418 63276 31424
rect 61948 31210 61976 31418
rect 62132 31278 62160 31418
rect 62120 31272 62172 31278
rect 62120 31214 62172 31220
rect 61936 31204 61988 31210
rect 61936 31146 61988 31152
rect 62212 31204 62264 31210
rect 62212 31146 62264 31152
rect 62396 31204 62448 31210
rect 62396 31146 62448 31152
rect 62028 31136 62080 31142
rect 62028 31078 62080 31084
rect 61660 30796 61712 30802
rect 61660 30738 61712 30744
rect 61936 30796 61988 30802
rect 61936 30738 61988 30744
rect 61672 30598 61700 30738
rect 61948 30598 61976 30738
rect 61660 30592 61712 30598
rect 61660 30534 61712 30540
rect 61936 30592 61988 30598
rect 61936 30534 61988 30540
rect 61948 30326 61976 30534
rect 61936 30320 61988 30326
rect 61936 30262 61988 30268
rect 61948 30025 61976 30262
rect 62040 30190 62068 31078
rect 62224 30938 62252 31146
rect 62212 30932 62264 30938
rect 62212 30874 62264 30880
rect 62408 30870 62436 31146
rect 62396 30864 62448 30870
rect 62396 30806 62448 30812
rect 62028 30184 62080 30190
rect 62028 30126 62080 30132
rect 61934 30016 61990 30025
rect 61934 29951 61990 29960
rect 61292 29776 61344 29782
rect 61292 29718 61344 29724
rect 60556 29708 60608 29714
rect 60556 29650 60608 29656
rect 60188 29640 60240 29646
rect 60188 29582 60240 29588
rect 61304 29510 61332 29718
rect 61292 29504 61344 29510
rect 61292 29446 61344 29452
rect 61568 29504 61620 29510
rect 61568 29446 61620 29452
rect 60004 29232 60056 29238
rect 60004 29174 60056 29180
rect 61580 29170 61608 29446
rect 63512 29238 63540 32302
rect 63604 31482 63632 39063
rect 65168 38894 65196 39850
rect 64972 38888 65024 38894
rect 64972 38830 65024 38836
rect 65156 38888 65208 38894
rect 65156 38830 65208 38836
rect 64236 38820 64288 38826
rect 64236 38762 64288 38768
rect 64248 38418 64276 38762
rect 64984 38758 65012 38830
rect 64972 38752 65024 38758
rect 64972 38694 65024 38700
rect 64984 38486 65012 38694
rect 64972 38480 65024 38486
rect 64972 38422 65024 38428
rect 64236 38412 64288 38418
rect 64236 38354 64288 38360
rect 64696 37868 64748 37874
rect 64696 37810 64748 37816
rect 64708 37670 64736 37810
rect 65168 37806 65196 38830
rect 65444 38214 65472 40666
rect 65660 40284 65956 40304
rect 65716 40282 65740 40284
rect 65796 40282 65820 40284
rect 65876 40282 65900 40284
rect 65738 40230 65740 40282
rect 65802 40230 65814 40282
rect 65876 40230 65878 40282
rect 65716 40228 65740 40230
rect 65796 40228 65820 40230
rect 65876 40228 65900 40230
rect 65660 40208 65956 40228
rect 66088 39914 66116 42026
rect 66444 42016 66496 42022
rect 66444 41958 66496 41964
rect 66456 41206 66484 41958
rect 66628 41472 66680 41478
rect 66628 41414 66680 41420
rect 66444 41200 66496 41206
rect 66444 41142 66496 41148
rect 66640 41070 66668 41414
rect 66628 41064 66680 41070
rect 66628 41006 66680 41012
rect 66732 41002 66760 42162
rect 66824 41834 66852 42502
rect 66916 42022 66944 43182
rect 67008 43110 67036 43794
rect 67086 43344 67142 43353
rect 67086 43279 67142 43288
rect 67100 43246 67128 43279
rect 67088 43240 67140 43246
rect 67088 43182 67140 43188
rect 66996 43104 67048 43110
rect 66996 43046 67048 43052
rect 68756 42770 68784 44134
rect 71044 43376 71096 43382
rect 71044 43318 71096 43324
rect 71056 43246 71084 43318
rect 71044 43240 71096 43246
rect 71044 43182 71096 43188
rect 71228 43240 71280 43246
rect 71228 43182 71280 43188
rect 71240 42770 71268 43182
rect 66996 42764 67048 42770
rect 66996 42706 67048 42712
rect 68744 42764 68796 42770
rect 68744 42706 68796 42712
rect 71228 42764 71280 42770
rect 71228 42706 71280 42712
rect 67008 42362 67036 42706
rect 71424 42702 71452 44406
rect 72884 44328 72936 44334
rect 72884 44270 72936 44276
rect 72896 43994 72924 44270
rect 72976 44192 73028 44198
rect 72976 44134 73028 44140
rect 72884 43988 72936 43994
rect 72884 43930 72936 43936
rect 72516 43920 72568 43926
rect 72516 43862 72568 43868
rect 71596 43852 71648 43858
rect 71596 43794 71648 43800
rect 71608 42838 71636 43794
rect 71780 43784 71832 43790
rect 71780 43726 71832 43732
rect 71596 42832 71648 42838
rect 71596 42774 71648 42780
rect 71412 42696 71464 42702
rect 71412 42638 71464 42644
rect 67456 42628 67508 42634
rect 67456 42570 67508 42576
rect 66996 42356 67048 42362
rect 66996 42298 67048 42304
rect 67468 42158 67496 42570
rect 69204 42560 69256 42566
rect 69204 42502 69256 42508
rect 69216 42158 69244 42502
rect 70492 42356 70544 42362
rect 70492 42298 70544 42304
rect 67456 42152 67508 42158
rect 67456 42094 67508 42100
rect 69204 42152 69256 42158
rect 69204 42094 69256 42100
rect 67468 42022 67496 42094
rect 66904 42016 66956 42022
rect 66904 41958 66956 41964
rect 67456 42016 67508 42022
rect 67456 41958 67508 41964
rect 66824 41806 66944 41834
rect 66812 41676 66864 41682
rect 66812 41618 66864 41624
rect 66720 40996 66772 41002
rect 66720 40938 66772 40944
rect 66824 40526 66852 41618
rect 66916 41138 66944 41806
rect 70504 41750 70532 42298
rect 71792 42022 71820 43726
rect 71872 43240 71924 43246
rect 71872 43182 71924 43188
rect 71884 42090 71912 43182
rect 71964 43172 72016 43178
rect 71964 43114 72016 43120
rect 71976 42158 72004 43114
rect 72424 43104 72476 43110
rect 72424 43046 72476 43052
rect 72436 42770 72464 43046
rect 72528 42770 72556 43862
rect 72792 43852 72844 43858
rect 72792 43794 72844 43800
rect 72056 42764 72108 42770
rect 72056 42706 72108 42712
rect 72424 42764 72476 42770
rect 72424 42706 72476 42712
rect 72516 42764 72568 42770
rect 72516 42706 72568 42712
rect 72068 42362 72096 42706
rect 72056 42356 72108 42362
rect 72056 42298 72108 42304
rect 72528 42226 72556 42706
rect 72804 42634 72832 43794
rect 72988 43382 73016 44134
rect 72976 43376 73028 43382
rect 72976 43318 73028 43324
rect 72792 42628 72844 42634
rect 72792 42570 72844 42576
rect 72516 42220 72568 42226
rect 72516 42162 72568 42168
rect 71964 42152 72016 42158
rect 71964 42094 72016 42100
rect 71872 42084 71924 42090
rect 71872 42026 71924 42032
rect 71780 42016 71832 42022
rect 71780 41958 71832 41964
rect 70492 41744 70544 41750
rect 70492 41686 70544 41692
rect 71872 41676 71924 41682
rect 71872 41618 71924 41624
rect 67362 41168 67418 41177
rect 66904 41132 66956 41138
rect 67362 41103 67418 41112
rect 71594 41168 71650 41177
rect 71884 41138 71912 41618
rect 71594 41103 71650 41112
rect 71872 41132 71924 41138
rect 66904 41074 66956 41080
rect 66916 40934 66944 41074
rect 67376 41070 67404 41103
rect 71608 41070 71636 41103
rect 71872 41074 71924 41080
rect 67364 41064 67416 41070
rect 67364 41006 67416 41012
rect 71596 41064 71648 41070
rect 71596 41006 71648 41012
rect 71778 41032 71834 41041
rect 67088 40996 67140 41002
rect 67088 40938 67140 40944
rect 71688 40996 71740 41002
rect 71778 40967 71834 40976
rect 71688 40938 71740 40944
rect 66904 40928 66956 40934
rect 66904 40870 66956 40876
rect 67100 40594 67128 40938
rect 67640 40928 67692 40934
rect 67640 40870 67692 40876
rect 67088 40588 67140 40594
rect 67088 40530 67140 40536
rect 66812 40520 66864 40526
rect 66812 40462 66864 40468
rect 67456 40520 67508 40526
rect 67456 40462 67508 40468
rect 66076 39908 66128 39914
rect 66076 39850 66128 39856
rect 66088 39574 66116 39850
rect 66076 39568 66128 39574
rect 66076 39510 66128 39516
rect 66824 39506 66852 40462
rect 67364 39840 67416 39846
rect 67364 39782 67416 39788
rect 67376 39642 67404 39782
rect 67364 39636 67416 39642
rect 67364 39578 67416 39584
rect 67468 39506 67496 40462
rect 67652 39914 67680 40870
rect 71700 40730 71728 40938
rect 71792 40934 71820 40967
rect 71780 40928 71832 40934
rect 71780 40870 71832 40876
rect 71688 40724 71740 40730
rect 71688 40666 71740 40672
rect 71136 39976 71188 39982
rect 71136 39918 71188 39924
rect 67640 39908 67692 39914
rect 67640 39850 67692 39856
rect 69756 39636 69808 39642
rect 69756 39578 69808 39584
rect 65524 39500 65576 39506
rect 65524 39442 65576 39448
rect 66812 39500 66864 39506
rect 66812 39442 66864 39448
rect 67456 39500 67508 39506
rect 67456 39442 67508 39448
rect 65536 38894 65564 39442
rect 68836 39432 68888 39438
rect 68836 39374 68888 39380
rect 66076 39364 66128 39370
rect 66076 39306 66128 39312
rect 65660 39196 65956 39216
rect 65716 39194 65740 39196
rect 65796 39194 65820 39196
rect 65876 39194 65900 39196
rect 65738 39142 65740 39194
rect 65802 39142 65814 39194
rect 65876 39142 65878 39194
rect 65716 39140 65740 39142
rect 65796 39140 65820 39142
rect 65876 39140 65900 39142
rect 65660 39120 65956 39140
rect 66088 38962 66116 39306
rect 66904 39296 66956 39302
rect 66904 39238 66956 39244
rect 66916 39001 66944 39238
rect 68848 39030 68876 39374
rect 69768 39030 69796 39578
rect 71148 39370 71176 39918
rect 71688 39840 71740 39846
rect 71688 39782 71740 39788
rect 71700 39642 71728 39782
rect 71688 39636 71740 39642
rect 71688 39578 71740 39584
rect 71596 39568 71648 39574
rect 71596 39510 71648 39516
rect 71412 39500 71464 39506
rect 71412 39442 71464 39448
rect 71136 39364 71188 39370
rect 71136 39306 71188 39312
rect 71424 39302 71452 39442
rect 71608 39438 71636 39510
rect 71596 39432 71648 39438
rect 71596 39374 71648 39380
rect 71412 39296 71464 39302
rect 71412 39238 71464 39244
rect 68376 39024 68428 39030
rect 66902 38992 66958 39001
rect 65984 38956 66036 38962
rect 65984 38898 66036 38904
rect 66076 38956 66128 38962
rect 68376 38966 68428 38972
rect 68836 39024 68888 39030
rect 68836 38966 68888 38972
rect 69756 39024 69808 39030
rect 69756 38966 69808 38972
rect 66902 38927 66958 38936
rect 66076 38898 66128 38904
rect 65524 38888 65576 38894
rect 65524 38830 65576 38836
rect 65432 38208 65484 38214
rect 65432 38150 65484 38156
rect 64880 37800 64932 37806
rect 65156 37800 65208 37806
rect 64932 37748 65104 37754
rect 64880 37742 65104 37748
rect 65156 37742 65208 37748
rect 64892 37738 65104 37742
rect 64892 37732 65116 37738
rect 64892 37726 65064 37732
rect 65064 37674 65116 37680
rect 64696 37664 64748 37670
rect 64696 37606 64748 37612
rect 64604 37324 64656 37330
rect 64604 37266 64656 37272
rect 65340 37324 65392 37330
rect 65340 37266 65392 37272
rect 64616 36718 64644 37266
rect 65248 37256 65300 37262
rect 65248 37198 65300 37204
rect 64880 37188 64932 37194
rect 64880 37130 64932 37136
rect 64892 36922 64920 37130
rect 65260 37126 65288 37198
rect 65248 37120 65300 37126
rect 65248 37062 65300 37068
rect 65260 36922 65288 37062
rect 64880 36916 64932 36922
rect 64880 36858 64932 36864
rect 65248 36916 65300 36922
rect 65248 36858 65300 36864
rect 65260 36718 65288 36858
rect 65352 36854 65380 37266
rect 65340 36848 65392 36854
rect 65340 36790 65392 36796
rect 64420 36712 64472 36718
rect 64420 36654 64472 36660
rect 64604 36712 64656 36718
rect 64604 36654 64656 36660
rect 65248 36712 65300 36718
rect 65248 36654 65300 36660
rect 64432 36310 64460 36654
rect 65444 36650 65472 38150
rect 65536 37806 65564 38830
rect 65660 38108 65956 38128
rect 65716 38106 65740 38108
rect 65796 38106 65820 38108
rect 65876 38106 65900 38108
rect 65738 38054 65740 38106
rect 65802 38054 65814 38106
rect 65876 38054 65878 38106
rect 65716 38052 65740 38054
rect 65796 38052 65820 38054
rect 65876 38052 65900 38054
rect 65660 38032 65956 38052
rect 65524 37800 65576 37806
rect 65524 37742 65576 37748
rect 65996 37330 66024 38898
rect 66916 38894 66944 38927
rect 66904 38888 66956 38894
rect 66904 38830 66956 38836
rect 68284 38752 68336 38758
rect 68284 38694 68336 38700
rect 66260 38276 66312 38282
rect 66260 38218 66312 38224
rect 66168 37664 66220 37670
rect 66168 37606 66220 37612
rect 66076 37460 66128 37466
rect 66076 37402 66128 37408
rect 65984 37324 66036 37330
rect 65984 37266 66036 37272
rect 65660 37020 65956 37040
rect 65716 37018 65740 37020
rect 65796 37018 65820 37020
rect 65876 37018 65900 37020
rect 65738 36966 65740 37018
rect 65802 36966 65814 37018
rect 65876 36966 65878 37018
rect 65716 36964 65740 36966
rect 65796 36964 65820 36966
rect 65876 36964 65900 36966
rect 65660 36944 65956 36964
rect 66088 36854 66116 37402
rect 66076 36848 66128 36854
rect 66076 36790 66128 36796
rect 66180 36718 66208 37606
rect 66272 37466 66300 38218
rect 66444 37732 66496 37738
rect 66444 37674 66496 37680
rect 66260 37460 66312 37466
rect 66260 37402 66312 37408
rect 66456 36786 66484 37674
rect 66996 37392 67048 37398
rect 66996 37334 67048 37340
rect 66444 36780 66496 36786
rect 66444 36722 66496 36728
rect 65984 36712 66036 36718
rect 65984 36654 66036 36660
rect 66168 36712 66220 36718
rect 66168 36654 66220 36660
rect 65432 36644 65484 36650
rect 65432 36586 65484 36592
rect 64420 36304 64472 36310
rect 64420 36246 64472 36252
rect 65660 35932 65956 35952
rect 65716 35930 65740 35932
rect 65796 35930 65820 35932
rect 65876 35930 65900 35932
rect 65738 35878 65740 35930
rect 65802 35878 65814 35930
rect 65876 35878 65878 35930
rect 65716 35876 65740 35878
rect 65796 35876 65820 35878
rect 65876 35876 65900 35878
rect 65660 35856 65956 35876
rect 65996 35834 66024 36654
rect 67008 36310 67036 37334
rect 68100 36576 68152 36582
rect 68100 36518 68152 36524
rect 66996 36304 67048 36310
rect 66996 36246 67048 36252
rect 67640 36236 67692 36242
rect 67640 36178 67692 36184
rect 68008 36236 68060 36242
rect 68008 36178 68060 36184
rect 65984 35828 66036 35834
rect 65984 35770 66036 35776
rect 66812 35828 66864 35834
rect 66812 35770 66864 35776
rect 66824 35630 66852 35770
rect 67652 35698 67680 36178
rect 67732 36168 67784 36174
rect 67732 36110 67784 36116
rect 67916 36168 67968 36174
rect 67916 36110 67968 36116
rect 67640 35692 67692 35698
rect 67640 35634 67692 35640
rect 66812 35624 66864 35630
rect 66812 35566 66864 35572
rect 65984 35556 66036 35562
rect 65984 35498 66036 35504
rect 65524 35488 65576 35494
rect 65524 35430 65576 35436
rect 64708 35278 64828 35306
rect 64708 35193 64736 35278
rect 64800 35222 64828 35278
rect 64788 35216 64840 35222
rect 64694 35184 64750 35193
rect 64788 35158 64840 35164
rect 64694 35119 64750 35128
rect 65536 34474 65564 35430
rect 65660 34844 65956 34864
rect 65716 34842 65740 34844
rect 65796 34842 65820 34844
rect 65876 34842 65900 34844
rect 65738 34790 65740 34842
rect 65802 34790 65814 34842
rect 65876 34790 65878 34842
rect 65716 34788 65740 34790
rect 65796 34788 65820 34790
rect 65876 34788 65900 34790
rect 65660 34768 65956 34788
rect 65996 34542 66024 35498
rect 67744 34950 67772 36110
rect 67928 35154 67956 36110
rect 68020 35834 68048 36178
rect 68008 35828 68060 35834
rect 68008 35770 68060 35776
rect 67916 35148 67968 35154
rect 67916 35090 67968 35096
rect 67732 34944 67784 34950
rect 67732 34886 67784 34892
rect 68008 34944 68060 34950
rect 68008 34886 68060 34892
rect 65984 34536 66036 34542
rect 65984 34478 66036 34484
rect 65524 34468 65576 34474
rect 65524 34410 65576 34416
rect 65996 34134 66024 34478
rect 65984 34128 66036 34134
rect 65984 34070 66036 34076
rect 67640 33992 67692 33998
rect 67640 33934 67692 33940
rect 65660 33756 65956 33776
rect 65716 33754 65740 33756
rect 65796 33754 65820 33756
rect 65876 33754 65900 33756
rect 65738 33702 65740 33754
rect 65802 33702 65814 33754
rect 65876 33702 65878 33754
rect 65716 33700 65740 33702
rect 65796 33700 65820 33702
rect 65876 33700 65900 33702
rect 65660 33680 65956 33700
rect 66996 33040 67048 33046
rect 66994 33008 66996 33017
rect 67048 33008 67050 33017
rect 66994 32943 67050 32952
rect 67456 32972 67508 32978
rect 67008 32774 67036 32943
rect 67456 32914 67508 32920
rect 66996 32768 67048 32774
rect 66996 32710 67048 32716
rect 65660 32668 65956 32688
rect 65716 32666 65740 32668
rect 65796 32666 65820 32668
rect 65876 32666 65900 32668
rect 65738 32614 65740 32666
rect 65802 32614 65814 32666
rect 65876 32614 65878 32666
rect 65716 32612 65740 32614
rect 65796 32612 65820 32614
rect 65876 32612 65900 32614
rect 65660 32592 65956 32612
rect 67468 32434 67496 32914
rect 67088 32428 67140 32434
rect 67088 32370 67140 32376
rect 67456 32428 67508 32434
rect 67456 32370 67508 32376
rect 66904 31816 66956 31822
rect 66904 31758 66956 31764
rect 65660 31580 65956 31600
rect 65716 31578 65740 31580
rect 65796 31578 65820 31580
rect 65876 31578 65900 31580
rect 65738 31526 65740 31578
rect 65802 31526 65814 31578
rect 65876 31526 65878 31578
rect 65716 31524 65740 31526
rect 65796 31524 65820 31526
rect 65876 31524 65900 31526
rect 65660 31504 65956 31524
rect 63592 31476 63644 31482
rect 63592 31418 63644 31424
rect 66916 31414 66944 31758
rect 66904 31408 66956 31414
rect 66904 31350 66956 31356
rect 66996 30796 67048 30802
rect 66996 30738 67048 30744
rect 67008 30598 67036 30738
rect 66996 30592 67048 30598
rect 66996 30534 67048 30540
rect 65660 30492 65956 30512
rect 65716 30490 65740 30492
rect 65796 30490 65820 30492
rect 65876 30490 65900 30492
rect 65738 30438 65740 30490
rect 65802 30438 65814 30490
rect 65876 30438 65878 30490
rect 65716 30436 65740 30438
rect 65796 30436 65820 30438
rect 65876 30436 65900 30438
rect 65660 30416 65956 30436
rect 66076 30252 66128 30258
rect 66076 30194 66128 30200
rect 66088 30054 66116 30194
rect 67100 30190 67128 32370
rect 67548 32224 67600 32230
rect 67548 32166 67600 32172
rect 67560 31958 67588 32166
rect 67548 31952 67600 31958
rect 67548 31894 67600 31900
rect 67180 31884 67232 31890
rect 67180 31826 67232 31832
rect 67192 31142 67220 31826
rect 67272 31816 67324 31822
rect 67272 31758 67324 31764
rect 67284 31686 67312 31758
rect 67272 31680 67324 31686
rect 67272 31622 67324 31628
rect 67548 31680 67600 31686
rect 67548 31622 67600 31628
rect 67456 31204 67508 31210
rect 67456 31146 67508 31152
rect 67180 31136 67232 31142
rect 67180 31078 67232 31084
rect 67468 30938 67496 31146
rect 67560 30938 67588 31622
rect 67456 30932 67508 30938
rect 67456 30874 67508 30880
rect 67548 30932 67600 30938
rect 67548 30874 67600 30880
rect 67088 30184 67140 30190
rect 67088 30126 67140 30132
rect 66076 30048 66128 30054
rect 66076 29990 66128 29996
rect 65660 29404 65956 29424
rect 65716 29402 65740 29404
rect 65796 29402 65820 29404
rect 65876 29402 65900 29404
rect 65738 29350 65740 29402
rect 65802 29350 65814 29402
rect 65876 29350 65878 29402
rect 65716 29348 65740 29350
rect 65796 29348 65820 29350
rect 65876 29348 65900 29350
rect 65660 29328 65956 29348
rect 66088 29306 66116 29990
rect 67652 29850 67680 33934
rect 68020 33658 68048 34886
rect 68112 34746 68140 36518
rect 68100 34740 68152 34746
rect 68100 34682 68152 34688
rect 68296 34678 68324 38694
rect 68284 34672 68336 34678
rect 68284 34614 68336 34620
rect 68100 34604 68152 34610
rect 68100 34546 68152 34552
rect 68008 33652 68060 33658
rect 68008 33594 68060 33600
rect 67916 33108 67968 33114
rect 67916 33050 67968 33056
rect 67928 32978 67956 33050
rect 68112 32978 68140 34546
rect 67916 32972 67968 32978
rect 67916 32914 67968 32920
rect 68100 32972 68152 32978
rect 68100 32914 68152 32920
rect 68112 32774 68140 32914
rect 68100 32768 68152 32774
rect 68100 32710 68152 32716
rect 68388 31414 68416 38966
rect 71424 38962 71452 39238
rect 69296 38956 69348 38962
rect 69296 38898 69348 38904
rect 71412 38956 71464 38962
rect 71412 38898 71464 38904
rect 68560 37732 68612 37738
rect 68560 37674 68612 37680
rect 68572 36378 68600 37674
rect 68652 36644 68704 36650
rect 68652 36586 68704 36592
rect 68664 36378 68692 36586
rect 68560 36372 68612 36378
rect 68560 36314 68612 36320
rect 68652 36372 68704 36378
rect 68652 36314 68704 36320
rect 68652 36032 68704 36038
rect 68652 35974 68704 35980
rect 68664 35601 68692 35974
rect 68650 35592 68706 35601
rect 68650 35527 68706 35536
rect 68560 35148 68612 35154
rect 68560 35090 68612 35096
rect 68572 33998 68600 35090
rect 68928 34740 68980 34746
rect 68928 34682 68980 34688
rect 68652 34672 68704 34678
rect 68704 34620 68876 34626
rect 68652 34614 68876 34620
rect 68664 34598 68876 34614
rect 68848 34542 68876 34598
rect 68940 34542 68968 34682
rect 68836 34536 68888 34542
rect 68836 34478 68888 34484
rect 68928 34536 68980 34542
rect 68928 34478 68980 34484
rect 68744 34400 68796 34406
rect 68744 34342 68796 34348
rect 68560 33992 68612 33998
rect 68560 33934 68612 33940
rect 68756 33114 68784 34342
rect 69308 33454 69336 38898
rect 71424 38758 71452 38898
rect 71700 38894 71728 39578
rect 71792 39506 71820 40870
rect 71976 39642 72004 42094
rect 72700 42084 72752 42090
rect 72700 42026 72752 42032
rect 72148 41676 72200 41682
rect 72148 41618 72200 41624
rect 72424 41676 72476 41682
rect 72424 41618 72476 41624
rect 72160 39982 72188 41618
rect 72436 41138 72464 41618
rect 72608 41472 72660 41478
rect 72608 41414 72660 41420
rect 72514 41168 72570 41177
rect 72424 41132 72476 41138
rect 72514 41103 72570 41112
rect 72424 41074 72476 41080
rect 72332 41064 72384 41070
rect 72330 41032 72332 41041
rect 72384 41032 72386 41041
rect 72528 41002 72556 41103
rect 72330 40967 72386 40976
rect 72516 40996 72568 41002
rect 72516 40938 72568 40944
rect 72620 40526 72648 41414
rect 72712 41138 72740 42026
rect 72792 41608 72844 41614
rect 72792 41550 72844 41556
rect 72804 41274 72832 41550
rect 72792 41268 72844 41274
rect 72792 41210 72844 41216
rect 72700 41132 72752 41138
rect 72700 41074 72752 41080
rect 72424 40520 72476 40526
rect 72424 40462 72476 40468
rect 72608 40520 72660 40526
rect 72608 40462 72660 40468
rect 72436 40186 72464 40462
rect 72424 40180 72476 40186
rect 72424 40122 72476 40128
rect 72148 39976 72200 39982
rect 72148 39918 72200 39924
rect 72516 39976 72568 39982
rect 72516 39918 72568 39924
rect 71964 39636 72016 39642
rect 71964 39578 72016 39584
rect 71780 39500 71832 39506
rect 71780 39442 71832 39448
rect 71976 39438 72004 39578
rect 72160 39506 72188 39918
rect 72528 39642 72556 39918
rect 72620 39914 72648 40462
rect 72608 39908 72660 39914
rect 72608 39850 72660 39856
rect 72516 39636 72568 39642
rect 72516 39578 72568 39584
rect 72148 39500 72200 39506
rect 72148 39442 72200 39448
rect 71964 39432 72016 39438
rect 71964 39374 72016 39380
rect 71976 38962 72004 39374
rect 72424 39364 72476 39370
rect 72424 39306 72476 39312
rect 71964 38956 72016 38962
rect 71964 38898 72016 38904
rect 71688 38888 71740 38894
rect 71688 38830 71740 38836
rect 71412 38752 71464 38758
rect 71412 38694 71464 38700
rect 72436 38554 72464 39306
rect 73080 39098 73108 48282
rect 81020 47356 81316 47376
rect 81076 47354 81100 47356
rect 81156 47354 81180 47356
rect 81236 47354 81260 47356
rect 81098 47302 81100 47354
rect 81162 47302 81174 47354
rect 81236 47302 81238 47354
rect 81076 47300 81100 47302
rect 81156 47300 81180 47302
rect 81236 47300 81260 47302
rect 81020 47280 81316 47300
rect 90836 46374 90864 49248
rect 96380 47900 96676 47920
rect 96436 47898 96460 47900
rect 96516 47898 96540 47900
rect 96596 47898 96620 47900
rect 96458 47846 96460 47898
rect 96522 47846 96534 47898
rect 96596 47846 96598 47898
rect 96436 47844 96460 47846
rect 96516 47844 96540 47846
rect 96596 47844 96620 47846
rect 96380 47824 96676 47844
rect 96380 46812 96676 46832
rect 96436 46810 96460 46812
rect 96516 46810 96540 46812
rect 96596 46810 96620 46812
rect 96458 46758 96460 46810
rect 96522 46758 96534 46810
rect 96596 46758 96598 46810
rect 96436 46756 96460 46758
rect 96516 46756 96540 46758
rect 96596 46756 96620 46758
rect 96380 46736 96676 46756
rect 83832 46368 83884 46374
rect 83832 46310 83884 46316
rect 90824 46368 90876 46374
rect 90824 46310 90876 46316
rect 81020 46268 81316 46288
rect 81076 46266 81100 46268
rect 81156 46266 81180 46268
rect 81236 46266 81260 46268
rect 81098 46214 81100 46266
rect 81162 46214 81174 46266
rect 81236 46214 81238 46266
rect 81076 46212 81100 46214
rect 81156 46212 81180 46214
rect 81236 46212 81260 46214
rect 81020 46192 81316 46212
rect 81020 45180 81316 45200
rect 81076 45178 81100 45180
rect 81156 45178 81180 45180
rect 81236 45178 81260 45180
rect 81098 45126 81100 45178
rect 81162 45126 81174 45178
rect 81236 45126 81238 45178
rect 81076 45124 81100 45126
rect 81156 45124 81180 45126
rect 81236 45124 81260 45126
rect 81020 45104 81316 45124
rect 73620 44532 73672 44538
rect 73620 44474 73672 44480
rect 73632 42702 73660 44474
rect 77392 44260 77444 44266
rect 77392 44202 77444 44208
rect 77404 43994 77432 44202
rect 81020 44092 81316 44112
rect 81076 44090 81100 44092
rect 81156 44090 81180 44092
rect 81236 44090 81260 44092
rect 81098 44038 81100 44090
rect 81162 44038 81174 44090
rect 81236 44038 81238 44090
rect 81076 44036 81100 44038
rect 81156 44036 81180 44038
rect 81236 44036 81260 44038
rect 81020 44016 81316 44036
rect 77392 43988 77444 43994
rect 77392 43930 77444 43936
rect 73344 42696 73396 42702
rect 73344 42638 73396 42644
rect 73620 42696 73672 42702
rect 73620 42638 73672 42644
rect 73068 39092 73120 39098
rect 73068 39034 73120 39040
rect 73080 38894 73108 39034
rect 72792 38888 72844 38894
rect 72792 38830 72844 38836
rect 73068 38888 73120 38894
rect 73068 38830 73120 38836
rect 72608 38752 72660 38758
rect 72608 38694 72660 38700
rect 72424 38548 72476 38554
rect 72424 38490 72476 38496
rect 71688 38480 71740 38486
rect 71688 38422 71740 38428
rect 70124 38004 70176 38010
rect 70124 37946 70176 37952
rect 70136 37330 70164 37946
rect 71700 37466 71728 38422
rect 72332 38004 72384 38010
rect 72332 37946 72384 37952
rect 72344 37806 72372 37946
rect 72332 37800 72384 37806
rect 72332 37742 72384 37748
rect 72620 37670 72648 38694
rect 72516 37664 72568 37670
rect 72516 37606 72568 37612
rect 72608 37664 72660 37670
rect 72608 37606 72660 37612
rect 71688 37460 71740 37466
rect 71688 37402 71740 37408
rect 70124 37324 70176 37330
rect 70124 37266 70176 37272
rect 71136 37324 71188 37330
rect 71136 37266 71188 37272
rect 71148 36786 71176 37266
rect 71136 36780 71188 36786
rect 71136 36722 71188 36728
rect 71700 35834 71728 37402
rect 72528 37330 72556 37606
rect 72516 37324 72568 37330
rect 72516 37266 72568 37272
rect 72804 36650 72832 38830
rect 73080 38010 73108 38830
rect 73160 38752 73212 38758
rect 73160 38694 73212 38700
rect 73172 38418 73200 38694
rect 73160 38412 73212 38418
rect 73160 38354 73212 38360
rect 73068 38004 73120 38010
rect 73068 37946 73120 37952
rect 73172 37806 73200 38354
rect 73356 38282 73384 42638
rect 73528 40384 73580 40390
rect 73528 40326 73580 40332
rect 73540 39982 73568 40326
rect 73528 39976 73580 39982
rect 73528 39918 73580 39924
rect 73540 38486 73568 39918
rect 73528 38480 73580 38486
rect 73528 38422 73580 38428
rect 73344 38276 73396 38282
rect 73264 38236 73344 38264
rect 73160 37800 73212 37806
rect 73160 37742 73212 37748
rect 73172 37330 73200 37742
rect 73160 37324 73212 37330
rect 73160 37266 73212 37272
rect 72792 36644 72844 36650
rect 72792 36586 72844 36592
rect 72424 36576 72476 36582
rect 72424 36518 72476 36524
rect 71964 36168 72016 36174
rect 71964 36110 72016 36116
rect 71688 35828 71740 35834
rect 71688 35770 71740 35776
rect 71976 35698 72004 36110
rect 71964 35692 72016 35698
rect 71964 35634 72016 35640
rect 72148 35624 72200 35630
rect 72148 35566 72200 35572
rect 72160 35494 72188 35566
rect 72148 35488 72200 35494
rect 72148 35430 72200 35436
rect 72160 35018 72188 35430
rect 72148 35012 72200 35018
rect 72148 34954 72200 34960
rect 69756 34400 69808 34406
rect 70124 34400 70176 34406
rect 69756 34342 69808 34348
rect 70122 34368 70124 34377
rect 70176 34368 70178 34377
rect 69480 33652 69532 33658
rect 69480 33594 69532 33600
rect 69296 33448 69348 33454
rect 69296 33390 69348 33396
rect 68744 33108 68796 33114
rect 68744 33050 68796 33056
rect 69296 33040 69348 33046
rect 69296 32982 69348 32988
rect 68836 32904 68888 32910
rect 68836 32846 68888 32852
rect 68468 31680 68520 31686
rect 68468 31622 68520 31628
rect 68480 31482 68508 31622
rect 68848 31482 68876 32846
rect 69308 32366 69336 32982
rect 69296 32360 69348 32366
rect 69296 32302 69348 32308
rect 69020 31884 69072 31890
rect 69020 31826 69072 31832
rect 69032 31686 69060 31826
rect 69020 31680 69072 31686
rect 69020 31622 69072 31628
rect 68468 31476 68520 31482
rect 68468 31418 68520 31424
rect 68836 31476 68888 31482
rect 68836 31418 68888 31424
rect 68376 31408 68428 31414
rect 68376 31350 68428 31356
rect 69032 31142 69060 31622
rect 69020 31136 69072 31142
rect 69072 31096 69244 31124
rect 69020 31078 69072 31084
rect 69216 30802 69244 31096
rect 69492 30938 69520 33594
rect 69664 33584 69716 33590
rect 69664 33526 69716 33532
rect 69676 32502 69704 33526
rect 69768 33522 69796 34342
rect 70122 34303 70178 34312
rect 72436 34202 72464 36518
rect 72884 36032 72936 36038
rect 72884 35974 72936 35980
rect 72896 35630 72924 35974
rect 72884 35624 72936 35630
rect 72884 35566 72936 35572
rect 72896 35154 72924 35566
rect 72884 35148 72936 35154
rect 72884 35090 72936 35096
rect 72424 34196 72476 34202
rect 72424 34138 72476 34144
rect 73264 34066 73292 38236
rect 73344 38218 73396 38224
rect 73632 37466 73660 42638
rect 77404 41750 77432 43930
rect 79600 43852 79652 43858
rect 79600 43794 79652 43800
rect 77760 43784 77812 43790
rect 77760 43726 77812 43732
rect 77772 43314 77800 43726
rect 77760 43308 77812 43314
rect 77760 43250 77812 43256
rect 77852 43240 77904 43246
rect 77852 43182 77904 43188
rect 78404 43240 78456 43246
rect 78404 43182 78456 43188
rect 78588 43240 78640 43246
rect 78588 43182 78640 43188
rect 77484 43104 77536 43110
rect 77484 43046 77536 43052
rect 77496 42838 77524 43046
rect 77864 42906 77892 43182
rect 77852 42900 77904 42906
rect 77852 42842 77904 42848
rect 77484 42832 77536 42838
rect 77484 42774 77536 42780
rect 77496 42566 77524 42774
rect 78416 42702 78444 43182
rect 78600 42838 78628 43182
rect 78588 42832 78640 42838
rect 78588 42774 78640 42780
rect 78404 42696 78456 42702
rect 78404 42638 78456 42644
rect 77760 42628 77812 42634
rect 77760 42570 77812 42576
rect 77484 42560 77536 42566
rect 77484 42502 77536 42508
rect 77392 41744 77444 41750
rect 77392 41686 77444 41692
rect 74264 41676 74316 41682
rect 74264 41618 74316 41624
rect 77116 41676 77168 41682
rect 77116 41618 77168 41624
rect 74276 40186 74304 41618
rect 76196 41064 76248 41070
rect 76196 41006 76248 41012
rect 76208 40934 76236 41006
rect 76196 40928 76248 40934
rect 76196 40870 76248 40876
rect 76208 40730 76236 40870
rect 76196 40724 76248 40730
rect 76196 40666 76248 40672
rect 74264 40180 74316 40186
rect 74264 40122 74316 40128
rect 77128 39030 77156 41618
rect 77496 41546 77524 42502
rect 77576 42220 77628 42226
rect 77576 42162 77628 42168
rect 77484 41540 77536 41546
rect 77484 41482 77536 41488
rect 77208 41064 77260 41070
rect 77208 41006 77260 41012
rect 77484 41064 77536 41070
rect 77484 41006 77536 41012
rect 77220 40526 77248 41006
rect 77496 40594 77524 41006
rect 77484 40588 77536 40594
rect 77484 40530 77536 40536
rect 77208 40520 77260 40526
rect 77208 40462 77260 40468
rect 77208 39976 77260 39982
rect 77208 39918 77260 39924
rect 77116 39024 77168 39030
rect 77116 38966 77168 38972
rect 77128 38894 77156 38966
rect 77116 38888 77168 38894
rect 77116 38830 77168 38836
rect 77128 38554 77156 38830
rect 76656 38548 76708 38554
rect 76656 38490 76708 38496
rect 77116 38548 77168 38554
rect 77116 38490 77168 38496
rect 76012 38412 76064 38418
rect 76012 38354 76064 38360
rect 73620 37460 73672 37466
rect 73620 37402 73672 37408
rect 75920 36712 75972 36718
rect 75920 36654 75972 36660
rect 73344 36576 73396 36582
rect 73344 36518 73396 36524
rect 75000 36576 75052 36582
rect 75000 36518 75052 36524
rect 73356 36242 73384 36518
rect 73344 36236 73396 36242
rect 73344 36178 73396 36184
rect 73356 36038 73384 36178
rect 73344 36032 73396 36038
rect 73344 35974 73396 35980
rect 74170 35592 74226 35601
rect 74170 35527 74172 35536
rect 74224 35527 74226 35536
rect 74172 35498 74224 35504
rect 75012 35494 75040 36518
rect 75184 36236 75236 36242
rect 75184 36178 75236 36184
rect 75368 36236 75420 36242
rect 75368 36178 75420 36184
rect 75000 35488 75052 35494
rect 75000 35430 75052 35436
rect 75196 35170 75224 36178
rect 75380 35698 75408 36178
rect 75828 36168 75880 36174
rect 75828 36110 75880 36116
rect 75840 35698 75868 36110
rect 75932 35834 75960 36654
rect 76024 36378 76052 38354
rect 76012 36372 76064 36378
rect 76012 36314 76064 36320
rect 75920 35828 75972 35834
rect 75920 35770 75972 35776
rect 75368 35692 75420 35698
rect 75368 35634 75420 35640
rect 75828 35692 75880 35698
rect 75828 35634 75880 35640
rect 75012 35154 75224 35170
rect 75000 35148 75224 35154
rect 75052 35142 75224 35148
rect 75000 35090 75052 35096
rect 75012 34678 75040 35090
rect 75552 35080 75604 35086
rect 75552 35022 75604 35028
rect 75184 35012 75236 35018
rect 75184 34954 75236 34960
rect 75000 34672 75052 34678
rect 75000 34614 75052 34620
rect 75196 34202 75224 34954
rect 75184 34196 75236 34202
rect 75184 34138 75236 34144
rect 75564 34066 75592 35022
rect 75828 34944 75880 34950
rect 75828 34886 75880 34892
rect 75736 34740 75788 34746
rect 75736 34682 75788 34688
rect 75748 34202 75776 34682
rect 75840 34542 75868 34886
rect 75828 34536 75880 34542
rect 75828 34478 75880 34484
rect 75840 34406 75868 34478
rect 75828 34400 75880 34406
rect 75828 34342 75880 34348
rect 75736 34196 75788 34202
rect 75736 34138 75788 34144
rect 73252 34060 73304 34066
rect 73252 34002 73304 34008
rect 74448 34060 74500 34066
rect 74448 34002 74500 34008
rect 75552 34060 75604 34066
rect 75552 34002 75604 34008
rect 74264 33992 74316 33998
rect 74264 33934 74316 33940
rect 73988 33924 74040 33930
rect 73988 33866 74040 33872
rect 69756 33516 69808 33522
rect 69756 33458 69808 33464
rect 74000 32978 74028 33866
rect 74276 32978 74304 33934
rect 74460 32978 74488 34002
rect 75748 33998 75776 34138
rect 75736 33992 75788 33998
rect 75736 33934 75788 33940
rect 75840 33862 75868 34342
rect 75552 33856 75604 33862
rect 75552 33798 75604 33804
rect 75828 33856 75880 33862
rect 75828 33798 75880 33804
rect 75564 33386 75592 33798
rect 75920 33448 75972 33454
rect 75920 33390 75972 33396
rect 75552 33380 75604 33386
rect 75552 33322 75604 33328
rect 75564 33114 75592 33322
rect 75552 33108 75604 33114
rect 75552 33050 75604 33056
rect 73988 32972 74040 32978
rect 73988 32914 74040 32920
rect 74264 32972 74316 32978
rect 74264 32914 74316 32920
rect 74448 32972 74500 32978
rect 74448 32914 74500 32920
rect 74264 32836 74316 32842
rect 74264 32778 74316 32784
rect 69940 32768 69992 32774
rect 69940 32710 69992 32716
rect 69952 32570 69980 32710
rect 69940 32564 69992 32570
rect 69940 32506 69992 32512
rect 69664 32496 69716 32502
rect 69664 32438 69716 32444
rect 74276 32366 74304 32778
rect 74264 32360 74316 32366
rect 74264 32302 74316 32308
rect 74460 32026 74488 32914
rect 75184 32836 75236 32842
rect 75184 32778 75236 32784
rect 74448 32020 74500 32026
rect 74448 31962 74500 31968
rect 75196 31958 75224 32778
rect 75932 32298 75960 33390
rect 76024 33046 76052 36314
rect 76668 36038 76696 38490
rect 77220 37330 77248 39918
rect 77588 39846 77616 42162
rect 77668 42152 77720 42158
rect 77668 42094 77720 42100
rect 77680 41138 77708 42094
rect 77772 42090 77800 42570
rect 77852 42356 77904 42362
rect 77852 42298 77904 42304
rect 77760 42084 77812 42090
rect 77760 42026 77812 42032
rect 77668 41132 77720 41138
rect 77668 41074 77720 41080
rect 77772 40730 77800 42026
rect 77864 41682 77892 42298
rect 77852 41676 77904 41682
rect 77852 41618 77904 41624
rect 78956 41472 79008 41478
rect 78956 41414 79008 41420
rect 78968 40934 78996 41414
rect 78956 40928 79008 40934
rect 78956 40870 79008 40876
rect 77760 40724 77812 40730
rect 77760 40666 77812 40672
rect 77576 39840 77628 39846
rect 77576 39782 77628 39788
rect 77760 39840 77812 39846
rect 77760 39782 77812 39788
rect 77772 39642 77800 39782
rect 77760 39636 77812 39642
rect 77760 39578 77812 39584
rect 78220 39500 78272 39506
rect 78220 39442 78272 39448
rect 77760 39092 77812 39098
rect 77760 39034 77812 39040
rect 77484 38344 77536 38350
rect 77484 38286 77536 38292
rect 77496 38010 77524 38286
rect 77772 38010 77800 39034
rect 78232 38350 78260 39442
rect 78404 39296 78456 39302
rect 78404 39238 78456 39244
rect 78416 38962 78444 39238
rect 78404 38956 78456 38962
rect 78404 38898 78456 38904
rect 79612 38894 79640 43794
rect 79692 43648 79744 43654
rect 79692 43590 79744 43596
rect 79704 42770 79732 43590
rect 81020 43004 81316 43024
rect 81076 43002 81100 43004
rect 81156 43002 81180 43004
rect 81236 43002 81260 43004
rect 81098 42950 81100 43002
rect 81162 42950 81174 43002
rect 81236 42950 81238 43002
rect 81076 42948 81100 42950
rect 81156 42948 81180 42950
rect 81236 42948 81260 42950
rect 81020 42928 81316 42948
rect 79692 42764 79744 42770
rect 79692 42706 79744 42712
rect 82176 42696 82228 42702
rect 82176 42638 82228 42644
rect 79784 42560 79836 42566
rect 79784 42502 79836 42508
rect 79796 41818 79824 42502
rect 81020 41916 81316 41936
rect 81076 41914 81100 41916
rect 81156 41914 81180 41916
rect 81236 41914 81260 41916
rect 81098 41862 81100 41914
rect 81162 41862 81174 41914
rect 81236 41862 81238 41914
rect 81076 41860 81100 41862
rect 81156 41860 81180 41862
rect 81236 41860 81260 41862
rect 81020 41840 81316 41860
rect 79784 41812 79836 41818
rect 79784 41754 79836 41760
rect 81020 40828 81316 40848
rect 81076 40826 81100 40828
rect 81156 40826 81180 40828
rect 81236 40826 81260 40828
rect 81098 40774 81100 40826
rect 81162 40774 81174 40826
rect 81236 40774 81238 40826
rect 81076 40772 81100 40774
rect 81156 40772 81180 40774
rect 81236 40772 81260 40774
rect 81020 40752 81316 40772
rect 79692 40044 79744 40050
rect 79692 39986 79744 39992
rect 79704 39574 79732 39986
rect 82188 39982 82216 42638
rect 83372 41608 83424 41614
rect 83372 41550 83424 41556
rect 83648 41608 83700 41614
rect 83648 41550 83700 41556
rect 83280 40520 83332 40526
rect 83280 40462 83332 40468
rect 83292 40118 83320 40462
rect 83280 40112 83332 40118
rect 83280 40054 83332 40060
rect 82176 39976 82228 39982
rect 82176 39918 82228 39924
rect 82268 39908 82320 39914
rect 82268 39850 82320 39856
rect 81020 39740 81316 39760
rect 81076 39738 81100 39740
rect 81156 39738 81180 39740
rect 81236 39738 81260 39740
rect 81098 39686 81100 39738
rect 81162 39686 81174 39738
rect 81236 39686 81238 39738
rect 81076 39684 81100 39686
rect 81156 39684 81180 39686
rect 81236 39684 81260 39686
rect 81020 39664 81316 39684
rect 79692 39568 79744 39574
rect 79692 39510 79744 39516
rect 79048 38888 79100 38894
rect 79048 38830 79100 38836
rect 79600 38888 79652 38894
rect 79600 38830 79652 38836
rect 79060 38554 79088 38830
rect 79048 38548 79100 38554
rect 79048 38490 79100 38496
rect 79060 38350 79088 38490
rect 79704 38486 79732 39510
rect 82280 38894 82308 39850
rect 82360 39840 82412 39846
rect 82360 39782 82412 39788
rect 82268 38888 82320 38894
rect 82268 38830 82320 38836
rect 79876 38752 79928 38758
rect 79876 38694 79928 38700
rect 79140 38480 79192 38486
rect 79140 38422 79192 38428
rect 79692 38480 79744 38486
rect 79692 38422 79744 38428
rect 78220 38344 78272 38350
rect 78220 38286 78272 38292
rect 79048 38344 79100 38350
rect 79048 38286 79100 38292
rect 78956 38276 79008 38282
rect 78956 38218 79008 38224
rect 78772 38208 78824 38214
rect 78772 38150 78824 38156
rect 77484 38004 77536 38010
rect 77484 37946 77536 37952
rect 77760 38004 77812 38010
rect 77760 37946 77812 37952
rect 77772 37806 77800 37946
rect 77760 37800 77812 37806
rect 77760 37742 77812 37748
rect 78784 37398 78812 38150
rect 78968 37466 78996 38218
rect 78956 37460 79008 37466
rect 78956 37402 79008 37408
rect 78772 37392 78824 37398
rect 78772 37334 78824 37340
rect 77208 37324 77260 37330
rect 77208 37266 77260 37272
rect 77220 36106 77248 37266
rect 78784 36922 78812 37334
rect 78968 37194 78996 37402
rect 78956 37188 79008 37194
rect 78956 37130 79008 37136
rect 79152 36922 79180 38422
rect 79784 38412 79836 38418
rect 79784 38354 79836 38360
rect 79416 38276 79468 38282
rect 79416 38218 79468 38224
rect 79324 37732 79376 37738
rect 79324 37674 79376 37680
rect 79336 37398 79364 37674
rect 79428 37670 79456 38218
rect 79796 37806 79824 38354
rect 79888 37874 79916 38694
rect 81020 38652 81316 38672
rect 81076 38650 81100 38652
rect 81156 38650 81180 38652
rect 81236 38650 81260 38652
rect 81098 38598 81100 38650
rect 81162 38598 81174 38650
rect 81236 38598 81238 38650
rect 81076 38596 81100 38598
rect 81156 38596 81180 38598
rect 81236 38596 81260 38598
rect 81020 38576 81316 38596
rect 79968 38548 80020 38554
rect 79968 38490 80020 38496
rect 79980 38214 80008 38490
rect 80336 38412 80388 38418
rect 80336 38354 80388 38360
rect 80888 38412 80940 38418
rect 80888 38354 80940 38360
rect 79968 38208 80020 38214
rect 79968 38150 80020 38156
rect 79876 37868 79928 37874
rect 79876 37810 79928 37816
rect 79784 37800 79836 37806
rect 79784 37742 79836 37748
rect 79416 37664 79468 37670
rect 79416 37606 79468 37612
rect 79324 37392 79376 37398
rect 79324 37334 79376 37340
rect 79888 37330 79916 37810
rect 79980 37806 80008 38150
rect 79968 37800 80020 37806
rect 79968 37742 80020 37748
rect 80348 37738 80376 38354
rect 80336 37732 80388 37738
rect 80336 37674 80388 37680
rect 79876 37324 79928 37330
rect 79876 37266 79928 37272
rect 79692 37256 79744 37262
rect 79692 37198 79744 37204
rect 79784 37256 79836 37262
rect 79784 37198 79836 37204
rect 78772 36916 78824 36922
rect 78772 36858 78824 36864
rect 79140 36916 79192 36922
rect 79140 36858 79192 36864
rect 79704 36650 79732 37198
rect 79796 36854 79824 37198
rect 79968 37120 80020 37126
rect 79968 37062 80020 37068
rect 79876 36916 79928 36922
rect 79876 36858 79928 36864
rect 79784 36848 79836 36854
rect 79784 36790 79836 36796
rect 79692 36644 79744 36650
rect 79692 36586 79744 36592
rect 79888 36242 79916 36858
rect 79980 36854 80008 37062
rect 79968 36848 80020 36854
rect 79968 36790 80020 36796
rect 80348 36786 80376 37674
rect 80900 37398 80928 38354
rect 81020 37564 81316 37584
rect 81076 37562 81100 37564
rect 81156 37562 81180 37564
rect 81236 37562 81260 37564
rect 81098 37510 81100 37562
rect 81162 37510 81174 37562
rect 81236 37510 81238 37562
rect 81076 37508 81100 37510
rect 81156 37508 81180 37510
rect 81236 37508 81260 37510
rect 81020 37488 81316 37508
rect 80888 37392 80940 37398
rect 80888 37334 80940 37340
rect 81348 37324 81400 37330
rect 81348 37266 81400 37272
rect 80428 37120 80480 37126
rect 80428 37062 80480 37068
rect 80336 36780 80388 36786
rect 80336 36722 80388 36728
rect 80440 36242 80468 37062
rect 81020 36476 81316 36496
rect 81076 36474 81100 36476
rect 81156 36474 81180 36476
rect 81236 36474 81260 36476
rect 81098 36422 81100 36474
rect 81162 36422 81174 36474
rect 81236 36422 81238 36474
rect 81076 36420 81100 36422
rect 81156 36420 81180 36422
rect 81236 36420 81260 36422
rect 81020 36400 81316 36420
rect 79876 36236 79928 36242
rect 79876 36178 79928 36184
rect 80428 36236 80480 36242
rect 80428 36178 80480 36184
rect 77208 36100 77260 36106
rect 77208 36042 77260 36048
rect 76656 36032 76708 36038
rect 76656 35974 76708 35980
rect 77024 35828 77076 35834
rect 77024 35770 77076 35776
rect 77036 35154 77064 35770
rect 77220 35154 77248 36042
rect 79508 36032 79560 36038
rect 79508 35974 79560 35980
rect 80244 36032 80296 36038
rect 80244 35974 80296 35980
rect 77300 35488 77352 35494
rect 77300 35430 77352 35436
rect 77024 35148 77076 35154
rect 77024 35090 77076 35096
rect 77208 35148 77260 35154
rect 77208 35090 77260 35096
rect 76840 34944 76892 34950
rect 76840 34886 76892 34892
rect 76852 34474 76880 34886
rect 77024 34740 77076 34746
rect 77024 34682 77076 34688
rect 77036 34542 77064 34682
rect 77116 34604 77168 34610
rect 77116 34546 77168 34552
rect 77024 34536 77076 34542
rect 77024 34478 77076 34484
rect 76840 34468 76892 34474
rect 76840 34410 76892 34416
rect 76288 34400 76340 34406
rect 76286 34368 76288 34377
rect 76340 34368 76342 34377
rect 76286 34303 76342 34312
rect 76852 33930 76880 34410
rect 77128 34134 77156 34546
rect 77116 34128 77168 34134
rect 77116 34070 77168 34076
rect 77220 33930 77248 35090
rect 76840 33924 76892 33930
rect 76840 33866 76892 33872
rect 77208 33924 77260 33930
rect 77208 33866 77260 33872
rect 77312 33454 77340 35430
rect 79520 35290 79548 35974
rect 80256 35698 80284 35974
rect 81360 35834 81388 37266
rect 81440 36712 81492 36718
rect 81440 36654 81492 36660
rect 81348 35828 81400 35834
rect 81348 35770 81400 35776
rect 80244 35692 80296 35698
rect 80244 35634 80296 35640
rect 81452 35630 81480 36654
rect 81440 35624 81492 35630
rect 81440 35566 81492 35572
rect 81020 35388 81316 35408
rect 81076 35386 81100 35388
rect 81156 35386 81180 35388
rect 81236 35386 81260 35388
rect 81098 35334 81100 35386
rect 81162 35334 81174 35386
rect 81236 35334 81238 35386
rect 81076 35332 81100 35334
rect 81156 35332 81180 35334
rect 81236 35332 81260 35334
rect 81020 35312 81316 35332
rect 79508 35284 79560 35290
rect 79508 35226 79560 35232
rect 81020 34300 81316 34320
rect 81076 34298 81100 34300
rect 81156 34298 81180 34300
rect 81236 34298 81260 34300
rect 81098 34246 81100 34298
rect 81162 34246 81174 34298
rect 81236 34246 81238 34298
rect 81076 34244 81100 34246
rect 81156 34244 81180 34246
rect 81236 34244 81260 34246
rect 81020 34224 81316 34244
rect 78680 33992 78732 33998
rect 78680 33934 78732 33940
rect 77484 33856 77536 33862
rect 77484 33798 77536 33804
rect 77496 33522 77524 33798
rect 77484 33516 77536 33522
rect 77484 33458 77536 33464
rect 77300 33448 77352 33454
rect 77300 33390 77352 33396
rect 77760 33448 77812 33454
rect 77760 33390 77812 33396
rect 77392 33312 77444 33318
rect 77392 33254 77444 33260
rect 76012 33040 76064 33046
rect 76012 32982 76064 32988
rect 77404 32978 77432 33254
rect 77772 33114 77800 33390
rect 77760 33108 77812 33114
rect 77760 33050 77812 33056
rect 77392 32972 77444 32978
rect 77392 32914 77444 32920
rect 76012 32496 76064 32502
rect 76012 32438 76064 32444
rect 75920 32292 75972 32298
rect 75920 32234 75972 32240
rect 75552 32224 75604 32230
rect 75552 32166 75604 32172
rect 75184 31952 75236 31958
rect 75184 31894 75236 31900
rect 75564 31890 75592 32166
rect 75552 31884 75604 31890
rect 75552 31826 75604 31832
rect 75736 31884 75788 31890
rect 75736 31826 75788 31832
rect 75748 31482 75776 31826
rect 75736 31476 75788 31482
rect 75736 31418 75788 31424
rect 73620 31408 73672 31414
rect 73620 31350 73672 31356
rect 72516 31204 72568 31210
rect 72516 31146 72568 31152
rect 69480 30932 69532 30938
rect 69480 30874 69532 30880
rect 69756 30932 69808 30938
rect 69756 30874 69808 30880
rect 67732 30796 67784 30802
rect 67732 30738 67784 30744
rect 69204 30796 69256 30802
rect 69204 30738 69256 30744
rect 67744 30598 67772 30738
rect 68008 30728 68060 30734
rect 68008 30670 68060 30676
rect 68020 30598 68048 30670
rect 69664 30660 69716 30666
rect 69664 30602 69716 30608
rect 67732 30592 67784 30598
rect 67732 30534 67784 30540
rect 68008 30592 68060 30598
rect 68008 30534 68060 30540
rect 67744 30394 67772 30534
rect 69676 30394 69704 30602
rect 69768 30598 69796 30874
rect 72528 30870 72556 31146
rect 73632 31142 73660 31350
rect 73620 31136 73672 31142
rect 73620 31078 73672 31084
rect 70032 30864 70084 30870
rect 70032 30806 70084 30812
rect 72516 30864 72568 30870
rect 72516 30806 72568 30812
rect 70044 30598 70072 30806
rect 73160 30728 73212 30734
rect 73160 30670 73212 30676
rect 73172 30598 73200 30670
rect 69756 30592 69808 30598
rect 69756 30534 69808 30540
rect 70032 30592 70084 30598
rect 70032 30534 70084 30540
rect 73160 30592 73212 30598
rect 73160 30534 73212 30540
rect 70044 30394 70072 30534
rect 67732 30388 67784 30394
rect 67732 30330 67784 30336
rect 69664 30388 69716 30394
rect 69664 30330 69716 30336
rect 70032 30388 70084 30394
rect 70032 30330 70084 30336
rect 71596 30320 71648 30326
rect 71596 30262 71648 30268
rect 68836 30184 68888 30190
rect 68836 30126 68888 30132
rect 68848 30054 68876 30126
rect 67916 30048 67968 30054
rect 67916 29990 67968 29996
rect 68836 30048 68888 30054
rect 68836 29990 68888 29996
rect 67640 29844 67692 29850
rect 67640 29786 67692 29792
rect 67652 29646 67680 29786
rect 67928 29714 67956 29990
rect 67916 29708 67968 29714
rect 67916 29650 67968 29656
rect 67640 29640 67692 29646
rect 67640 29582 67692 29588
rect 68848 29510 68876 29990
rect 69480 29844 69532 29850
rect 69480 29786 69532 29792
rect 67916 29504 67968 29510
rect 67916 29446 67968 29452
rect 68836 29504 68888 29510
rect 68836 29446 68888 29452
rect 66076 29300 66128 29306
rect 66076 29242 66128 29248
rect 63500 29232 63552 29238
rect 63500 29174 63552 29180
rect 61568 29164 61620 29170
rect 61568 29106 61620 29112
rect 63512 26586 63540 29174
rect 67928 27946 67956 29446
rect 69492 29238 69520 29786
rect 71608 29646 71636 30262
rect 73172 30258 73200 30534
rect 73160 30252 73212 30258
rect 73160 30194 73212 30200
rect 73160 30048 73212 30054
rect 73160 29990 73212 29996
rect 73172 29850 73200 29990
rect 73160 29844 73212 29850
rect 73160 29786 73212 29792
rect 71596 29640 71648 29646
rect 71596 29582 71648 29588
rect 69480 29232 69532 29238
rect 69480 29174 69532 29180
rect 73632 29170 73660 31078
rect 73724 30802 74304 30818
rect 73712 30796 74316 30802
rect 73764 30790 74264 30796
rect 73712 30738 73764 30744
rect 74264 30738 74316 30744
rect 74356 30184 74408 30190
rect 74356 30126 74408 30132
rect 74368 29850 74396 30126
rect 75932 30122 75960 32234
rect 76024 32026 76052 32438
rect 76012 32020 76064 32026
rect 76012 31962 76064 31968
rect 76024 31482 76052 31962
rect 78692 31890 78720 33934
rect 81020 33212 81316 33232
rect 81076 33210 81100 33212
rect 81156 33210 81180 33212
rect 81236 33210 81260 33212
rect 81098 33158 81100 33210
rect 81162 33158 81174 33210
rect 81236 33158 81238 33210
rect 81076 33156 81100 33158
rect 81156 33156 81180 33158
rect 81236 33156 81260 33158
rect 81020 33136 81316 33156
rect 80520 32972 80572 32978
rect 80520 32914 80572 32920
rect 80532 32434 80560 32914
rect 80520 32428 80572 32434
rect 80520 32370 80572 32376
rect 78680 31884 78732 31890
rect 78680 31826 78732 31832
rect 79784 31884 79836 31890
rect 79784 31826 79836 31832
rect 76012 31476 76064 31482
rect 76012 31418 76064 31424
rect 79600 31476 79652 31482
rect 79600 31418 79652 31424
rect 76024 30870 76052 31418
rect 76012 30864 76064 30870
rect 76012 30806 76064 30812
rect 79612 30802 79640 31418
rect 79796 31278 79824 31826
rect 80532 31686 80560 32370
rect 80888 32224 80940 32230
rect 80888 32166 80940 32172
rect 80900 32026 80928 32166
rect 81020 32124 81316 32144
rect 81076 32122 81100 32124
rect 81156 32122 81180 32124
rect 81236 32122 81260 32124
rect 81098 32070 81100 32122
rect 81162 32070 81174 32122
rect 81236 32070 81238 32122
rect 81076 32068 81100 32070
rect 81156 32068 81180 32070
rect 81236 32068 81260 32070
rect 81020 32048 81316 32068
rect 81452 32026 81480 35566
rect 81532 33448 81584 33454
rect 81532 33390 81584 33396
rect 81544 32434 81572 33390
rect 82268 33312 82320 33318
rect 82268 33254 82320 33260
rect 82280 33046 82308 33254
rect 82268 33040 82320 33046
rect 82268 32982 82320 32988
rect 82372 32978 82400 39782
rect 83384 39642 83412 41550
rect 83660 40662 83688 41550
rect 83740 41200 83792 41206
rect 83740 41142 83792 41148
rect 83648 40656 83700 40662
rect 83648 40598 83700 40604
rect 83752 40594 83780 41142
rect 83556 40588 83608 40594
rect 83556 40530 83608 40536
rect 83740 40588 83792 40594
rect 83740 40530 83792 40536
rect 83568 40050 83596 40530
rect 83752 40186 83780 40530
rect 83740 40180 83792 40186
rect 83740 40122 83792 40128
rect 83556 40044 83608 40050
rect 83556 39986 83608 39992
rect 83752 39982 83780 40122
rect 83740 39976 83792 39982
rect 83740 39918 83792 39924
rect 83372 39636 83424 39642
rect 83372 39578 83424 39584
rect 83372 38752 83424 38758
rect 83372 38694 83424 38700
rect 83384 38554 83412 38694
rect 83372 38548 83424 38554
rect 83372 38490 83424 38496
rect 83384 38214 83412 38490
rect 83372 38208 83424 38214
rect 83372 38150 83424 38156
rect 82912 34196 82964 34202
rect 82912 34138 82964 34144
rect 82544 33040 82596 33046
rect 82544 32982 82596 32988
rect 82360 32972 82412 32978
rect 82360 32914 82412 32920
rect 82452 32904 82504 32910
rect 82452 32846 82504 32852
rect 82084 32836 82136 32842
rect 82084 32778 82136 32784
rect 82096 32434 82124 32778
rect 81532 32428 81584 32434
rect 81532 32370 81584 32376
rect 82084 32428 82136 32434
rect 82084 32370 82136 32376
rect 82464 32366 82492 32846
rect 82556 32774 82584 32982
rect 82544 32768 82596 32774
rect 82544 32710 82596 32716
rect 82556 32434 82584 32710
rect 82544 32428 82596 32434
rect 82544 32370 82596 32376
rect 82452 32360 82504 32366
rect 82452 32302 82504 32308
rect 82728 32292 82780 32298
rect 82728 32234 82780 32240
rect 80888 32020 80940 32026
rect 80888 31962 80940 31968
rect 81440 32020 81492 32026
rect 81440 31962 81492 31968
rect 82268 31952 82320 31958
rect 82268 31894 82320 31900
rect 80888 31816 80940 31822
rect 80888 31758 80940 31764
rect 80520 31680 80572 31686
rect 80520 31622 80572 31628
rect 79784 31272 79836 31278
rect 79784 31214 79836 31220
rect 79876 31272 79928 31278
rect 79876 31214 79928 31220
rect 79600 30796 79652 30802
rect 79600 30738 79652 30744
rect 79796 30734 79824 31214
rect 79888 30802 79916 31214
rect 80900 30802 80928 31758
rect 82280 31362 82308 31894
rect 82740 31414 82768 32234
rect 82820 31816 82872 31822
rect 82820 31758 82872 31764
rect 82728 31408 82780 31414
rect 82280 31334 82400 31362
rect 82728 31350 82780 31356
rect 82372 31278 82400 31334
rect 82740 31278 82768 31350
rect 82360 31272 82412 31278
rect 82360 31214 82412 31220
rect 82728 31272 82780 31278
rect 82728 31214 82780 31220
rect 81020 31036 81316 31056
rect 81076 31034 81100 31036
rect 81156 31034 81180 31036
rect 81236 31034 81260 31036
rect 81098 30982 81100 31034
rect 81162 30982 81174 31034
rect 81236 30982 81238 31034
rect 81076 30980 81100 30982
rect 81156 30980 81180 30982
rect 81236 30980 81260 30982
rect 81020 30960 81316 30980
rect 79876 30796 79928 30802
rect 79876 30738 79928 30744
rect 80888 30796 80940 30802
rect 80888 30738 80940 30744
rect 79784 30728 79836 30734
rect 79784 30670 79836 30676
rect 80704 30728 80756 30734
rect 80704 30670 80756 30676
rect 79232 30592 79284 30598
rect 79232 30534 79284 30540
rect 75920 30116 75972 30122
rect 75920 30058 75972 30064
rect 74356 29844 74408 29850
rect 74356 29786 74408 29792
rect 75932 29646 75960 30058
rect 79244 29714 79272 30534
rect 80716 30394 80744 30670
rect 82372 30666 82400 31214
rect 82832 30870 82860 31758
rect 82820 30864 82872 30870
rect 82820 30806 82872 30812
rect 82360 30660 82412 30666
rect 82360 30602 82412 30608
rect 80704 30388 80756 30394
rect 80704 30330 80756 30336
rect 80060 30184 80112 30190
rect 80060 30126 80112 30132
rect 80072 29850 80100 30126
rect 80520 30048 80572 30054
rect 80520 29990 80572 29996
rect 80060 29844 80112 29850
rect 80060 29786 80112 29792
rect 80532 29714 80560 29990
rect 80716 29850 80744 30330
rect 81020 29948 81316 29968
rect 81076 29946 81100 29948
rect 81156 29946 81180 29948
rect 81236 29946 81260 29948
rect 81098 29894 81100 29946
rect 81162 29894 81174 29946
rect 81236 29894 81238 29946
rect 81076 29892 81100 29894
rect 81156 29892 81180 29894
rect 81236 29892 81260 29894
rect 81020 29872 81316 29892
rect 80704 29844 80756 29850
rect 80704 29786 80756 29792
rect 79232 29708 79284 29714
rect 79232 29650 79284 29656
rect 80520 29708 80572 29714
rect 80520 29650 80572 29656
rect 75920 29640 75972 29646
rect 75920 29582 75972 29588
rect 82924 29578 82952 34138
rect 83188 33856 83240 33862
rect 83188 33798 83240 33804
rect 83200 33522 83228 33798
rect 83188 33516 83240 33522
rect 83188 33458 83240 33464
rect 83200 30870 83228 33458
rect 83188 30864 83240 30870
rect 83188 30806 83240 30812
rect 82912 29572 82964 29578
rect 82912 29514 82964 29520
rect 73620 29164 73672 29170
rect 73620 29106 73672 29112
rect 67916 27940 67968 27946
rect 67916 27882 67968 27888
rect 63500 26580 63552 26586
rect 63500 26522 63552 26528
rect 83844 26081 83872 46310
rect 96380 45724 96676 45744
rect 96436 45722 96460 45724
rect 96516 45722 96540 45724
rect 96596 45722 96620 45724
rect 96458 45670 96460 45722
rect 96522 45670 96534 45722
rect 96596 45670 96598 45722
rect 96436 45668 96460 45670
rect 96516 45668 96540 45670
rect 96596 45668 96620 45670
rect 96380 45648 96676 45668
rect 96380 44636 96676 44656
rect 96436 44634 96460 44636
rect 96516 44634 96540 44636
rect 96596 44634 96620 44636
rect 96458 44582 96460 44634
rect 96522 44582 96534 44634
rect 96596 44582 96598 44634
rect 96436 44580 96460 44582
rect 96516 44580 96540 44582
rect 96596 44580 96620 44582
rect 96380 44560 96676 44580
rect 96380 43548 96676 43568
rect 96436 43546 96460 43548
rect 96516 43546 96540 43548
rect 96596 43546 96620 43548
rect 96458 43494 96460 43546
rect 96522 43494 96534 43546
rect 96596 43494 96598 43546
rect 96436 43492 96460 43494
rect 96516 43492 96540 43494
rect 96596 43492 96620 43494
rect 96380 43472 96676 43492
rect 96380 42460 96676 42480
rect 96436 42458 96460 42460
rect 96516 42458 96540 42460
rect 96596 42458 96620 42460
rect 96458 42406 96460 42458
rect 96522 42406 96534 42458
rect 96596 42406 96598 42458
rect 96436 42404 96460 42406
rect 96516 42404 96540 42406
rect 96596 42404 96620 42406
rect 96380 42384 96676 42404
rect 84568 41472 84620 41478
rect 84568 41414 84620 41420
rect 84108 40996 84160 41002
rect 84108 40938 84160 40944
rect 84120 40730 84148 40938
rect 84108 40724 84160 40730
rect 84108 40666 84160 40672
rect 84120 36582 84148 40666
rect 84580 40594 84608 41414
rect 96380 41372 96676 41392
rect 96436 41370 96460 41372
rect 96516 41370 96540 41372
rect 96596 41370 96620 41372
rect 96458 41318 96460 41370
rect 96522 41318 96534 41370
rect 96596 41318 96598 41370
rect 96436 41316 96460 41318
rect 96516 41316 96540 41318
rect 96596 41316 96620 41318
rect 96380 41296 96676 41316
rect 84568 40588 84620 40594
rect 84568 40530 84620 40536
rect 96380 40284 96676 40304
rect 96436 40282 96460 40284
rect 96516 40282 96540 40284
rect 96596 40282 96620 40284
rect 96458 40230 96460 40282
rect 96522 40230 96534 40282
rect 96596 40230 96598 40282
rect 96436 40228 96460 40230
rect 96516 40228 96540 40230
rect 96596 40228 96620 40230
rect 96380 40208 96676 40228
rect 86316 39500 86368 39506
rect 86316 39442 86368 39448
rect 84384 39432 84436 39438
rect 84384 39374 84436 39380
rect 84396 39098 84424 39374
rect 85396 39296 85448 39302
rect 85396 39238 85448 39244
rect 84384 39092 84436 39098
rect 84384 39034 84436 39040
rect 85408 38894 85436 39238
rect 86328 39098 86356 39442
rect 96380 39196 96676 39216
rect 96436 39194 96460 39196
rect 96516 39194 96540 39196
rect 96596 39194 96620 39196
rect 96458 39142 96460 39194
rect 96522 39142 96534 39194
rect 96596 39142 96598 39194
rect 96436 39140 96460 39142
rect 96516 39140 96540 39142
rect 96596 39140 96620 39142
rect 96380 39120 96676 39140
rect 86316 39092 86368 39098
rect 86316 39034 86368 39040
rect 86328 38894 86356 39034
rect 84292 38888 84344 38894
rect 84292 38830 84344 38836
rect 85396 38888 85448 38894
rect 85396 38830 85448 38836
rect 86316 38888 86368 38894
rect 86316 38830 86368 38836
rect 86776 38888 86828 38894
rect 86776 38830 86828 38836
rect 84304 38486 84332 38830
rect 84752 38820 84804 38826
rect 84752 38762 84804 38768
rect 84292 38480 84344 38486
rect 84292 38422 84344 38428
rect 84200 38344 84252 38350
rect 84200 38286 84252 38292
rect 84212 37670 84240 38286
rect 84200 37664 84252 37670
rect 84200 37606 84252 37612
rect 84212 37466 84240 37606
rect 84200 37460 84252 37466
rect 84200 37402 84252 37408
rect 84764 36922 84792 38762
rect 85396 38276 85448 38282
rect 85396 38218 85448 38224
rect 85408 36922 85436 38218
rect 85580 37936 85632 37942
rect 85580 37878 85632 37884
rect 85592 37398 85620 37878
rect 85580 37392 85632 37398
rect 85580 37334 85632 37340
rect 85856 37324 85908 37330
rect 85856 37266 85908 37272
rect 85948 37324 86000 37330
rect 85948 37266 86000 37272
rect 85764 37256 85816 37262
rect 85764 37198 85816 37204
rect 84752 36916 84804 36922
rect 85396 36916 85448 36922
rect 84752 36858 84804 36864
rect 85224 36876 85396 36904
rect 84108 36576 84160 36582
rect 84108 36518 84160 36524
rect 85028 34536 85080 34542
rect 85028 34478 85080 34484
rect 85040 34134 85068 34478
rect 85028 34128 85080 34134
rect 85028 34070 85080 34076
rect 85224 33114 85252 36876
rect 85396 36858 85448 36864
rect 85488 36848 85540 36854
rect 85488 36790 85540 36796
rect 85304 36576 85356 36582
rect 85304 36518 85356 36524
rect 85316 35698 85344 36518
rect 85500 35766 85528 36790
rect 85776 36106 85804 37198
rect 85868 36310 85896 37266
rect 85960 36922 85988 37266
rect 85948 36916 86000 36922
rect 85948 36858 86000 36864
rect 85960 36378 85988 36858
rect 85948 36372 86000 36378
rect 85948 36314 86000 36320
rect 85856 36304 85908 36310
rect 85856 36246 85908 36252
rect 85764 36100 85816 36106
rect 85764 36042 85816 36048
rect 85488 35760 85540 35766
rect 85488 35702 85540 35708
rect 85304 35692 85356 35698
rect 85304 35634 85356 35640
rect 85316 35578 85344 35634
rect 85316 35550 85436 35578
rect 85408 34678 85436 35550
rect 85396 34672 85448 34678
rect 85396 34614 85448 34620
rect 85212 33108 85264 33114
rect 85212 33050 85264 33056
rect 85028 32904 85080 32910
rect 85028 32846 85080 32852
rect 84200 31476 84252 31482
rect 84200 31418 84252 31424
rect 83924 30864 83976 30870
rect 83924 30806 83976 30812
rect 83936 30734 83964 30806
rect 84212 30802 84240 31418
rect 85040 31414 85068 32846
rect 85408 32230 85436 34614
rect 85500 34542 85528 35702
rect 85868 35698 85896 36246
rect 86328 36038 86356 38830
rect 86788 38010 86816 38830
rect 96380 38108 96676 38128
rect 96436 38106 96460 38108
rect 96516 38106 96540 38108
rect 96596 38106 96620 38108
rect 96458 38054 96460 38106
rect 96522 38054 96534 38106
rect 96596 38054 96598 38106
rect 96436 38052 96460 38054
rect 96516 38052 96540 38054
rect 96596 38052 96620 38054
rect 96380 38032 96676 38052
rect 86776 38004 86828 38010
rect 86776 37946 86828 37952
rect 86592 37800 86644 37806
rect 86592 37742 86644 37748
rect 86604 36922 86632 37742
rect 87328 37324 87380 37330
rect 87328 37266 87380 37272
rect 86592 36916 86644 36922
rect 86592 36858 86644 36864
rect 86776 36916 86828 36922
rect 86776 36858 86828 36864
rect 86788 36310 86816 36858
rect 86960 36712 87012 36718
rect 86880 36660 86960 36666
rect 86880 36654 87012 36660
rect 86880 36638 87000 36654
rect 86880 36378 86908 36638
rect 86868 36372 86920 36378
rect 86868 36314 86920 36320
rect 87340 36310 87368 37266
rect 88432 37120 88484 37126
rect 88432 37062 88484 37068
rect 88444 36718 88472 37062
rect 96380 37020 96676 37040
rect 96436 37018 96460 37020
rect 96516 37018 96540 37020
rect 96596 37018 96620 37020
rect 96458 36966 96460 37018
rect 96522 36966 96534 37018
rect 96596 36966 96598 37018
rect 96436 36964 96460 36966
rect 96516 36964 96540 36966
rect 96596 36964 96620 36966
rect 96380 36944 96676 36964
rect 88432 36712 88484 36718
rect 88432 36654 88484 36660
rect 87880 36644 87932 36650
rect 87880 36586 87932 36592
rect 88340 36644 88392 36650
rect 88340 36586 88392 36592
rect 88708 36644 88760 36650
rect 88708 36586 88760 36592
rect 86776 36304 86828 36310
rect 86776 36246 86828 36252
rect 87328 36304 87380 36310
rect 87328 36246 87380 36252
rect 86316 36032 86368 36038
rect 86316 35974 86368 35980
rect 85856 35692 85908 35698
rect 85856 35634 85908 35640
rect 86776 35556 86828 35562
rect 86776 35498 86828 35504
rect 85488 34536 85540 34542
rect 85488 34478 85540 34484
rect 85488 33992 85540 33998
rect 85488 33934 85540 33940
rect 85500 33658 85528 33934
rect 85488 33652 85540 33658
rect 85488 33594 85540 33600
rect 85672 33448 85724 33454
rect 85672 33390 85724 33396
rect 85684 33046 85712 33390
rect 86788 33386 86816 35498
rect 87340 35154 87368 36246
rect 87892 35630 87920 36586
rect 87972 36576 88024 36582
rect 87972 36518 88024 36524
rect 87984 36106 88012 36518
rect 88064 36168 88116 36174
rect 88064 36110 88116 36116
rect 87972 36100 88024 36106
rect 87972 36042 88024 36048
rect 87880 35624 87932 35630
rect 87880 35566 87932 35572
rect 87892 35290 87920 35566
rect 87880 35284 87932 35290
rect 87880 35226 87932 35232
rect 87328 35148 87380 35154
rect 87328 35090 87380 35096
rect 87144 34468 87196 34474
rect 87144 34410 87196 34416
rect 87156 34066 87184 34410
rect 87984 34202 88012 36042
rect 88076 35630 88104 36110
rect 88352 35698 88380 36586
rect 88720 36242 88748 36586
rect 88708 36236 88760 36242
rect 88708 36178 88760 36184
rect 96380 35932 96676 35952
rect 96436 35930 96460 35932
rect 96516 35930 96540 35932
rect 96596 35930 96620 35932
rect 96458 35878 96460 35930
rect 96522 35878 96534 35930
rect 96596 35878 96598 35930
rect 96436 35876 96460 35878
rect 96516 35876 96540 35878
rect 96596 35876 96620 35878
rect 96380 35856 96676 35876
rect 88340 35692 88392 35698
rect 88340 35634 88392 35640
rect 88064 35624 88116 35630
rect 88064 35566 88116 35572
rect 96380 34844 96676 34864
rect 96436 34842 96460 34844
rect 96516 34842 96540 34844
rect 96596 34842 96620 34844
rect 96458 34790 96460 34842
rect 96522 34790 96534 34842
rect 96596 34790 96598 34842
rect 96436 34788 96460 34790
rect 96516 34788 96540 34790
rect 96596 34788 96620 34790
rect 96380 34768 96676 34788
rect 89812 34536 89864 34542
rect 89812 34478 89864 34484
rect 88524 34468 88576 34474
rect 88524 34410 88576 34416
rect 88340 34400 88392 34406
rect 88340 34342 88392 34348
rect 87972 34196 88024 34202
rect 87972 34138 88024 34144
rect 87144 34060 87196 34066
rect 87144 34002 87196 34008
rect 87420 34060 87472 34066
rect 87420 34002 87472 34008
rect 87156 33658 87184 34002
rect 87236 33856 87288 33862
rect 87236 33798 87288 33804
rect 87144 33652 87196 33658
rect 87144 33594 87196 33600
rect 86776 33380 86828 33386
rect 86776 33322 86828 33328
rect 86684 33312 86736 33318
rect 86684 33254 86736 33260
rect 85672 33040 85724 33046
rect 85672 32982 85724 32988
rect 86696 32978 86724 33254
rect 86788 32978 86816 33322
rect 87248 33046 87276 33798
rect 87236 33040 87288 33046
rect 87236 32982 87288 32988
rect 86684 32972 86736 32978
rect 86684 32914 86736 32920
rect 86776 32972 86828 32978
rect 86776 32914 86828 32920
rect 85580 32768 85632 32774
rect 85580 32710 85632 32716
rect 85592 32502 85620 32710
rect 86960 32564 87012 32570
rect 86960 32506 87012 32512
rect 85580 32496 85632 32502
rect 85580 32438 85632 32444
rect 85396 32224 85448 32230
rect 85396 32166 85448 32172
rect 86972 31890 87000 32506
rect 85396 31884 85448 31890
rect 85396 31826 85448 31832
rect 86960 31884 87012 31890
rect 86960 31826 87012 31832
rect 85120 31680 85172 31686
rect 85120 31622 85172 31628
rect 85132 31482 85160 31622
rect 85120 31476 85172 31482
rect 85120 31418 85172 31424
rect 85028 31408 85080 31414
rect 85028 31350 85080 31356
rect 85132 30938 85160 31418
rect 85408 31210 85436 31826
rect 87432 31278 87460 34002
rect 88352 33930 88380 34342
rect 88536 34066 88564 34410
rect 89824 34066 89852 34478
rect 88432 34060 88484 34066
rect 88432 34002 88484 34008
rect 88524 34060 88576 34066
rect 88524 34002 88576 34008
rect 89812 34060 89864 34066
rect 89812 34002 89864 34008
rect 88340 33924 88392 33930
rect 88340 33866 88392 33872
rect 87972 33312 88024 33318
rect 87972 33254 88024 33260
rect 87696 31884 87748 31890
rect 87696 31826 87748 31832
rect 87708 31278 87736 31826
rect 87420 31272 87472 31278
rect 87420 31214 87472 31220
rect 87696 31272 87748 31278
rect 87696 31214 87748 31220
rect 85396 31204 85448 31210
rect 85396 31146 85448 31152
rect 86684 31204 86736 31210
rect 86684 31146 86736 31152
rect 84660 30932 84712 30938
rect 84660 30874 84712 30880
rect 85120 30932 85172 30938
rect 85120 30874 85172 30880
rect 84200 30796 84252 30802
rect 84200 30738 84252 30744
rect 83924 30728 83976 30734
rect 83924 30670 83976 30676
rect 84672 30394 84700 30874
rect 84660 30388 84712 30394
rect 84660 30330 84712 30336
rect 84672 30190 84700 30330
rect 85132 30326 85160 30874
rect 85304 30592 85356 30598
rect 85304 30534 85356 30540
rect 85316 30394 85344 30534
rect 85304 30388 85356 30394
rect 85304 30330 85356 30336
rect 85120 30320 85172 30326
rect 85120 30262 85172 30268
rect 85408 30190 85436 31146
rect 86592 30796 86644 30802
rect 86592 30738 86644 30744
rect 86604 30258 86632 30738
rect 86592 30252 86644 30258
rect 86592 30194 86644 30200
rect 86696 30190 86724 31146
rect 87432 31142 87460 31214
rect 87420 31136 87472 31142
rect 87420 31078 87472 31084
rect 87984 30938 88012 33254
rect 88352 32978 88380 33866
rect 88444 33114 88472 34002
rect 88524 33856 88576 33862
rect 88524 33798 88576 33804
rect 88536 33522 88564 33798
rect 89824 33658 89852 34002
rect 96380 33756 96676 33776
rect 96436 33754 96460 33756
rect 96516 33754 96540 33756
rect 96596 33754 96620 33756
rect 96458 33702 96460 33754
rect 96522 33702 96534 33754
rect 96596 33702 96598 33754
rect 96436 33700 96460 33702
rect 96516 33700 96540 33702
rect 96596 33700 96620 33702
rect 96380 33680 96676 33700
rect 89812 33652 89864 33658
rect 89812 33594 89864 33600
rect 88524 33516 88576 33522
rect 88524 33458 88576 33464
rect 88432 33108 88484 33114
rect 88432 33050 88484 33056
rect 88340 32972 88392 32978
rect 88340 32914 88392 32920
rect 96380 32668 96676 32688
rect 96436 32666 96460 32668
rect 96516 32666 96540 32668
rect 96596 32666 96620 32668
rect 96458 32614 96460 32666
rect 96522 32614 96534 32666
rect 96596 32614 96598 32666
rect 96436 32612 96460 32614
rect 96516 32612 96540 32614
rect 96596 32612 96620 32614
rect 96380 32592 96676 32612
rect 88248 31884 88300 31890
rect 88248 31826 88300 31832
rect 88260 30938 88288 31826
rect 96380 31580 96676 31600
rect 96436 31578 96460 31580
rect 96516 31578 96540 31580
rect 96596 31578 96620 31580
rect 96458 31526 96460 31578
rect 96522 31526 96534 31578
rect 96596 31526 96598 31578
rect 96436 31524 96460 31526
rect 96516 31524 96540 31526
rect 96596 31524 96620 31526
rect 96380 31504 96676 31524
rect 88616 31204 88668 31210
rect 88616 31146 88668 31152
rect 87972 30932 88024 30938
rect 87972 30874 88024 30880
rect 88248 30932 88300 30938
rect 88248 30874 88300 30880
rect 88260 30190 88288 30874
rect 88628 30802 88656 31146
rect 88616 30796 88668 30802
rect 88616 30738 88668 30744
rect 96380 30492 96676 30512
rect 96436 30490 96460 30492
rect 96516 30490 96540 30492
rect 96596 30490 96620 30492
rect 96458 30438 96460 30490
rect 96522 30438 96534 30490
rect 96596 30438 96598 30490
rect 96436 30436 96460 30438
rect 96516 30436 96540 30438
rect 96596 30436 96620 30438
rect 96380 30416 96676 30436
rect 84660 30184 84712 30190
rect 84660 30126 84712 30132
rect 85396 30184 85448 30190
rect 85396 30126 85448 30132
rect 86684 30184 86736 30190
rect 86684 30126 86736 30132
rect 88248 30184 88300 30190
rect 88248 30126 88300 30132
rect 86960 30116 87012 30122
rect 86960 30058 87012 30064
rect 83924 29572 83976 29578
rect 83924 29514 83976 29520
rect 83830 26072 83886 26081
rect 83830 26007 83886 26016
rect 59912 20800 59964 20806
rect 59912 20742 59964 20748
rect 83646 17776 83702 17785
rect 83646 17711 83702 17720
rect 59636 17400 59688 17406
rect 59636 17342 59688 17348
rect 83660 16697 83688 17711
rect 83646 16688 83702 16697
rect 83646 16623 83702 16632
rect 83660 12889 83688 16623
rect 83646 12880 83702 12889
rect 83646 12815 83702 12824
rect 83936 4729 83964 29514
rect 86316 29504 86368 29510
rect 86316 29446 86368 29452
rect 86500 29504 86552 29510
rect 86500 29446 86552 29452
rect 86592 29504 86644 29510
rect 86592 29446 86644 29452
rect 86328 23905 86356 29446
rect 86512 25537 86540 29446
rect 86498 25528 86554 25537
rect 86498 25463 86554 25472
rect 86314 23896 86370 23905
rect 86314 23831 86370 23840
rect 86604 21797 86632 29446
rect 86682 24984 86738 24993
rect 86972 24970 87000 30058
rect 87052 30048 87104 30054
rect 87052 29990 87104 29996
rect 86738 24942 87000 24970
rect 86682 24919 86738 24928
rect 87064 22930 87092 29990
rect 87144 29572 87196 29578
rect 87144 29514 87196 29520
rect 86972 22902 87092 22930
rect 86682 22876 86738 22885
rect 86972 22862 87000 22902
rect 86738 22834 87000 22862
rect 86682 22811 86738 22820
rect 86590 21788 86646 21797
rect 86590 21723 86646 21732
rect 86682 20700 86738 20709
rect 87156 20686 87184 29514
rect 87236 29504 87288 29510
rect 87236 29446 87288 29452
rect 87420 29504 87472 29510
rect 87420 29446 87472 29452
rect 87604 29504 87656 29510
rect 87604 29446 87656 29452
rect 86738 20658 87184 20686
rect 86682 20635 86738 20644
rect 87248 19650 87276 29446
rect 86684 19644 86736 19650
rect 86682 19612 86684 19621
rect 87236 19644 87288 19650
rect 86736 19612 86738 19621
rect 87236 19586 87288 19592
rect 86682 19547 86738 19556
rect 86684 17808 86736 17814
rect 86682 17776 86684 17785
rect 86736 17776 86738 17785
rect 86682 17711 86738 17720
rect 87432 17474 87460 29446
rect 87616 17814 87644 29446
rect 96380 29404 96676 29424
rect 96436 29402 96460 29404
rect 96516 29402 96540 29404
rect 96596 29402 96620 29404
rect 96458 29350 96460 29402
rect 96522 29350 96534 29402
rect 96596 29350 96598 29402
rect 96436 29348 96460 29350
rect 96516 29348 96540 29350
rect 96596 29348 96620 29350
rect 96380 29328 96676 29348
rect 87604 17808 87656 17814
rect 87604 17750 87656 17756
rect 86684 17468 86736 17474
rect 86682 17436 86684 17445
rect 87420 17468 87472 17474
rect 86736 17436 86738 17445
rect 87420 17410 87472 17416
rect 86682 17371 86738 17380
rect 59542 4720 59598 4729
rect 59542 4655 59598 4664
rect 83922 4720 83978 4729
rect 83922 4655 83978 4664
rect 53852 870 54616 898
rect 54588 800 54616 870
rect 3424 740 3476 746
rect 3424 682 3476 688
rect 8208 740 8260 746
rect 8208 682 8260 688
rect 3436 377 3464 682
rect 3422 368 3478 377
rect 3422 303 3478 312
rect 54574 0 54630 800
<< via2 >>
rect 3974 49680 4030 49736
rect 2778 49000 2834 49056
rect 4066 48356 4068 48376
rect 4068 48356 4120 48376
rect 4120 48356 4122 48376
rect 4066 48320 4122 48356
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 2870 39888 2926 39944
rect 2962 37304 3018 37360
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4066 45056 4122 45112
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 3974 43832 4030 43888
rect 3422 38528 3478 38584
rect 3054 29008 3110 29064
rect 2870 28192 2926 28248
rect 2778 24928 2834 24984
rect 2962 24248 3018 24304
rect 2870 22344 2926 22400
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4066 43152 4122 43208
rect 3974 42472 4030 42528
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4066 41792 4122 41848
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4066 41268 4122 41304
rect 4066 41248 4068 41268
rect 4068 41248 4120 41268
rect 4120 41248 4122 41268
rect 3790 39208 3846 39264
rect 3882 36624 3938 36680
rect 3698 34040 3754 34096
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4066 37984 4122 38040
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4066 35944 4122 36000
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4066 35400 4122 35456
rect 3974 34720 4030 34776
rect 3514 30776 3570 30832
rect 3330 27512 3386 27568
rect 3422 26832 3478 26888
rect 3238 26288 3294 26344
rect 3146 21664 3202 21720
rect 3330 19080 3386 19136
rect 3330 12008 3386 12064
rect 3790 32680 3846 32736
rect 3882 30096 3938 30152
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4066 33360 4122 33416
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4066 32136 4122 32192
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4066 31456 4122 31512
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4066 29552 4122 29608
rect 3974 28872 4030 28928
rect 3514 17176 3570 17232
rect 3882 25608 3938 25664
rect 3790 23024 3846 23080
rect 3698 18400 3754 18456
rect 3606 15816 3662 15872
rect 3514 9324 3516 9344
rect 3516 9324 3568 9344
rect 3568 9324 3570 9344
rect 3514 9288 3570 9324
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4066 23704 4122 23760
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4066 20984 4122 21040
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 3974 20476 3976 20496
rect 3976 20476 4028 20496
rect 4028 20476 4030 20496
rect 3974 20440 4030 20476
rect 3882 19760 3938 19816
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4066 17856 4122 17912
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4066 16496 4122 16552
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4066 15136 4122 15192
rect 3974 14592 4030 14648
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4066 13912 4122 13968
rect 3882 13232 3938 13288
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 3974 12552 4030 12608
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 3974 11328 4030 11384
rect 3974 10648 4030 10704
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3974 9968 4030 10024
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4066 8744 4122 8800
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 3790 8064 3846 8120
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 3974 7384 4030 7440
rect 3974 6740 3976 6760
rect 3976 6740 4028 6760
rect 4028 6740 4030 6760
rect 3974 6704 4030 6740
rect 3422 5480 3478 5536
rect 2962 4120 3018 4176
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4066 6160 4122 6216
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4066 4800 4122 4856
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4066 3440 4122 3496
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 5170 26188 5172 26208
rect 5172 26188 5224 26208
rect 5224 26188 5226 26208
rect 5170 26152 5226 26188
rect 6366 29008 6422 29064
rect 7838 40568 7894 40624
rect 9034 44376 9090 44432
rect 11150 41692 11152 41712
rect 11152 41692 11204 41712
rect 11204 41692 11206 41712
rect 11150 41656 11206 41692
rect 3330 2896 3386 2952
rect 2870 2252 2872 2272
rect 2872 2252 2924 2272
rect 2924 2252 2926 2272
rect 2870 2216 2926 2252
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 8298 26188 8300 26208
rect 8300 26188 8352 26208
rect 8352 26188 8354 26208
rect 8298 26152 8354 26188
rect 3238 1536 3294 1592
rect 2778 856 2834 912
rect 12530 37868 12586 37904
rect 12530 37848 12532 37868
rect 12532 37848 12584 37868
rect 12584 37848 12586 37868
rect 12898 33532 12900 33552
rect 12900 33532 12952 33552
rect 12952 33532 12954 33552
rect 12898 33496 12954 33532
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 50300 47354 50356 47356
rect 50380 47354 50436 47356
rect 50460 47354 50516 47356
rect 50540 47354 50596 47356
rect 50300 47302 50326 47354
rect 50326 47302 50356 47354
rect 50380 47302 50390 47354
rect 50390 47302 50436 47354
rect 50460 47302 50506 47354
rect 50506 47302 50516 47354
rect 50540 47302 50570 47354
rect 50570 47302 50596 47354
rect 50300 47300 50356 47302
rect 50380 47300 50436 47302
rect 50460 47300 50516 47302
rect 50540 47300 50596 47302
rect 12714 23468 12716 23488
rect 12716 23468 12768 23488
rect 12768 23468 12770 23488
rect 12714 23432 12770 23468
rect 13634 27532 13690 27568
rect 13634 27512 13636 27532
rect 13636 27512 13688 27532
rect 13688 27512 13690 27532
rect 14094 21256 14150 21312
rect 15290 27512 15346 27568
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 18694 41656 18750 41712
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 21822 40876 21824 40896
rect 21824 40876 21876 40896
rect 21876 40876 21878 40896
rect 21822 40840 21878 40876
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 20350 40704 20406 40760
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 14554 22752 14610 22808
rect 14186 17076 14188 17096
rect 14188 17076 14240 17096
rect 14240 17076 14242 17096
rect 14186 17040 14242 17076
rect 13450 16652 13506 16688
rect 13450 16632 13452 16652
rect 13452 16632 13504 16652
rect 13504 16632 13506 16652
rect 14830 23432 14886 23488
rect 15566 20032 15622 20088
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 18418 26152 18474 26208
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 22650 37884 22652 37904
rect 22652 37884 22704 37904
rect 22704 37884 22706 37904
rect 22650 37848 22706 37884
rect 21914 33924 21970 33960
rect 21914 33904 21916 33924
rect 21916 33904 21968 33924
rect 21968 33904 21970 33924
rect 22742 33496 22798 33552
rect 21730 32292 21786 32328
rect 21730 32272 21732 32292
rect 21732 32272 21784 32292
rect 21784 32272 21786 32292
rect 20258 29416 20314 29472
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 18786 23468 18788 23488
rect 18788 23468 18840 23488
rect 18840 23468 18842 23488
rect 18786 23432 18842 23468
rect 18970 20712 19026 20768
rect 19154 19352 19210 19408
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 22742 31340 22798 31376
rect 22742 31320 22744 31340
rect 22744 31320 22796 31340
rect 22796 31320 22798 31340
rect 22742 31204 22798 31240
rect 22742 31184 22744 31204
rect 22744 31184 22796 31204
rect 22796 31184 22798 31204
rect 23018 29300 23074 29336
rect 23018 29280 23020 29300
rect 23020 29280 23072 29300
rect 23072 29280 23074 29300
rect 20810 16632 20866 16688
rect 24214 29144 24270 29200
rect 21270 15972 21326 16008
rect 21270 15952 21272 15972
rect 21272 15952 21324 15972
rect 21324 15952 21326 15972
rect 28998 42220 29054 42256
rect 28998 42200 29000 42220
rect 29000 42200 29052 42220
rect 29052 42200 29054 42220
rect 26514 40704 26570 40760
rect 25134 29044 25136 29064
rect 25136 29044 25188 29064
rect 25188 29044 25190 29064
rect 25134 29008 25190 29044
rect 27434 40840 27490 40896
rect 27710 40296 27766 40352
rect 29090 40568 29146 40624
rect 29182 40332 29184 40352
rect 29184 40332 29236 40352
rect 29236 40332 29238 40352
rect 29182 40296 29238 40332
rect 25686 34484 25688 34504
rect 25688 34484 25740 34504
rect 25740 34484 25742 34504
rect 25686 34448 25742 34484
rect 26790 34448 26846 34504
rect 27066 34076 27068 34096
rect 27068 34076 27120 34096
rect 27120 34076 27122 34096
rect 27066 34040 27122 34076
rect 27526 34448 27582 34504
rect 27618 34076 27620 34096
rect 27620 34076 27672 34096
rect 27672 34076 27674 34096
rect 27618 34040 27674 34076
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 32770 43308 32826 43344
rect 32770 43288 32772 43308
rect 32772 43288 32824 43308
rect 32824 43288 32826 43308
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 32126 42236 32128 42256
rect 32128 42236 32180 42256
rect 32180 42236 32182 42256
rect 32126 42200 32182 42236
rect 30746 41540 30802 41576
rect 30746 41520 30748 41540
rect 30748 41520 30800 41540
rect 30800 41520 30802 41540
rect 35070 41556 35072 41576
rect 35072 41556 35124 41576
rect 35124 41556 35126 41576
rect 35070 41520 35126 41556
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34150 40604 34152 40624
rect 34152 40604 34204 40624
rect 34204 40604 34206 40624
rect 34150 40568 34206 40604
rect 27802 33924 27858 33960
rect 27802 33904 27804 33924
rect 27804 33904 27856 33924
rect 27856 33904 27858 33924
rect 27158 32308 27160 32328
rect 27160 32308 27212 32328
rect 27212 32308 27214 32328
rect 27158 32272 27214 32308
rect 25410 31340 25466 31376
rect 25410 31320 25412 31340
rect 25412 31320 25464 31340
rect 25464 31320 25466 31340
rect 25410 31204 25466 31240
rect 25410 31184 25412 31204
rect 25412 31184 25464 31204
rect 25464 31184 25466 31204
rect 25594 29280 25650 29336
rect 25410 29044 25412 29064
rect 25412 29044 25464 29064
rect 25464 29044 25466 29064
rect 25410 29008 25466 29044
rect 25410 21392 25466 21448
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 26422 29144 26478 29200
rect 26882 24012 26884 24032
rect 26884 24012 26936 24032
rect 26936 24012 26938 24032
rect 26882 23976 26938 24012
rect 31942 35692 31998 35728
rect 31942 35672 31944 35692
rect 31944 35672 31996 35692
rect 31996 35672 31998 35692
rect 32034 35572 32036 35592
rect 32036 35572 32088 35592
rect 32088 35572 32090 35592
rect 32034 35536 32090 35572
rect 31666 34992 31722 35048
rect 30654 33380 30710 33416
rect 30654 33360 30656 33380
rect 30656 33360 30708 33380
rect 30708 33360 30710 33380
rect 28170 29416 28226 29472
rect 31574 26042 31630 26098
rect 31666 25498 31722 25554
rect 31758 24998 31814 25054
rect 31574 23910 31630 23966
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 32586 35572 32588 35592
rect 32588 35572 32640 35592
rect 32640 35572 32642 35592
rect 32586 35536 32642 35572
rect 33782 35672 33838 35728
rect 33506 35536 33562 35592
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 37830 43308 37886 43344
rect 37830 43288 37832 43308
rect 37832 43288 37884 43308
rect 37884 43288 37886 43308
rect 38658 40840 38714 40896
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 35438 33396 35440 33416
rect 35440 33396 35492 33416
rect 35492 33396 35494 33416
rect 35438 33360 35494 33396
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 37462 34992 37518 35048
rect 39394 40588 39450 40624
rect 39394 40568 39396 40588
rect 39396 40568 39448 40588
rect 39448 40568 39450 40588
rect 40222 40604 40224 40624
rect 40224 40604 40276 40624
rect 40276 40604 40278 40624
rect 40222 40568 40278 40604
rect 40958 40840 41014 40896
rect 40590 40452 40646 40488
rect 40590 40432 40592 40452
rect 40592 40432 40644 40452
rect 40644 40432 40646 40452
rect 41602 40568 41658 40624
rect 40314 39616 40370 39672
rect 50300 46266 50356 46268
rect 50380 46266 50436 46268
rect 50460 46266 50516 46268
rect 50540 46266 50596 46268
rect 50300 46214 50326 46266
rect 50326 46214 50356 46266
rect 50380 46214 50390 46266
rect 50390 46214 50436 46266
rect 50460 46214 50506 46266
rect 50506 46214 50516 46266
rect 50540 46214 50570 46266
rect 50570 46214 50596 46266
rect 50300 46212 50356 46214
rect 50380 46212 50436 46214
rect 50460 46212 50516 46214
rect 50540 46212 50596 46214
rect 50300 45178 50356 45180
rect 50380 45178 50436 45180
rect 50460 45178 50516 45180
rect 50540 45178 50596 45180
rect 50300 45126 50326 45178
rect 50326 45126 50356 45178
rect 50380 45126 50390 45178
rect 50390 45126 50436 45178
rect 50460 45126 50506 45178
rect 50506 45126 50516 45178
rect 50540 45126 50570 45178
rect 50570 45126 50596 45178
rect 50300 45124 50356 45126
rect 50380 45124 50436 45126
rect 50460 45124 50516 45126
rect 50540 45124 50596 45126
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 44638 40452 44694 40488
rect 44638 40432 44640 40452
rect 44640 40432 44692 40452
rect 44692 40432 44694 40452
rect 42154 38972 42156 38992
rect 42156 38972 42208 38992
rect 42208 38972 42210 38992
rect 42154 38936 42210 38972
rect 39210 34584 39266 34640
rect 44546 37440 44602 37496
rect 44822 37440 44878 37496
rect 38750 33632 38806 33688
rect 38658 33516 38714 33552
rect 38658 33496 38660 33516
rect 38660 33496 38712 33516
rect 38712 33496 38714 33516
rect 38658 33360 38714 33416
rect 39486 33632 39542 33688
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 43534 34584 43590 34640
rect 43718 33496 43774 33552
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 41694 30640 41750 30696
rect 47582 39616 47638 39672
rect 47306 39344 47362 39400
rect 46662 37440 46718 37496
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 49054 39344 49110 39400
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 51170 38936 51226 38992
rect 50986 37340 50988 37360
rect 50988 37340 51040 37360
rect 51040 37340 51042 37360
rect 50986 37304 51042 37340
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 45282 29724 45284 29744
rect 45284 29724 45336 29744
rect 45336 29724 45338 29744
rect 45282 29688 45338 29724
rect 47030 29708 47086 29744
rect 47030 29688 47032 29708
rect 47032 29688 47084 29708
rect 47084 29688 47086 29708
rect 44178 29588 44180 29608
rect 44180 29588 44232 29608
rect 44232 29588 44234 29608
rect 44178 29552 44234 29588
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 65660 47898 65716 47900
rect 65740 47898 65796 47900
rect 65820 47898 65876 47900
rect 65900 47898 65956 47900
rect 65660 47846 65686 47898
rect 65686 47846 65716 47898
rect 65740 47846 65750 47898
rect 65750 47846 65796 47898
rect 65820 47846 65866 47898
rect 65866 47846 65876 47898
rect 65900 47846 65930 47898
rect 65930 47846 65956 47898
rect 65660 47844 65716 47846
rect 65740 47844 65796 47846
rect 65820 47844 65876 47846
rect 65900 47844 65956 47846
rect 54206 39924 54208 39944
rect 54208 39924 54260 39944
rect 54260 39924 54262 39944
rect 54206 39888 54262 39924
rect 50300 33210 50356 33212
rect 50380 33210 50436 33212
rect 50460 33210 50516 33212
rect 50540 33210 50596 33212
rect 50300 33158 50326 33210
rect 50326 33158 50356 33210
rect 50380 33158 50390 33210
rect 50390 33158 50436 33210
rect 50460 33158 50506 33210
rect 50506 33158 50516 33210
rect 50540 33158 50570 33210
rect 50570 33158 50596 33210
rect 50300 33156 50356 33158
rect 50380 33156 50436 33158
rect 50460 33156 50516 33158
rect 50540 33156 50596 33158
rect 51814 33380 51870 33416
rect 51814 33360 51816 33380
rect 51816 33360 51868 33380
rect 51868 33360 51870 33380
rect 48134 30640 48190 30696
rect 50300 32122 50356 32124
rect 50380 32122 50436 32124
rect 50460 32122 50516 32124
rect 50540 32122 50596 32124
rect 50300 32070 50326 32122
rect 50326 32070 50356 32122
rect 50380 32070 50390 32122
rect 50390 32070 50436 32122
rect 50460 32070 50506 32122
rect 50506 32070 50516 32122
rect 50540 32070 50570 32122
rect 50570 32070 50596 32122
rect 50300 32068 50356 32070
rect 50380 32068 50436 32070
rect 50460 32068 50516 32070
rect 50540 32068 50596 32070
rect 50300 31034 50356 31036
rect 50380 31034 50436 31036
rect 50460 31034 50516 31036
rect 50540 31034 50596 31036
rect 50300 30982 50326 31034
rect 50326 30982 50356 31034
rect 50380 30982 50390 31034
rect 50390 30982 50436 31034
rect 50460 30982 50506 31034
rect 50506 30982 50516 31034
rect 50540 30982 50570 31034
rect 50570 30982 50596 31034
rect 50300 30980 50356 30982
rect 50380 30980 50436 30982
rect 50460 30980 50516 30982
rect 50540 30980 50596 30982
rect 48962 29552 49018 29608
rect 48870 29452 48872 29472
rect 48872 29452 48924 29472
rect 48924 29452 48926 29472
rect 48870 29416 48926 29452
rect 50300 29946 50356 29948
rect 50380 29946 50436 29948
rect 50460 29946 50516 29948
rect 50540 29946 50596 29948
rect 50300 29894 50326 29946
rect 50326 29894 50356 29946
rect 50380 29894 50390 29946
rect 50390 29894 50436 29946
rect 50460 29894 50506 29946
rect 50506 29894 50516 29946
rect 50540 29894 50570 29946
rect 50570 29894 50596 29946
rect 50300 29892 50356 29894
rect 50380 29892 50436 29894
rect 50460 29892 50516 29894
rect 50540 29892 50596 29894
rect 54850 39888 54906 39944
rect 53194 29416 53250 29472
rect 31574 22778 31630 22834
rect 28998 21664 29054 21720
rect 28998 20576 29054 20632
rect 28906 19488 28962 19544
rect 28906 17312 28962 17368
rect 31758 13030 31814 13086
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 29918 4800 29974 4856
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 55310 37304 55366 37360
rect 55218 35164 55220 35184
rect 55220 35164 55272 35184
rect 55272 35164 55274 35184
rect 55218 35128 55274 35164
rect 56598 35284 56654 35320
rect 56598 35264 56600 35284
rect 56600 35264 56652 35284
rect 56652 35264 56654 35284
rect 56966 35264 57022 35320
rect 58714 43308 58770 43344
rect 58714 43288 58716 43308
rect 58716 43288 58768 43308
rect 58768 43288 58770 43308
rect 59174 41148 59176 41168
rect 59176 41148 59228 41168
rect 59228 41148 59230 41168
rect 59174 41112 59230 41148
rect 60830 39072 60886 39128
rect 60738 38936 60794 38992
rect 65660 46810 65716 46812
rect 65740 46810 65796 46812
rect 65820 46810 65876 46812
rect 65900 46810 65956 46812
rect 65660 46758 65686 46810
rect 65686 46758 65716 46810
rect 65740 46758 65750 46810
rect 65750 46758 65796 46810
rect 65820 46758 65866 46810
rect 65866 46758 65876 46810
rect 65900 46758 65930 46810
rect 65930 46758 65956 46810
rect 65660 46756 65716 46758
rect 65740 46756 65796 46758
rect 65820 46756 65876 46758
rect 65900 46756 65956 46758
rect 65660 45722 65716 45724
rect 65740 45722 65796 45724
rect 65820 45722 65876 45724
rect 65900 45722 65956 45724
rect 65660 45670 65686 45722
rect 65686 45670 65716 45722
rect 65740 45670 65750 45722
rect 65750 45670 65796 45722
rect 65820 45670 65866 45722
rect 65866 45670 65876 45722
rect 65900 45670 65930 45722
rect 65930 45670 65956 45722
rect 65660 45668 65716 45670
rect 65740 45668 65796 45670
rect 65820 45668 65876 45670
rect 65900 45668 65956 45670
rect 65660 44634 65716 44636
rect 65740 44634 65796 44636
rect 65820 44634 65876 44636
rect 65900 44634 65956 44636
rect 65660 44582 65686 44634
rect 65686 44582 65716 44634
rect 65740 44582 65750 44634
rect 65750 44582 65796 44634
rect 65820 44582 65866 44634
rect 65866 44582 65876 44634
rect 65900 44582 65930 44634
rect 65930 44582 65956 44634
rect 65660 44580 65716 44582
rect 65740 44580 65796 44582
rect 65820 44580 65876 44582
rect 65900 44580 65956 44582
rect 65660 43546 65716 43548
rect 65740 43546 65796 43548
rect 65820 43546 65876 43548
rect 65900 43546 65956 43548
rect 65660 43494 65686 43546
rect 65686 43494 65716 43546
rect 65740 43494 65750 43546
rect 65750 43494 65796 43546
rect 65820 43494 65866 43546
rect 65866 43494 65876 43546
rect 65900 43494 65930 43546
rect 65930 43494 65956 43546
rect 65660 43492 65716 43494
rect 65740 43492 65796 43494
rect 65820 43492 65876 43494
rect 65900 43492 65956 43494
rect 65660 42458 65716 42460
rect 65740 42458 65796 42460
rect 65820 42458 65876 42460
rect 65900 42458 65956 42460
rect 65660 42406 65686 42458
rect 65686 42406 65716 42458
rect 65740 42406 65750 42458
rect 65750 42406 65796 42458
rect 65820 42406 65866 42458
rect 65866 42406 65876 42458
rect 65900 42406 65930 42458
rect 65930 42406 65956 42458
rect 65660 42404 65716 42406
rect 65740 42404 65796 42406
rect 65820 42404 65876 42406
rect 65900 42404 65956 42406
rect 65660 41370 65716 41372
rect 65740 41370 65796 41372
rect 65820 41370 65876 41372
rect 65900 41370 65956 41372
rect 65660 41318 65686 41370
rect 65686 41318 65716 41370
rect 65740 41318 65750 41370
rect 65750 41318 65796 41370
rect 65820 41318 65866 41370
rect 65866 41318 65876 41370
rect 65900 41318 65930 41370
rect 65930 41318 65956 41370
rect 65660 41316 65716 41318
rect 65740 41316 65796 41318
rect 65820 41316 65876 41318
rect 65900 41316 65956 41318
rect 56598 26188 56600 26208
rect 56600 26188 56652 26208
rect 56652 26188 56654 26208
rect 56598 26152 56654 26188
rect 56690 25608 56746 25664
rect 59174 29008 59230 29064
rect 59082 25004 59138 25060
rect 58990 22828 59046 22884
rect 57794 21800 57850 21856
rect 59358 25548 59414 25604
rect 59358 23860 59414 23916
rect 59358 21392 59414 21448
rect 59266 20652 59322 20708
rect 59358 19564 59414 19620
rect 59358 17348 59360 17394
rect 59360 17348 59412 17394
rect 59412 17348 59414 17394
rect 59358 17338 59414 17348
rect 60646 29996 60648 30016
rect 60648 29996 60700 30016
rect 60700 29996 60702 30016
rect 60646 29960 60702 29996
rect 63590 39072 63646 39128
rect 61566 32972 61622 33008
rect 61566 32952 61568 32972
rect 61568 32952 61620 32972
rect 61620 32952 61622 32972
rect 61934 29960 61990 30016
rect 65660 40282 65716 40284
rect 65740 40282 65796 40284
rect 65820 40282 65876 40284
rect 65900 40282 65956 40284
rect 65660 40230 65686 40282
rect 65686 40230 65716 40282
rect 65740 40230 65750 40282
rect 65750 40230 65796 40282
rect 65820 40230 65866 40282
rect 65866 40230 65876 40282
rect 65900 40230 65930 40282
rect 65930 40230 65956 40282
rect 65660 40228 65716 40230
rect 65740 40228 65796 40230
rect 65820 40228 65876 40230
rect 65900 40228 65956 40230
rect 67086 43288 67142 43344
rect 67362 41112 67418 41168
rect 71594 41112 71650 41168
rect 71778 40976 71834 41032
rect 65660 39194 65716 39196
rect 65740 39194 65796 39196
rect 65820 39194 65876 39196
rect 65900 39194 65956 39196
rect 65660 39142 65686 39194
rect 65686 39142 65716 39194
rect 65740 39142 65750 39194
rect 65750 39142 65796 39194
rect 65820 39142 65866 39194
rect 65866 39142 65876 39194
rect 65900 39142 65930 39194
rect 65930 39142 65956 39194
rect 65660 39140 65716 39142
rect 65740 39140 65796 39142
rect 65820 39140 65876 39142
rect 65900 39140 65956 39142
rect 66902 38936 66958 38992
rect 65660 38106 65716 38108
rect 65740 38106 65796 38108
rect 65820 38106 65876 38108
rect 65900 38106 65956 38108
rect 65660 38054 65686 38106
rect 65686 38054 65716 38106
rect 65740 38054 65750 38106
rect 65750 38054 65796 38106
rect 65820 38054 65866 38106
rect 65866 38054 65876 38106
rect 65900 38054 65930 38106
rect 65930 38054 65956 38106
rect 65660 38052 65716 38054
rect 65740 38052 65796 38054
rect 65820 38052 65876 38054
rect 65900 38052 65956 38054
rect 65660 37018 65716 37020
rect 65740 37018 65796 37020
rect 65820 37018 65876 37020
rect 65900 37018 65956 37020
rect 65660 36966 65686 37018
rect 65686 36966 65716 37018
rect 65740 36966 65750 37018
rect 65750 36966 65796 37018
rect 65820 36966 65866 37018
rect 65866 36966 65876 37018
rect 65900 36966 65930 37018
rect 65930 36966 65956 37018
rect 65660 36964 65716 36966
rect 65740 36964 65796 36966
rect 65820 36964 65876 36966
rect 65900 36964 65956 36966
rect 65660 35930 65716 35932
rect 65740 35930 65796 35932
rect 65820 35930 65876 35932
rect 65900 35930 65956 35932
rect 65660 35878 65686 35930
rect 65686 35878 65716 35930
rect 65740 35878 65750 35930
rect 65750 35878 65796 35930
rect 65820 35878 65866 35930
rect 65866 35878 65876 35930
rect 65900 35878 65930 35930
rect 65930 35878 65956 35930
rect 65660 35876 65716 35878
rect 65740 35876 65796 35878
rect 65820 35876 65876 35878
rect 65900 35876 65956 35878
rect 64694 35128 64750 35184
rect 65660 34842 65716 34844
rect 65740 34842 65796 34844
rect 65820 34842 65876 34844
rect 65900 34842 65956 34844
rect 65660 34790 65686 34842
rect 65686 34790 65716 34842
rect 65740 34790 65750 34842
rect 65750 34790 65796 34842
rect 65820 34790 65866 34842
rect 65866 34790 65876 34842
rect 65900 34790 65930 34842
rect 65930 34790 65956 34842
rect 65660 34788 65716 34790
rect 65740 34788 65796 34790
rect 65820 34788 65876 34790
rect 65900 34788 65956 34790
rect 65660 33754 65716 33756
rect 65740 33754 65796 33756
rect 65820 33754 65876 33756
rect 65900 33754 65956 33756
rect 65660 33702 65686 33754
rect 65686 33702 65716 33754
rect 65740 33702 65750 33754
rect 65750 33702 65796 33754
rect 65820 33702 65866 33754
rect 65866 33702 65876 33754
rect 65900 33702 65930 33754
rect 65930 33702 65956 33754
rect 65660 33700 65716 33702
rect 65740 33700 65796 33702
rect 65820 33700 65876 33702
rect 65900 33700 65956 33702
rect 66994 32988 66996 33008
rect 66996 32988 67048 33008
rect 67048 32988 67050 33008
rect 66994 32952 67050 32988
rect 65660 32666 65716 32668
rect 65740 32666 65796 32668
rect 65820 32666 65876 32668
rect 65900 32666 65956 32668
rect 65660 32614 65686 32666
rect 65686 32614 65716 32666
rect 65740 32614 65750 32666
rect 65750 32614 65796 32666
rect 65820 32614 65866 32666
rect 65866 32614 65876 32666
rect 65900 32614 65930 32666
rect 65930 32614 65956 32666
rect 65660 32612 65716 32614
rect 65740 32612 65796 32614
rect 65820 32612 65876 32614
rect 65900 32612 65956 32614
rect 65660 31578 65716 31580
rect 65740 31578 65796 31580
rect 65820 31578 65876 31580
rect 65900 31578 65956 31580
rect 65660 31526 65686 31578
rect 65686 31526 65716 31578
rect 65740 31526 65750 31578
rect 65750 31526 65796 31578
rect 65820 31526 65866 31578
rect 65866 31526 65876 31578
rect 65900 31526 65930 31578
rect 65930 31526 65956 31578
rect 65660 31524 65716 31526
rect 65740 31524 65796 31526
rect 65820 31524 65876 31526
rect 65900 31524 65956 31526
rect 65660 30490 65716 30492
rect 65740 30490 65796 30492
rect 65820 30490 65876 30492
rect 65900 30490 65956 30492
rect 65660 30438 65686 30490
rect 65686 30438 65716 30490
rect 65740 30438 65750 30490
rect 65750 30438 65796 30490
rect 65820 30438 65866 30490
rect 65866 30438 65876 30490
rect 65900 30438 65930 30490
rect 65930 30438 65956 30490
rect 65660 30436 65716 30438
rect 65740 30436 65796 30438
rect 65820 30436 65876 30438
rect 65900 30436 65956 30438
rect 65660 29402 65716 29404
rect 65740 29402 65796 29404
rect 65820 29402 65876 29404
rect 65900 29402 65956 29404
rect 65660 29350 65686 29402
rect 65686 29350 65716 29402
rect 65740 29350 65750 29402
rect 65750 29350 65796 29402
rect 65820 29350 65866 29402
rect 65866 29350 65876 29402
rect 65900 29350 65930 29402
rect 65930 29350 65956 29402
rect 65660 29348 65716 29350
rect 65740 29348 65796 29350
rect 65820 29348 65876 29350
rect 65900 29348 65956 29350
rect 68650 35536 68706 35592
rect 72514 41112 72570 41168
rect 72330 41012 72332 41032
rect 72332 41012 72384 41032
rect 72384 41012 72386 41032
rect 72330 40976 72386 41012
rect 81020 47354 81076 47356
rect 81100 47354 81156 47356
rect 81180 47354 81236 47356
rect 81260 47354 81316 47356
rect 81020 47302 81046 47354
rect 81046 47302 81076 47354
rect 81100 47302 81110 47354
rect 81110 47302 81156 47354
rect 81180 47302 81226 47354
rect 81226 47302 81236 47354
rect 81260 47302 81290 47354
rect 81290 47302 81316 47354
rect 81020 47300 81076 47302
rect 81100 47300 81156 47302
rect 81180 47300 81236 47302
rect 81260 47300 81316 47302
rect 96380 47898 96436 47900
rect 96460 47898 96516 47900
rect 96540 47898 96596 47900
rect 96620 47898 96676 47900
rect 96380 47846 96406 47898
rect 96406 47846 96436 47898
rect 96460 47846 96470 47898
rect 96470 47846 96516 47898
rect 96540 47846 96586 47898
rect 96586 47846 96596 47898
rect 96620 47846 96650 47898
rect 96650 47846 96676 47898
rect 96380 47844 96436 47846
rect 96460 47844 96516 47846
rect 96540 47844 96596 47846
rect 96620 47844 96676 47846
rect 96380 46810 96436 46812
rect 96460 46810 96516 46812
rect 96540 46810 96596 46812
rect 96620 46810 96676 46812
rect 96380 46758 96406 46810
rect 96406 46758 96436 46810
rect 96460 46758 96470 46810
rect 96470 46758 96516 46810
rect 96540 46758 96586 46810
rect 96586 46758 96596 46810
rect 96620 46758 96650 46810
rect 96650 46758 96676 46810
rect 96380 46756 96436 46758
rect 96460 46756 96516 46758
rect 96540 46756 96596 46758
rect 96620 46756 96676 46758
rect 81020 46266 81076 46268
rect 81100 46266 81156 46268
rect 81180 46266 81236 46268
rect 81260 46266 81316 46268
rect 81020 46214 81046 46266
rect 81046 46214 81076 46266
rect 81100 46214 81110 46266
rect 81110 46214 81156 46266
rect 81180 46214 81226 46266
rect 81226 46214 81236 46266
rect 81260 46214 81290 46266
rect 81290 46214 81316 46266
rect 81020 46212 81076 46214
rect 81100 46212 81156 46214
rect 81180 46212 81236 46214
rect 81260 46212 81316 46214
rect 81020 45178 81076 45180
rect 81100 45178 81156 45180
rect 81180 45178 81236 45180
rect 81260 45178 81316 45180
rect 81020 45126 81046 45178
rect 81046 45126 81076 45178
rect 81100 45126 81110 45178
rect 81110 45126 81156 45178
rect 81180 45126 81226 45178
rect 81226 45126 81236 45178
rect 81260 45126 81290 45178
rect 81290 45126 81316 45178
rect 81020 45124 81076 45126
rect 81100 45124 81156 45126
rect 81180 45124 81236 45126
rect 81260 45124 81316 45126
rect 81020 44090 81076 44092
rect 81100 44090 81156 44092
rect 81180 44090 81236 44092
rect 81260 44090 81316 44092
rect 81020 44038 81046 44090
rect 81046 44038 81076 44090
rect 81100 44038 81110 44090
rect 81110 44038 81156 44090
rect 81180 44038 81226 44090
rect 81226 44038 81236 44090
rect 81260 44038 81290 44090
rect 81290 44038 81316 44090
rect 81020 44036 81076 44038
rect 81100 44036 81156 44038
rect 81180 44036 81236 44038
rect 81260 44036 81316 44038
rect 70122 34348 70124 34368
rect 70124 34348 70176 34368
rect 70176 34348 70178 34368
rect 70122 34312 70178 34348
rect 74170 35556 74226 35592
rect 74170 35536 74172 35556
rect 74172 35536 74224 35556
rect 74224 35536 74226 35556
rect 81020 43002 81076 43004
rect 81100 43002 81156 43004
rect 81180 43002 81236 43004
rect 81260 43002 81316 43004
rect 81020 42950 81046 43002
rect 81046 42950 81076 43002
rect 81100 42950 81110 43002
rect 81110 42950 81156 43002
rect 81180 42950 81226 43002
rect 81226 42950 81236 43002
rect 81260 42950 81290 43002
rect 81290 42950 81316 43002
rect 81020 42948 81076 42950
rect 81100 42948 81156 42950
rect 81180 42948 81236 42950
rect 81260 42948 81316 42950
rect 81020 41914 81076 41916
rect 81100 41914 81156 41916
rect 81180 41914 81236 41916
rect 81260 41914 81316 41916
rect 81020 41862 81046 41914
rect 81046 41862 81076 41914
rect 81100 41862 81110 41914
rect 81110 41862 81156 41914
rect 81180 41862 81226 41914
rect 81226 41862 81236 41914
rect 81260 41862 81290 41914
rect 81290 41862 81316 41914
rect 81020 41860 81076 41862
rect 81100 41860 81156 41862
rect 81180 41860 81236 41862
rect 81260 41860 81316 41862
rect 81020 40826 81076 40828
rect 81100 40826 81156 40828
rect 81180 40826 81236 40828
rect 81260 40826 81316 40828
rect 81020 40774 81046 40826
rect 81046 40774 81076 40826
rect 81100 40774 81110 40826
rect 81110 40774 81156 40826
rect 81180 40774 81226 40826
rect 81226 40774 81236 40826
rect 81260 40774 81290 40826
rect 81290 40774 81316 40826
rect 81020 40772 81076 40774
rect 81100 40772 81156 40774
rect 81180 40772 81236 40774
rect 81260 40772 81316 40774
rect 81020 39738 81076 39740
rect 81100 39738 81156 39740
rect 81180 39738 81236 39740
rect 81260 39738 81316 39740
rect 81020 39686 81046 39738
rect 81046 39686 81076 39738
rect 81100 39686 81110 39738
rect 81110 39686 81156 39738
rect 81180 39686 81226 39738
rect 81226 39686 81236 39738
rect 81260 39686 81290 39738
rect 81290 39686 81316 39738
rect 81020 39684 81076 39686
rect 81100 39684 81156 39686
rect 81180 39684 81236 39686
rect 81260 39684 81316 39686
rect 81020 38650 81076 38652
rect 81100 38650 81156 38652
rect 81180 38650 81236 38652
rect 81260 38650 81316 38652
rect 81020 38598 81046 38650
rect 81046 38598 81076 38650
rect 81100 38598 81110 38650
rect 81110 38598 81156 38650
rect 81180 38598 81226 38650
rect 81226 38598 81236 38650
rect 81260 38598 81290 38650
rect 81290 38598 81316 38650
rect 81020 38596 81076 38598
rect 81100 38596 81156 38598
rect 81180 38596 81236 38598
rect 81260 38596 81316 38598
rect 81020 37562 81076 37564
rect 81100 37562 81156 37564
rect 81180 37562 81236 37564
rect 81260 37562 81316 37564
rect 81020 37510 81046 37562
rect 81046 37510 81076 37562
rect 81100 37510 81110 37562
rect 81110 37510 81156 37562
rect 81180 37510 81226 37562
rect 81226 37510 81236 37562
rect 81260 37510 81290 37562
rect 81290 37510 81316 37562
rect 81020 37508 81076 37510
rect 81100 37508 81156 37510
rect 81180 37508 81236 37510
rect 81260 37508 81316 37510
rect 81020 36474 81076 36476
rect 81100 36474 81156 36476
rect 81180 36474 81236 36476
rect 81260 36474 81316 36476
rect 81020 36422 81046 36474
rect 81046 36422 81076 36474
rect 81100 36422 81110 36474
rect 81110 36422 81156 36474
rect 81180 36422 81226 36474
rect 81226 36422 81236 36474
rect 81260 36422 81290 36474
rect 81290 36422 81316 36474
rect 81020 36420 81076 36422
rect 81100 36420 81156 36422
rect 81180 36420 81236 36422
rect 81260 36420 81316 36422
rect 76286 34348 76288 34368
rect 76288 34348 76340 34368
rect 76340 34348 76342 34368
rect 76286 34312 76342 34348
rect 81020 35386 81076 35388
rect 81100 35386 81156 35388
rect 81180 35386 81236 35388
rect 81260 35386 81316 35388
rect 81020 35334 81046 35386
rect 81046 35334 81076 35386
rect 81100 35334 81110 35386
rect 81110 35334 81156 35386
rect 81180 35334 81226 35386
rect 81226 35334 81236 35386
rect 81260 35334 81290 35386
rect 81290 35334 81316 35386
rect 81020 35332 81076 35334
rect 81100 35332 81156 35334
rect 81180 35332 81236 35334
rect 81260 35332 81316 35334
rect 81020 34298 81076 34300
rect 81100 34298 81156 34300
rect 81180 34298 81236 34300
rect 81260 34298 81316 34300
rect 81020 34246 81046 34298
rect 81046 34246 81076 34298
rect 81100 34246 81110 34298
rect 81110 34246 81156 34298
rect 81180 34246 81226 34298
rect 81226 34246 81236 34298
rect 81260 34246 81290 34298
rect 81290 34246 81316 34298
rect 81020 34244 81076 34246
rect 81100 34244 81156 34246
rect 81180 34244 81236 34246
rect 81260 34244 81316 34246
rect 81020 33210 81076 33212
rect 81100 33210 81156 33212
rect 81180 33210 81236 33212
rect 81260 33210 81316 33212
rect 81020 33158 81046 33210
rect 81046 33158 81076 33210
rect 81100 33158 81110 33210
rect 81110 33158 81156 33210
rect 81180 33158 81226 33210
rect 81226 33158 81236 33210
rect 81260 33158 81290 33210
rect 81290 33158 81316 33210
rect 81020 33156 81076 33158
rect 81100 33156 81156 33158
rect 81180 33156 81236 33158
rect 81260 33156 81316 33158
rect 81020 32122 81076 32124
rect 81100 32122 81156 32124
rect 81180 32122 81236 32124
rect 81260 32122 81316 32124
rect 81020 32070 81046 32122
rect 81046 32070 81076 32122
rect 81100 32070 81110 32122
rect 81110 32070 81156 32122
rect 81180 32070 81226 32122
rect 81226 32070 81236 32122
rect 81260 32070 81290 32122
rect 81290 32070 81316 32122
rect 81020 32068 81076 32070
rect 81100 32068 81156 32070
rect 81180 32068 81236 32070
rect 81260 32068 81316 32070
rect 81020 31034 81076 31036
rect 81100 31034 81156 31036
rect 81180 31034 81236 31036
rect 81260 31034 81316 31036
rect 81020 30982 81046 31034
rect 81046 30982 81076 31034
rect 81100 30982 81110 31034
rect 81110 30982 81156 31034
rect 81180 30982 81226 31034
rect 81226 30982 81236 31034
rect 81260 30982 81290 31034
rect 81290 30982 81316 31034
rect 81020 30980 81076 30982
rect 81100 30980 81156 30982
rect 81180 30980 81236 30982
rect 81260 30980 81316 30982
rect 81020 29946 81076 29948
rect 81100 29946 81156 29948
rect 81180 29946 81236 29948
rect 81260 29946 81316 29948
rect 81020 29894 81046 29946
rect 81046 29894 81076 29946
rect 81100 29894 81110 29946
rect 81110 29894 81156 29946
rect 81180 29894 81226 29946
rect 81226 29894 81236 29946
rect 81260 29894 81290 29946
rect 81290 29894 81316 29946
rect 81020 29892 81076 29894
rect 81100 29892 81156 29894
rect 81180 29892 81236 29894
rect 81260 29892 81316 29894
rect 96380 45722 96436 45724
rect 96460 45722 96516 45724
rect 96540 45722 96596 45724
rect 96620 45722 96676 45724
rect 96380 45670 96406 45722
rect 96406 45670 96436 45722
rect 96460 45670 96470 45722
rect 96470 45670 96516 45722
rect 96540 45670 96586 45722
rect 96586 45670 96596 45722
rect 96620 45670 96650 45722
rect 96650 45670 96676 45722
rect 96380 45668 96436 45670
rect 96460 45668 96516 45670
rect 96540 45668 96596 45670
rect 96620 45668 96676 45670
rect 96380 44634 96436 44636
rect 96460 44634 96516 44636
rect 96540 44634 96596 44636
rect 96620 44634 96676 44636
rect 96380 44582 96406 44634
rect 96406 44582 96436 44634
rect 96460 44582 96470 44634
rect 96470 44582 96516 44634
rect 96540 44582 96586 44634
rect 96586 44582 96596 44634
rect 96620 44582 96650 44634
rect 96650 44582 96676 44634
rect 96380 44580 96436 44582
rect 96460 44580 96516 44582
rect 96540 44580 96596 44582
rect 96620 44580 96676 44582
rect 96380 43546 96436 43548
rect 96460 43546 96516 43548
rect 96540 43546 96596 43548
rect 96620 43546 96676 43548
rect 96380 43494 96406 43546
rect 96406 43494 96436 43546
rect 96460 43494 96470 43546
rect 96470 43494 96516 43546
rect 96540 43494 96586 43546
rect 96586 43494 96596 43546
rect 96620 43494 96650 43546
rect 96650 43494 96676 43546
rect 96380 43492 96436 43494
rect 96460 43492 96516 43494
rect 96540 43492 96596 43494
rect 96620 43492 96676 43494
rect 96380 42458 96436 42460
rect 96460 42458 96516 42460
rect 96540 42458 96596 42460
rect 96620 42458 96676 42460
rect 96380 42406 96406 42458
rect 96406 42406 96436 42458
rect 96460 42406 96470 42458
rect 96470 42406 96516 42458
rect 96540 42406 96586 42458
rect 96586 42406 96596 42458
rect 96620 42406 96650 42458
rect 96650 42406 96676 42458
rect 96380 42404 96436 42406
rect 96460 42404 96516 42406
rect 96540 42404 96596 42406
rect 96620 42404 96676 42406
rect 96380 41370 96436 41372
rect 96460 41370 96516 41372
rect 96540 41370 96596 41372
rect 96620 41370 96676 41372
rect 96380 41318 96406 41370
rect 96406 41318 96436 41370
rect 96460 41318 96470 41370
rect 96470 41318 96516 41370
rect 96540 41318 96586 41370
rect 96586 41318 96596 41370
rect 96620 41318 96650 41370
rect 96650 41318 96676 41370
rect 96380 41316 96436 41318
rect 96460 41316 96516 41318
rect 96540 41316 96596 41318
rect 96620 41316 96676 41318
rect 96380 40282 96436 40284
rect 96460 40282 96516 40284
rect 96540 40282 96596 40284
rect 96620 40282 96676 40284
rect 96380 40230 96406 40282
rect 96406 40230 96436 40282
rect 96460 40230 96470 40282
rect 96470 40230 96516 40282
rect 96540 40230 96586 40282
rect 96586 40230 96596 40282
rect 96620 40230 96650 40282
rect 96650 40230 96676 40282
rect 96380 40228 96436 40230
rect 96460 40228 96516 40230
rect 96540 40228 96596 40230
rect 96620 40228 96676 40230
rect 96380 39194 96436 39196
rect 96460 39194 96516 39196
rect 96540 39194 96596 39196
rect 96620 39194 96676 39196
rect 96380 39142 96406 39194
rect 96406 39142 96436 39194
rect 96460 39142 96470 39194
rect 96470 39142 96516 39194
rect 96540 39142 96586 39194
rect 96586 39142 96596 39194
rect 96620 39142 96650 39194
rect 96650 39142 96676 39194
rect 96380 39140 96436 39142
rect 96460 39140 96516 39142
rect 96540 39140 96596 39142
rect 96620 39140 96676 39142
rect 96380 38106 96436 38108
rect 96460 38106 96516 38108
rect 96540 38106 96596 38108
rect 96620 38106 96676 38108
rect 96380 38054 96406 38106
rect 96406 38054 96436 38106
rect 96460 38054 96470 38106
rect 96470 38054 96516 38106
rect 96540 38054 96586 38106
rect 96586 38054 96596 38106
rect 96620 38054 96650 38106
rect 96650 38054 96676 38106
rect 96380 38052 96436 38054
rect 96460 38052 96516 38054
rect 96540 38052 96596 38054
rect 96620 38052 96676 38054
rect 96380 37018 96436 37020
rect 96460 37018 96516 37020
rect 96540 37018 96596 37020
rect 96620 37018 96676 37020
rect 96380 36966 96406 37018
rect 96406 36966 96436 37018
rect 96460 36966 96470 37018
rect 96470 36966 96516 37018
rect 96540 36966 96586 37018
rect 96586 36966 96596 37018
rect 96620 36966 96650 37018
rect 96650 36966 96676 37018
rect 96380 36964 96436 36966
rect 96460 36964 96516 36966
rect 96540 36964 96596 36966
rect 96620 36964 96676 36966
rect 96380 35930 96436 35932
rect 96460 35930 96516 35932
rect 96540 35930 96596 35932
rect 96620 35930 96676 35932
rect 96380 35878 96406 35930
rect 96406 35878 96436 35930
rect 96460 35878 96470 35930
rect 96470 35878 96516 35930
rect 96540 35878 96586 35930
rect 96586 35878 96596 35930
rect 96620 35878 96650 35930
rect 96650 35878 96676 35930
rect 96380 35876 96436 35878
rect 96460 35876 96516 35878
rect 96540 35876 96596 35878
rect 96620 35876 96676 35878
rect 96380 34842 96436 34844
rect 96460 34842 96516 34844
rect 96540 34842 96596 34844
rect 96620 34842 96676 34844
rect 96380 34790 96406 34842
rect 96406 34790 96436 34842
rect 96460 34790 96470 34842
rect 96470 34790 96516 34842
rect 96540 34790 96586 34842
rect 96586 34790 96596 34842
rect 96620 34790 96650 34842
rect 96650 34790 96676 34842
rect 96380 34788 96436 34790
rect 96460 34788 96516 34790
rect 96540 34788 96596 34790
rect 96620 34788 96676 34790
rect 96380 33754 96436 33756
rect 96460 33754 96516 33756
rect 96540 33754 96596 33756
rect 96620 33754 96676 33756
rect 96380 33702 96406 33754
rect 96406 33702 96436 33754
rect 96460 33702 96470 33754
rect 96470 33702 96516 33754
rect 96540 33702 96586 33754
rect 96586 33702 96596 33754
rect 96620 33702 96650 33754
rect 96650 33702 96676 33754
rect 96380 33700 96436 33702
rect 96460 33700 96516 33702
rect 96540 33700 96596 33702
rect 96620 33700 96676 33702
rect 96380 32666 96436 32668
rect 96460 32666 96516 32668
rect 96540 32666 96596 32668
rect 96620 32666 96676 32668
rect 96380 32614 96406 32666
rect 96406 32614 96436 32666
rect 96460 32614 96470 32666
rect 96470 32614 96516 32666
rect 96540 32614 96586 32666
rect 96586 32614 96596 32666
rect 96620 32614 96650 32666
rect 96650 32614 96676 32666
rect 96380 32612 96436 32614
rect 96460 32612 96516 32614
rect 96540 32612 96596 32614
rect 96620 32612 96676 32614
rect 96380 31578 96436 31580
rect 96460 31578 96516 31580
rect 96540 31578 96596 31580
rect 96620 31578 96676 31580
rect 96380 31526 96406 31578
rect 96406 31526 96436 31578
rect 96460 31526 96470 31578
rect 96470 31526 96516 31578
rect 96540 31526 96586 31578
rect 96586 31526 96596 31578
rect 96620 31526 96650 31578
rect 96650 31526 96676 31578
rect 96380 31524 96436 31526
rect 96460 31524 96516 31526
rect 96540 31524 96596 31526
rect 96620 31524 96676 31526
rect 96380 30490 96436 30492
rect 96460 30490 96516 30492
rect 96540 30490 96596 30492
rect 96620 30490 96676 30492
rect 96380 30438 96406 30490
rect 96406 30438 96436 30490
rect 96460 30438 96470 30490
rect 96470 30438 96516 30490
rect 96540 30438 96586 30490
rect 96586 30438 96596 30490
rect 96620 30438 96650 30490
rect 96650 30438 96676 30490
rect 96380 30436 96436 30438
rect 96460 30436 96516 30438
rect 96540 30436 96596 30438
rect 96620 30436 96676 30438
rect 83830 26016 83886 26072
rect 83646 17720 83702 17776
rect 83646 16632 83702 16688
rect 83646 12824 83702 12880
rect 86498 25472 86554 25528
rect 86314 23840 86370 23896
rect 86682 24928 86738 24984
rect 86682 22820 86738 22876
rect 86590 21732 86646 21788
rect 86682 20644 86738 20700
rect 86682 19592 86684 19612
rect 86684 19592 86736 19612
rect 86736 19592 86738 19612
rect 86682 19556 86738 19592
rect 86682 17756 86684 17776
rect 86684 17756 86736 17776
rect 86736 17756 86738 17776
rect 86682 17720 86738 17756
rect 96380 29402 96436 29404
rect 96460 29402 96516 29404
rect 96540 29402 96596 29404
rect 96620 29402 96676 29404
rect 96380 29350 96406 29402
rect 96406 29350 96436 29402
rect 96460 29350 96470 29402
rect 96470 29350 96516 29402
rect 96540 29350 96586 29402
rect 96586 29350 96596 29402
rect 96620 29350 96650 29402
rect 96650 29350 96676 29402
rect 96380 29348 96436 29350
rect 96460 29348 96516 29350
rect 96540 29348 96596 29350
rect 96620 29348 96676 29350
rect 86682 17416 86684 17436
rect 86684 17416 86736 17436
rect 86736 17416 86738 17436
rect 86682 17380 86738 17416
rect 59542 4664 59598 4720
rect 83922 4664 83978 4720
rect 3422 312 3478 368
<< metal3 >>
rect 0 49738 800 49768
rect 3969 49738 4035 49741
rect 0 49736 4035 49738
rect 0 49680 3974 49736
rect 4030 49680 4035 49736
rect 0 49678 4035 49680
rect 0 49648 800 49678
rect 3969 49675 4035 49678
rect 0 49058 800 49088
rect 2773 49058 2839 49061
rect 0 49056 2839 49058
rect 0 49000 2778 49056
rect 2834 49000 2839 49056
rect 0 48998 2839 49000
rect 0 48968 800 48998
rect 2773 48995 2839 48998
rect 0 48378 800 48408
rect 4061 48378 4127 48381
rect 0 48376 4127 48378
rect 0 48320 4066 48376
rect 4122 48320 4127 48376
rect 0 48318 4127 48320
rect 0 48288 800 48318
rect 4061 48315 4127 48318
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 65648 47904 65968 47905
rect 65648 47840 65656 47904
rect 65720 47840 65736 47904
rect 65800 47840 65816 47904
rect 65880 47840 65896 47904
rect 65960 47840 65968 47904
rect 65648 47839 65968 47840
rect 96368 47904 96688 47905
rect 96368 47840 96376 47904
rect 96440 47840 96456 47904
rect 96520 47840 96536 47904
rect 96600 47840 96616 47904
rect 96680 47840 96688 47904
rect 96368 47839 96688 47840
rect 0 47608 800 47728
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 50288 47360 50608 47361
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 47295 50608 47296
rect 81008 47360 81328 47361
rect 81008 47296 81016 47360
rect 81080 47296 81096 47360
rect 81160 47296 81176 47360
rect 81240 47296 81256 47360
rect 81320 47296 81328 47360
rect 81008 47295 81328 47296
rect 0 47064 800 47184
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 65648 46816 65968 46817
rect 65648 46752 65656 46816
rect 65720 46752 65736 46816
rect 65800 46752 65816 46816
rect 65880 46752 65896 46816
rect 65960 46752 65968 46816
rect 65648 46751 65968 46752
rect 96368 46816 96688 46817
rect 96368 46752 96376 46816
rect 96440 46752 96456 46816
rect 96520 46752 96536 46816
rect 96600 46752 96616 46816
rect 96680 46752 96688 46816
rect 96368 46751 96688 46752
rect 0 46384 800 46504
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 50288 46272 50608 46273
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 46207 50608 46208
rect 81008 46272 81328 46273
rect 81008 46208 81016 46272
rect 81080 46208 81096 46272
rect 81160 46208 81176 46272
rect 81240 46208 81256 46272
rect 81320 46208 81328 46272
rect 81008 46207 81328 46208
rect 0 45704 800 45824
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 65648 45728 65968 45729
rect 65648 45664 65656 45728
rect 65720 45664 65736 45728
rect 65800 45664 65816 45728
rect 65880 45664 65896 45728
rect 65960 45664 65968 45728
rect 65648 45663 65968 45664
rect 96368 45728 96688 45729
rect 96368 45664 96376 45728
rect 96440 45664 96456 45728
rect 96520 45664 96536 45728
rect 96600 45664 96616 45728
rect 96680 45664 96688 45728
rect 96368 45663 96688 45664
rect 19568 45184 19888 45185
rect 0 45114 800 45144
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 50288 45184 50608 45185
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 45119 50608 45120
rect 81008 45184 81328 45185
rect 81008 45120 81016 45184
rect 81080 45120 81096 45184
rect 81160 45120 81176 45184
rect 81240 45120 81256 45184
rect 81320 45120 81328 45184
rect 81008 45119 81328 45120
rect 4061 45114 4127 45117
rect 0 45112 4127 45114
rect 0 45056 4066 45112
rect 4122 45056 4127 45112
rect 0 45054 4127 45056
rect 0 45024 800 45054
rect 4061 45051 4127 45054
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 65648 44640 65968 44641
rect 65648 44576 65656 44640
rect 65720 44576 65736 44640
rect 65800 44576 65816 44640
rect 65880 44576 65896 44640
rect 65960 44576 65968 44640
rect 65648 44575 65968 44576
rect 96368 44640 96688 44641
rect 96368 44576 96376 44640
rect 96440 44576 96456 44640
rect 96520 44576 96536 44640
rect 96600 44576 96616 44640
rect 96680 44576 96688 44640
rect 96368 44575 96688 44576
rect 0 44434 800 44464
rect 9029 44434 9095 44437
rect 0 44432 9095 44434
rect 0 44376 9034 44432
rect 9090 44376 9095 44432
rect 0 44374 9095 44376
rect 0 44344 800 44374
rect 9029 44371 9095 44374
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 44031 50608 44032
rect 81008 44096 81328 44097
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 44031 81328 44032
rect 0 43890 800 43920
rect 3969 43890 4035 43893
rect 0 43888 4035 43890
rect 0 43832 3974 43888
rect 4030 43832 4035 43888
rect 0 43830 4035 43832
rect 0 43800 800 43830
rect 3969 43827 4035 43830
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 65648 43552 65968 43553
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43487 65968 43488
rect 96368 43552 96688 43553
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43487 96688 43488
rect 32765 43346 32831 43349
rect 37825 43346 37891 43349
rect 32765 43344 37891 43346
rect 32765 43288 32770 43344
rect 32826 43288 37830 43344
rect 37886 43288 37891 43344
rect 32765 43286 37891 43288
rect 32765 43283 32831 43286
rect 37825 43283 37891 43286
rect 58709 43346 58775 43349
rect 67081 43346 67147 43349
rect 58709 43344 67147 43346
rect 58709 43288 58714 43344
rect 58770 43288 67086 43344
rect 67142 43288 67147 43344
rect 58709 43286 67147 43288
rect 58709 43283 58775 43286
rect 67081 43283 67147 43286
rect 0 43210 800 43240
rect 4061 43210 4127 43213
rect 0 43208 4127 43210
rect 0 43152 4066 43208
rect 4122 43152 4127 43208
rect 0 43150 4127 43152
rect 0 43120 800 43150
rect 4061 43147 4127 43150
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 42943 50608 42944
rect 81008 43008 81328 43009
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 42943 81328 42944
rect 0 42530 800 42560
rect 3969 42530 4035 42533
rect 0 42528 4035 42530
rect 0 42472 3974 42528
rect 4030 42472 4035 42528
rect 0 42470 4035 42472
rect 0 42440 800 42470
rect 3969 42467 4035 42470
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 65648 42464 65968 42465
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 42399 65968 42400
rect 96368 42464 96688 42465
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 42399 96688 42400
rect 28993 42258 29059 42261
rect 32121 42258 32187 42261
rect 28993 42256 32187 42258
rect 28993 42200 28998 42256
rect 29054 42200 32126 42256
rect 32182 42200 32187 42256
rect 28993 42198 32187 42200
rect 28993 42195 29059 42198
rect 32121 42195 32187 42198
rect 19568 41920 19888 41921
rect 0 41850 800 41880
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 41855 50608 41856
rect 81008 41920 81328 41921
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 41855 81328 41856
rect 4061 41850 4127 41853
rect 0 41848 4127 41850
rect 0 41792 4066 41848
rect 4122 41792 4127 41848
rect 0 41790 4127 41792
rect 0 41760 800 41790
rect 4061 41787 4127 41790
rect 11145 41714 11211 41717
rect 18689 41714 18755 41717
rect 11145 41712 18755 41714
rect 11145 41656 11150 41712
rect 11206 41656 18694 41712
rect 18750 41656 18755 41712
rect 11145 41654 18755 41656
rect 11145 41651 11211 41654
rect 18689 41651 18755 41654
rect 30741 41578 30807 41581
rect 35065 41578 35131 41581
rect 30741 41576 35131 41578
rect 30741 41520 30746 41576
rect 30802 41520 35070 41576
rect 35126 41520 35131 41576
rect 30741 41518 35131 41520
rect 30741 41515 30807 41518
rect 35065 41515 35131 41518
rect 4208 41376 4528 41377
rect 0 41306 800 41336
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 65648 41376 65968 41377
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 41311 65968 41312
rect 96368 41376 96688 41377
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 41311 96688 41312
rect 4061 41306 4127 41309
rect 0 41304 4127 41306
rect 0 41248 4066 41304
rect 4122 41248 4127 41304
rect 0 41246 4127 41248
rect 0 41216 800 41246
rect 4061 41243 4127 41246
rect 59169 41170 59235 41173
rect 67357 41170 67423 41173
rect 59169 41168 67423 41170
rect 59169 41112 59174 41168
rect 59230 41112 67362 41168
rect 67418 41112 67423 41168
rect 59169 41110 67423 41112
rect 59169 41107 59235 41110
rect 67357 41107 67423 41110
rect 71589 41170 71655 41173
rect 72509 41170 72575 41173
rect 71589 41168 72575 41170
rect 71589 41112 71594 41168
rect 71650 41112 72514 41168
rect 72570 41112 72575 41168
rect 71589 41110 72575 41112
rect 71589 41107 71655 41110
rect 72509 41107 72575 41110
rect 71773 41034 71839 41037
rect 72325 41034 72391 41037
rect 71773 41032 72391 41034
rect 71773 40976 71778 41032
rect 71834 40976 72330 41032
rect 72386 40976 72391 41032
rect 71773 40974 72391 40976
rect 71773 40971 71839 40974
rect 72325 40971 72391 40974
rect 21817 40898 21883 40901
rect 27429 40898 27495 40901
rect 21817 40896 27495 40898
rect 21817 40840 21822 40896
rect 21878 40840 27434 40896
rect 27490 40840 27495 40896
rect 21817 40838 27495 40840
rect 21817 40835 21883 40838
rect 27429 40835 27495 40838
rect 38653 40898 38719 40901
rect 40953 40898 41019 40901
rect 38653 40896 41019 40898
rect 38653 40840 38658 40896
rect 38714 40840 40958 40896
rect 41014 40840 41019 40896
rect 38653 40838 41019 40840
rect 38653 40835 38719 40838
rect 40953 40835 41019 40838
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 40767 50608 40768
rect 81008 40832 81328 40833
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 40767 81328 40768
rect 20345 40762 20411 40765
rect 26509 40762 26575 40765
rect 20345 40760 26575 40762
rect 20345 40704 20350 40760
rect 20406 40704 26514 40760
rect 26570 40704 26575 40760
rect 20345 40702 26575 40704
rect 20345 40699 20411 40702
rect 26509 40699 26575 40702
rect 0 40626 800 40656
rect 7833 40626 7899 40629
rect 0 40624 7899 40626
rect 0 40568 7838 40624
rect 7894 40568 7899 40624
rect 0 40566 7899 40568
rect 0 40536 800 40566
rect 7833 40563 7899 40566
rect 29085 40626 29151 40629
rect 34145 40626 34211 40629
rect 29085 40624 34211 40626
rect 29085 40568 29090 40624
rect 29146 40568 34150 40624
rect 34206 40568 34211 40624
rect 29085 40566 34211 40568
rect 29085 40563 29151 40566
rect 34145 40563 34211 40566
rect 39389 40626 39455 40629
rect 40217 40626 40283 40629
rect 41597 40626 41663 40629
rect 39389 40624 41663 40626
rect 39389 40568 39394 40624
rect 39450 40568 40222 40624
rect 40278 40568 41602 40624
rect 41658 40568 41663 40624
rect 39389 40566 41663 40568
rect 39389 40563 39455 40566
rect 40217 40563 40283 40566
rect 41597 40563 41663 40566
rect 40585 40490 40651 40493
rect 44633 40490 44699 40493
rect 40585 40488 44699 40490
rect 40585 40432 40590 40488
rect 40646 40432 44638 40488
rect 44694 40432 44699 40488
rect 40585 40430 44699 40432
rect 40585 40427 40651 40430
rect 44633 40427 44699 40430
rect 27705 40354 27771 40357
rect 29177 40354 29243 40357
rect 27705 40352 29243 40354
rect 27705 40296 27710 40352
rect 27766 40296 29182 40352
rect 29238 40296 29243 40352
rect 27705 40294 29243 40296
rect 27705 40291 27771 40294
rect 29177 40291 29243 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 65648 40288 65968 40289
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 40223 65968 40224
rect 96368 40288 96688 40289
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 40223 96688 40224
rect 0 39946 800 39976
rect 2865 39946 2931 39949
rect 0 39944 2931 39946
rect 0 39888 2870 39944
rect 2926 39888 2931 39944
rect 0 39886 2931 39888
rect 0 39856 800 39886
rect 2865 39883 2931 39886
rect 54201 39946 54267 39949
rect 54845 39946 54911 39949
rect 54201 39944 54911 39946
rect 54201 39888 54206 39944
rect 54262 39888 54850 39944
rect 54906 39888 54911 39944
rect 54201 39886 54911 39888
rect 54201 39883 54267 39886
rect 54845 39883 54911 39886
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 39679 50608 39680
rect 81008 39744 81328 39745
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 39679 81328 39680
rect 40309 39674 40375 39677
rect 47577 39674 47643 39677
rect 40309 39672 47643 39674
rect 40309 39616 40314 39672
rect 40370 39616 47582 39672
rect 47638 39616 47643 39672
rect 40309 39614 47643 39616
rect 40309 39611 40375 39614
rect 47577 39611 47643 39614
rect 47301 39402 47367 39405
rect 49049 39402 49115 39405
rect 47301 39400 49115 39402
rect 47301 39344 47306 39400
rect 47362 39344 49054 39400
rect 49110 39344 49115 39400
rect 47301 39342 49115 39344
rect 47301 39339 47367 39342
rect 49049 39339 49115 39342
rect 0 39266 800 39296
rect 3785 39266 3851 39269
rect 0 39264 3851 39266
rect 0 39208 3790 39264
rect 3846 39208 3851 39264
rect 0 39206 3851 39208
rect 0 39176 800 39206
rect 3785 39203 3851 39206
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 65648 39200 65968 39201
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 39135 65968 39136
rect 96368 39200 96688 39201
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 39135 96688 39136
rect 60825 39130 60891 39133
rect 63585 39130 63651 39133
rect 60825 39128 63651 39130
rect 60825 39072 60830 39128
rect 60886 39072 63590 39128
rect 63646 39072 63651 39128
rect 60825 39070 63651 39072
rect 60825 39067 60891 39070
rect 63585 39067 63651 39070
rect 42149 38994 42215 38997
rect 51165 38994 51231 38997
rect 42149 38992 51231 38994
rect 42149 38936 42154 38992
rect 42210 38936 51170 38992
rect 51226 38936 51231 38992
rect 42149 38934 51231 38936
rect 42149 38931 42215 38934
rect 51165 38931 51231 38934
rect 60733 38994 60799 38997
rect 66897 38994 66963 38997
rect 60733 38992 66963 38994
rect 60733 38936 60738 38992
rect 60794 38936 66902 38992
rect 66958 38936 66963 38992
rect 60733 38934 66963 38936
rect 60733 38931 60799 38934
rect 66897 38931 66963 38934
rect 19568 38656 19888 38657
rect 0 38586 800 38616
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 38591 50608 38592
rect 81008 38656 81328 38657
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 38591 81328 38592
rect 3417 38586 3483 38589
rect 0 38584 3483 38586
rect 0 38528 3422 38584
rect 3478 38528 3483 38584
rect 0 38526 3483 38528
rect 0 38496 800 38526
rect 3417 38523 3483 38526
rect 4208 38112 4528 38113
rect 0 38042 800 38072
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 65648 38112 65968 38113
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 38047 65968 38048
rect 96368 38112 96688 38113
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 38047 96688 38048
rect 4061 38042 4127 38045
rect 0 38040 4127 38042
rect 0 37984 4066 38040
rect 4122 37984 4127 38040
rect 0 37982 4127 37984
rect 0 37952 800 37982
rect 4061 37979 4127 37982
rect 12525 37906 12591 37909
rect 22645 37906 22711 37909
rect 12525 37904 22711 37906
rect 12525 37848 12530 37904
rect 12586 37848 22650 37904
rect 22706 37848 22711 37904
rect 12525 37846 22711 37848
rect 12525 37843 12591 37846
rect 22645 37843 22711 37846
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 81008 37568 81328 37569
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 37503 81328 37504
rect 44541 37498 44607 37501
rect 44817 37498 44883 37501
rect 46657 37498 46723 37501
rect 44541 37496 46723 37498
rect 44541 37440 44546 37496
rect 44602 37440 44822 37496
rect 44878 37440 46662 37496
rect 46718 37440 46723 37496
rect 44541 37438 46723 37440
rect 44541 37435 44607 37438
rect 44817 37435 44883 37438
rect 46657 37435 46723 37438
rect 0 37362 800 37392
rect 2957 37362 3023 37365
rect 0 37360 3023 37362
rect 0 37304 2962 37360
rect 3018 37304 3023 37360
rect 0 37302 3023 37304
rect 0 37272 800 37302
rect 2957 37299 3023 37302
rect 50981 37362 51047 37365
rect 55305 37362 55371 37365
rect 50981 37360 55371 37362
rect 50981 37304 50986 37360
rect 51042 37304 55310 37360
rect 55366 37304 55371 37360
rect 50981 37302 55371 37304
rect 50981 37299 51047 37302
rect 55305 37299 55371 37302
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 65648 37024 65968 37025
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 36959 65968 36960
rect 96368 37024 96688 37025
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 36959 96688 36960
rect 0 36682 800 36712
rect 3877 36682 3943 36685
rect 0 36680 3943 36682
rect 0 36624 3882 36680
rect 3938 36624 3943 36680
rect 0 36622 3943 36624
rect 0 36592 800 36622
rect 3877 36619 3943 36622
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 81008 36480 81328 36481
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 36415 81328 36416
rect 0 36002 800 36032
rect 4061 36002 4127 36005
rect 0 36000 4127 36002
rect 0 35944 4066 36000
rect 4122 35944 4127 36000
rect 0 35942 4127 35944
rect 0 35912 800 35942
rect 4061 35939 4127 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 65648 35936 65968 35937
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 35871 65968 35872
rect 96368 35936 96688 35937
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 35871 96688 35872
rect 31937 35730 32003 35733
rect 33777 35730 33843 35733
rect 31937 35728 33843 35730
rect 31937 35672 31942 35728
rect 31998 35672 33782 35728
rect 33838 35672 33843 35728
rect 31937 35670 33843 35672
rect 31937 35667 32003 35670
rect 33777 35667 33843 35670
rect 32029 35594 32095 35597
rect 32581 35594 32647 35597
rect 33501 35594 33567 35597
rect 32029 35592 33567 35594
rect 32029 35536 32034 35592
rect 32090 35536 32586 35592
rect 32642 35536 33506 35592
rect 33562 35536 33567 35592
rect 32029 35534 33567 35536
rect 32029 35531 32095 35534
rect 32581 35531 32647 35534
rect 33501 35531 33567 35534
rect 68645 35594 68711 35597
rect 74165 35594 74231 35597
rect 68645 35592 74231 35594
rect 68645 35536 68650 35592
rect 68706 35536 74170 35592
rect 74226 35536 74231 35592
rect 68645 35534 74231 35536
rect 68645 35531 68711 35534
rect 74165 35531 74231 35534
rect 0 35458 800 35488
rect 4061 35458 4127 35461
rect 0 35456 4127 35458
rect 0 35400 4066 35456
rect 4122 35400 4127 35456
rect 0 35398 4127 35400
rect 0 35368 800 35398
rect 4061 35395 4127 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 81008 35392 81328 35393
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 35327 81328 35328
rect 56593 35322 56659 35325
rect 56961 35322 57027 35325
rect 56593 35320 57027 35322
rect 56593 35264 56598 35320
rect 56654 35264 56966 35320
rect 57022 35264 57027 35320
rect 56593 35262 57027 35264
rect 56593 35259 56659 35262
rect 56961 35259 57027 35262
rect 55213 35186 55279 35189
rect 64689 35186 64755 35189
rect 55213 35184 64755 35186
rect 55213 35128 55218 35184
rect 55274 35128 64694 35184
rect 64750 35128 64755 35184
rect 55213 35126 64755 35128
rect 55213 35123 55279 35126
rect 64689 35123 64755 35126
rect 31661 35050 31727 35053
rect 37457 35050 37523 35053
rect 31661 35048 37523 35050
rect 31661 34992 31666 35048
rect 31722 34992 37462 35048
rect 37518 34992 37523 35048
rect 31661 34990 37523 34992
rect 31661 34987 31727 34990
rect 37457 34987 37523 34990
rect 4208 34848 4528 34849
rect 0 34778 800 34808
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 65648 34848 65968 34849
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 34783 65968 34784
rect 96368 34848 96688 34849
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 34783 96688 34784
rect 3969 34778 4035 34781
rect 0 34776 4035 34778
rect 0 34720 3974 34776
rect 4030 34720 4035 34776
rect 0 34718 4035 34720
rect 0 34688 800 34718
rect 3969 34715 4035 34718
rect 39205 34642 39271 34645
rect 43529 34642 43595 34645
rect 39205 34640 43595 34642
rect 39205 34584 39210 34640
rect 39266 34584 43534 34640
rect 43590 34584 43595 34640
rect 39205 34582 43595 34584
rect 39205 34579 39271 34582
rect 43529 34579 43595 34582
rect 25681 34506 25747 34509
rect 26785 34506 26851 34509
rect 27521 34506 27587 34509
rect 25681 34504 27587 34506
rect 25681 34448 25686 34504
rect 25742 34448 26790 34504
rect 26846 34448 27526 34504
rect 27582 34448 27587 34504
rect 25681 34446 27587 34448
rect 25681 34443 25747 34446
rect 26785 34443 26851 34446
rect 27521 34443 27587 34446
rect 70117 34370 70183 34373
rect 76281 34370 76347 34373
rect 70117 34368 76347 34370
rect 70117 34312 70122 34368
rect 70178 34312 76286 34368
rect 76342 34312 76347 34368
rect 70117 34310 76347 34312
rect 70117 34307 70183 34310
rect 76281 34307 76347 34310
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 81008 34304 81328 34305
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 34239 81328 34240
rect 0 34098 800 34128
rect 3693 34098 3759 34101
rect 0 34096 3759 34098
rect 0 34040 3698 34096
rect 3754 34040 3759 34096
rect 0 34038 3759 34040
rect 0 34008 800 34038
rect 3693 34035 3759 34038
rect 27061 34098 27127 34101
rect 27613 34098 27679 34101
rect 27061 34096 27679 34098
rect 27061 34040 27066 34096
rect 27122 34040 27618 34096
rect 27674 34040 27679 34096
rect 27061 34038 27679 34040
rect 27061 34035 27127 34038
rect 27613 34035 27679 34038
rect 21909 33962 21975 33965
rect 27797 33962 27863 33965
rect 21909 33960 27863 33962
rect 21909 33904 21914 33960
rect 21970 33904 27802 33960
rect 27858 33904 27863 33960
rect 21909 33902 27863 33904
rect 21909 33899 21975 33902
rect 27797 33899 27863 33902
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 65648 33760 65968 33761
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 33695 65968 33696
rect 96368 33760 96688 33761
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 33695 96688 33696
rect 38745 33690 38811 33693
rect 39481 33690 39547 33693
rect 38745 33688 39547 33690
rect 38745 33632 38750 33688
rect 38806 33632 39486 33688
rect 39542 33632 39547 33688
rect 38745 33630 39547 33632
rect 38745 33627 38811 33630
rect 39481 33627 39547 33630
rect 12893 33554 12959 33557
rect 22737 33554 22803 33557
rect 12893 33552 22803 33554
rect 12893 33496 12898 33552
rect 12954 33496 22742 33552
rect 22798 33496 22803 33552
rect 12893 33494 22803 33496
rect 12893 33491 12959 33494
rect 22737 33491 22803 33494
rect 38653 33554 38719 33557
rect 43713 33554 43779 33557
rect 38653 33552 43779 33554
rect 38653 33496 38658 33552
rect 38714 33496 43718 33552
rect 43774 33496 43779 33552
rect 38653 33494 43779 33496
rect 38653 33491 38719 33494
rect 43713 33491 43779 33494
rect 0 33418 800 33448
rect 4061 33418 4127 33421
rect 0 33416 4127 33418
rect 0 33360 4066 33416
rect 4122 33360 4127 33416
rect 0 33358 4127 33360
rect 0 33328 800 33358
rect 4061 33355 4127 33358
rect 30649 33418 30715 33421
rect 35433 33418 35499 33421
rect 30649 33416 35499 33418
rect 30649 33360 30654 33416
rect 30710 33360 35438 33416
rect 35494 33360 35499 33416
rect 30649 33358 35499 33360
rect 30649 33355 30715 33358
rect 35433 33355 35499 33358
rect 38653 33418 38719 33421
rect 51809 33418 51875 33421
rect 38653 33416 51875 33418
rect 38653 33360 38658 33416
rect 38714 33360 51814 33416
rect 51870 33360 51875 33416
rect 38653 33358 51875 33360
rect 38653 33355 38719 33358
rect 51809 33355 51875 33358
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 50288 33216 50608 33217
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 33151 50608 33152
rect 81008 33216 81328 33217
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 33151 81328 33152
rect 61561 33010 61627 33013
rect 66989 33010 67055 33013
rect 61561 33008 67055 33010
rect 61561 32952 61566 33008
rect 61622 32952 66994 33008
rect 67050 32952 67055 33008
rect 61561 32950 67055 32952
rect 61561 32947 61627 32950
rect 66989 32947 67055 32950
rect 0 32738 800 32768
rect 3785 32738 3851 32741
rect 0 32736 3851 32738
rect 0 32680 3790 32736
rect 3846 32680 3851 32736
rect 0 32678 3851 32680
rect 0 32648 800 32678
rect 3785 32675 3851 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 65648 32672 65968 32673
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 32607 65968 32608
rect 96368 32672 96688 32673
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 32607 96688 32608
rect 21725 32330 21791 32333
rect 27153 32330 27219 32333
rect 21725 32328 27219 32330
rect 21725 32272 21730 32328
rect 21786 32272 27158 32328
rect 27214 32272 27219 32328
rect 21725 32270 27219 32272
rect 21725 32267 21791 32270
rect 27153 32267 27219 32270
rect 0 32194 800 32224
rect 4061 32194 4127 32197
rect 0 32192 4127 32194
rect 0 32136 4066 32192
rect 4122 32136 4127 32192
rect 0 32134 4127 32136
rect 0 32104 800 32134
rect 4061 32131 4127 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 50288 32128 50608 32129
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 32063 50608 32064
rect 81008 32128 81328 32129
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 32063 81328 32064
rect 4208 31584 4528 31585
rect 0 31514 800 31544
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 65648 31584 65968 31585
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 31519 65968 31520
rect 96368 31584 96688 31585
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 31519 96688 31520
rect 4061 31514 4127 31517
rect 0 31512 4127 31514
rect 0 31456 4066 31512
rect 4122 31456 4127 31512
rect 0 31454 4127 31456
rect 0 31424 800 31454
rect 4061 31451 4127 31454
rect 22737 31378 22803 31381
rect 25405 31378 25471 31381
rect 22737 31376 25471 31378
rect 22737 31320 22742 31376
rect 22798 31320 25410 31376
rect 25466 31320 25471 31376
rect 22737 31318 25471 31320
rect 22737 31315 22803 31318
rect 25405 31315 25471 31318
rect 22737 31242 22803 31245
rect 25405 31242 25471 31245
rect 22737 31240 25471 31242
rect 22737 31184 22742 31240
rect 22798 31184 25410 31240
rect 25466 31184 25471 31240
rect 22737 31182 25471 31184
rect 22737 31179 22803 31182
rect 25405 31179 25471 31182
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 50288 31040 50608 31041
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 30975 50608 30976
rect 81008 31040 81328 31041
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 30975 81328 30976
rect 0 30834 800 30864
rect 3509 30834 3575 30837
rect 0 30832 3575 30834
rect 0 30776 3514 30832
rect 3570 30776 3575 30832
rect 0 30774 3575 30776
rect 0 30744 800 30774
rect 3509 30771 3575 30774
rect 41689 30698 41755 30701
rect 48129 30698 48195 30701
rect 41689 30696 48195 30698
rect 41689 30640 41694 30696
rect 41750 30640 48134 30696
rect 48190 30640 48195 30696
rect 41689 30638 48195 30640
rect 41689 30635 41755 30638
rect 48129 30635 48195 30638
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 65648 30496 65968 30497
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 30431 65968 30432
rect 96368 30496 96688 30497
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 30431 96688 30432
rect 0 30154 800 30184
rect 3877 30154 3943 30157
rect 0 30152 3943 30154
rect 0 30096 3882 30152
rect 3938 30096 3943 30152
rect 0 30094 3943 30096
rect 0 30064 800 30094
rect 3877 30091 3943 30094
rect 60641 30018 60707 30021
rect 61929 30018 61995 30021
rect 60641 30016 61995 30018
rect 60641 29960 60646 30016
rect 60702 29960 61934 30016
rect 61990 29960 61995 30016
rect 60641 29958 61995 29960
rect 60641 29955 60707 29958
rect 61929 29955 61995 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 50288 29952 50608 29953
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29887 50608 29888
rect 81008 29952 81328 29953
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 29887 81328 29888
rect 45277 29746 45343 29749
rect 47025 29746 47091 29749
rect 45277 29744 47091 29746
rect 45277 29688 45282 29744
rect 45338 29688 47030 29744
rect 47086 29688 47091 29744
rect 45277 29686 47091 29688
rect 45277 29683 45343 29686
rect 47025 29683 47091 29686
rect 0 29610 800 29640
rect 4061 29610 4127 29613
rect 0 29608 4127 29610
rect 0 29552 4066 29608
rect 4122 29552 4127 29608
rect 0 29550 4127 29552
rect 0 29520 800 29550
rect 4061 29547 4127 29550
rect 44173 29610 44239 29613
rect 48957 29610 49023 29613
rect 44173 29608 49023 29610
rect 44173 29552 44178 29608
rect 44234 29552 48962 29608
rect 49018 29552 49023 29608
rect 44173 29550 49023 29552
rect 44173 29547 44239 29550
rect 48957 29547 49023 29550
rect 20253 29474 20319 29477
rect 28165 29474 28231 29477
rect 20253 29472 28231 29474
rect 20253 29416 20258 29472
rect 20314 29416 28170 29472
rect 28226 29416 28231 29472
rect 20253 29414 28231 29416
rect 20253 29411 20319 29414
rect 28165 29411 28231 29414
rect 48865 29474 48931 29477
rect 53189 29474 53255 29477
rect 48865 29472 53255 29474
rect 48865 29416 48870 29472
rect 48926 29416 53194 29472
rect 53250 29416 53255 29472
rect 48865 29414 53255 29416
rect 48865 29411 48931 29414
rect 53189 29411 53255 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 65648 29408 65968 29409
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 29343 65968 29344
rect 96368 29408 96688 29409
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 29343 96688 29344
rect 23013 29338 23079 29341
rect 25589 29338 25655 29341
rect 23013 29336 25655 29338
rect 23013 29280 23018 29336
rect 23074 29280 25594 29336
rect 25650 29280 25655 29336
rect 23013 29278 25655 29280
rect 23013 29275 23079 29278
rect 25589 29275 25655 29278
rect 24209 29202 24275 29205
rect 26417 29202 26483 29205
rect 24209 29200 26483 29202
rect 24209 29144 24214 29200
rect 24270 29144 26422 29200
rect 26478 29144 26483 29200
rect 24209 29142 26483 29144
rect 24209 29139 24275 29142
rect 26417 29139 26483 29142
rect 3049 29066 3115 29069
rect 6361 29066 6427 29069
rect 3049 29064 6427 29066
rect 3049 29008 3054 29064
rect 3110 29008 6366 29064
rect 6422 29008 6427 29064
rect 3049 29006 6427 29008
rect 3049 29003 3115 29006
rect 6361 29003 6427 29006
rect 25129 29066 25195 29069
rect 25405 29066 25471 29069
rect 59169 29068 59235 29069
rect 59118 29066 59124 29068
rect 25129 29064 25471 29066
rect 25129 29008 25134 29064
rect 25190 29008 25410 29064
rect 25466 29008 25471 29064
rect 25129 29006 25471 29008
rect 59078 29006 59124 29066
rect 59188 29064 59235 29068
rect 59230 29008 59235 29064
rect 25129 29003 25195 29006
rect 25405 29003 25471 29006
rect 59118 29004 59124 29006
rect 59188 29004 59235 29008
rect 59169 29003 59235 29004
rect 0 28930 800 28960
rect 3969 28930 4035 28933
rect 0 28928 4035 28930
rect 0 28872 3974 28928
rect 4030 28872 4035 28928
rect 0 28870 4035 28872
rect 0 28840 800 28870
rect 3969 28867 4035 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 4208 28320 4528 28321
rect 0 28250 800 28280
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 2865 28250 2931 28253
rect 0 28248 2931 28250
rect 0 28192 2870 28248
rect 2926 28192 2931 28248
rect 0 28190 2931 28192
rect 0 28160 800 28190
rect 2865 28187 2931 28190
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 0 27570 800 27600
rect 3325 27570 3391 27573
rect 0 27568 3391 27570
rect 0 27512 3330 27568
rect 3386 27512 3391 27568
rect 0 27510 3391 27512
rect 0 27480 800 27510
rect 3325 27507 3391 27510
rect 13629 27570 13695 27573
rect 15285 27570 15351 27573
rect 13629 27568 15351 27570
rect 13629 27512 13634 27568
rect 13690 27512 15290 27568
rect 15346 27512 15351 27568
rect 13629 27510 15351 27512
rect 13629 27507 13695 27510
rect 15285 27507 15351 27510
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 0 26890 800 26920
rect 3417 26890 3483 26893
rect 0 26888 3483 26890
rect 0 26832 3422 26888
rect 3478 26832 3483 26888
rect 0 26830 3483 26832
rect 0 26800 800 26830
rect 3417 26827 3483 26830
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 0 26346 800 26376
rect 3233 26346 3299 26349
rect 0 26344 3299 26346
rect 0 26288 3238 26344
rect 3294 26288 3299 26344
rect 0 26286 3299 26288
rect 0 26256 800 26286
rect 3233 26283 3299 26286
rect 5165 26210 5231 26213
rect 8293 26210 8359 26213
rect 18413 26212 18479 26213
rect 18413 26210 18460 26212
rect 5165 26208 8359 26210
rect 5165 26152 5170 26208
rect 5226 26152 8298 26208
rect 8354 26152 8359 26208
rect 5165 26150 8359 26152
rect 18368 26208 18460 26210
rect 18368 26152 18418 26208
rect 18368 26150 18460 26152
rect 5165 26147 5231 26150
rect 8293 26147 8359 26150
rect 18413 26148 18460 26150
rect 18524 26148 18530 26212
rect 56593 26210 56659 26213
rect 56593 26208 59002 26210
rect 56593 26152 56598 26208
rect 56654 26152 59002 26208
rect 56593 26150 59002 26152
rect 18413 26147 18479 26148
rect 56593 26147 56659 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 31569 26100 31635 26103
rect 31569 26098 32108 26100
rect 31569 26042 31574 26098
rect 31630 26042 32108 26098
rect 58942 26090 59524 26150
rect 31569 26040 32108 26042
rect 83825 26074 83891 26077
rect 83825 26072 86940 26074
rect 31569 26037 31635 26040
rect 83825 26016 83830 26072
rect 83886 26016 86940 26072
rect 83825 26014 86940 26016
rect 83825 26011 83891 26014
rect 0 25666 800 25696
rect 3877 25666 3943 25669
rect 0 25664 3943 25666
rect 0 25608 3882 25664
rect 3938 25608 3943 25664
rect 0 25606 3943 25608
rect 0 25576 800 25606
rect 3877 25603 3943 25606
rect 56685 25666 56751 25669
rect 56685 25664 59002 25666
rect 56685 25608 56690 25664
rect 56746 25608 59002 25664
rect 56685 25606 59002 25608
rect 59353 25606 59419 25609
rect 56685 25603 56751 25606
rect 58942 25604 59524 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 31661 25556 31727 25559
rect 31661 25554 32108 25556
rect 31661 25498 31666 25554
rect 31722 25498 32108 25554
rect 58942 25548 59358 25604
rect 59414 25548 59524 25604
rect 58942 25546 59524 25548
rect 59353 25543 59419 25546
rect 31661 25496 32108 25498
rect 31661 25493 31727 25496
rect 82854 25468 82860 25532
rect 82924 25530 82930 25532
rect 86493 25530 86559 25533
rect 82924 25528 86940 25530
rect 82924 25472 86498 25528
rect 86554 25472 86940 25528
rect 82924 25470 86940 25472
rect 82924 25468 82930 25470
rect 86493 25467 86559 25470
rect 59077 25062 59143 25065
rect 58942 25060 59524 25062
rect 4208 25056 4528 25057
rect 0 24986 800 25016
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 31753 25056 31819 25059
rect 31753 25054 32108 25056
rect 31753 24998 31758 25054
rect 31814 24998 32108 25054
rect 31753 24996 32108 24998
rect 58942 25004 59082 25060
rect 59138 25004 59524 25060
rect 58942 25002 59524 25004
rect 31753 24993 31819 24996
rect 4208 24991 4528 24992
rect 2773 24986 2839 24989
rect 0 24984 2839 24986
rect 0 24928 2778 24984
rect 2834 24928 2839 24984
rect 0 24926 2839 24928
rect 0 24896 800 24926
rect 2773 24923 2839 24926
rect 57462 24924 57468 24988
rect 57532 24986 57538 24988
rect 58942 24986 59002 25002
rect 59077 24999 59143 25002
rect 57532 24926 59002 24986
rect 57532 24924 57538 24926
rect 83590 24924 83596 24988
rect 83660 24986 83666 24988
rect 86677 24986 86743 24989
rect 83660 24984 86940 24986
rect 83660 24928 86682 24984
rect 86738 24928 86940 24984
rect 83660 24926 86940 24928
rect 83660 24924 83666 24926
rect 86677 24923 86743 24926
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 0 24306 800 24336
rect 2957 24306 3023 24309
rect 0 24304 3023 24306
rect 0 24248 2962 24304
rect 3018 24248 3023 24304
rect 0 24246 3023 24248
rect 0 24216 800 24246
rect 2957 24243 3023 24246
rect 26877 24036 26943 24037
rect 26877 24034 26924 24036
rect 26832 24032 26924 24034
rect 26832 23976 26882 24032
rect 26832 23974 26924 23976
rect 26877 23972 26924 23974
rect 26988 23972 26994 24036
rect 26877 23971 26943 23972
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 31569 23968 31635 23971
rect 31569 23966 32108 23968
rect 31569 23910 31574 23966
rect 31630 23910 32108 23966
rect 59353 23918 59419 23921
rect 31569 23908 32108 23910
rect 58942 23916 59524 23918
rect 31569 23905 31635 23908
rect 4208 23903 4528 23904
rect 56542 23836 56548 23900
rect 56612 23898 56618 23900
rect 58942 23898 59358 23916
rect 56612 23860 59358 23898
rect 59414 23860 59524 23916
rect 56612 23858 59524 23860
rect 56612 23838 59002 23858
rect 59353 23855 59419 23858
rect 56612 23836 56618 23838
rect 82854 23836 82860 23900
rect 82924 23898 82930 23900
rect 86309 23898 86375 23901
rect 82924 23896 86940 23898
rect 82924 23840 86314 23896
rect 86370 23840 86940 23896
rect 82924 23838 86940 23840
rect 82924 23836 82930 23838
rect 86309 23835 86375 23838
rect 0 23762 800 23792
rect 4061 23762 4127 23765
rect 0 23760 4127 23762
rect 0 23704 4066 23760
rect 4122 23704 4127 23760
rect 0 23702 4127 23704
rect 0 23672 800 23702
rect 4061 23699 4127 23702
rect 12709 23492 12775 23493
rect 12709 23490 12756 23492
rect 12664 23488 12756 23490
rect 12664 23432 12714 23488
rect 12664 23430 12756 23432
rect 12709 23428 12756 23430
rect 12820 23428 12826 23492
rect 14825 23490 14891 23493
rect 18781 23492 18847 23493
rect 14958 23490 14964 23492
rect 14825 23488 14964 23490
rect 14825 23432 14830 23488
rect 14886 23432 14964 23488
rect 14825 23430 14964 23432
rect 12709 23427 12775 23428
rect 14825 23427 14891 23430
rect 14958 23428 14964 23430
rect 15028 23428 15034 23492
rect 18781 23488 18828 23492
rect 18892 23490 18898 23492
rect 18781 23432 18786 23488
rect 18781 23428 18828 23432
rect 18892 23430 18938 23490
rect 18892 23428 18898 23430
rect 18781 23427 18847 23428
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 0 23082 800 23112
rect 3785 23082 3851 23085
rect 0 23080 3851 23082
rect 0 23024 3790 23080
rect 3846 23024 3851 23080
rect 0 23022 3851 23024
rect 0 22992 800 23022
rect 3785 23019 3851 23022
rect 56910 22884 56916 22948
rect 56980 22946 56986 22948
rect 56980 22886 59186 22946
rect 56980 22884 56986 22886
rect 58985 22884 59524 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 31569 22836 31635 22839
rect 31569 22834 32108 22836
rect 14549 22812 14615 22813
rect 14549 22810 14596 22812
rect 14504 22808 14596 22810
rect 14504 22752 14554 22808
rect 14504 22750 14596 22752
rect 14549 22748 14596 22750
rect 14660 22748 14666 22812
rect 31569 22778 31574 22834
rect 31630 22778 32108 22834
rect 58985 22828 58990 22884
rect 59046 22828 59524 22884
rect 86677 22878 86743 22881
rect 58985 22826 59524 22828
rect 86358 22876 86940 22878
rect 58985 22823 59051 22826
rect 86358 22820 86682 22876
rect 86738 22820 86940 22876
rect 86358 22818 86940 22820
rect 31569 22776 32108 22778
rect 31569 22773 31635 22776
rect 82854 22748 82860 22812
rect 82924 22810 82930 22812
rect 86358 22810 86418 22818
rect 86677 22815 86743 22818
rect 82924 22750 86418 22810
rect 82924 22748 82930 22750
rect 14549 22747 14615 22748
rect 0 22402 800 22432
rect 2865 22402 2931 22405
rect 0 22400 2931 22402
rect 0 22344 2870 22400
rect 2926 22344 2931 22400
rect 0 22342 2931 22344
rect 0 22312 800 22342
rect 2865 22339 2931 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 57789 21858 57855 21861
rect 57789 21856 59002 21858
rect 57789 21800 57794 21856
rect 57850 21800 59002 21856
rect 57789 21798 59002 21800
rect 57789 21795 57855 21798
rect 4208 21792 4528 21793
rect 0 21722 800 21752
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 3141 21722 3207 21725
rect 0 21720 3207 21722
rect 0 21664 3146 21720
rect 3202 21664 3207 21720
rect 0 21662 3207 21664
rect 0 21632 800 21662
rect 3141 21659 3207 21662
rect 28993 21722 29059 21725
rect 31526 21722 32108 21742
rect 58942 21738 59524 21798
rect 86585 21790 86651 21793
rect 86358 21788 86940 21790
rect 86358 21732 86590 21788
rect 86646 21732 86940 21788
rect 86358 21730 86940 21732
rect 28993 21720 32108 21722
rect 28993 21664 28998 21720
rect 29054 21682 32108 21720
rect 29054 21664 31586 21682
rect 28993 21662 31586 21664
rect 28993 21659 29059 21662
rect 82854 21660 82860 21724
rect 82924 21722 82930 21724
rect 86358 21722 86418 21730
rect 86585 21727 86651 21730
rect 82924 21662 86418 21722
rect 82924 21660 82930 21662
rect 25405 21452 25471 21453
rect 25405 21450 25452 21452
rect 25360 21448 25452 21450
rect 25360 21392 25410 21448
rect 25360 21390 25452 21392
rect 25405 21388 25452 21390
rect 25516 21388 25522 21452
rect 57830 21388 57836 21452
rect 57900 21450 57906 21452
rect 59353 21450 59419 21453
rect 57900 21448 59419 21450
rect 57900 21392 59358 21448
rect 59414 21392 59419 21448
rect 57900 21390 59419 21392
rect 57900 21388 57906 21390
rect 25405 21387 25471 21388
rect 59353 21387 59419 21390
rect 14089 21314 14155 21317
rect 14222 21314 14228 21316
rect 14089 21312 14228 21314
rect 14089 21256 14094 21312
rect 14150 21256 14228 21312
rect 14089 21254 14228 21256
rect 14089 21251 14155 21254
rect 14222 21252 14228 21254
rect 14292 21252 14298 21316
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 0 21042 800 21072
rect 4061 21042 4127 21045
rect 0 21040 4127 21042
rect 0 20984 4066 21040
rect 4122 20984 4127 21040
rect 0 20982 4127 20984
rect 0 20952 800 20982
rect 4061 20979 4127 20982
rect 18965 20770 19031 20773
rect 19190 20770 19196 20772
rect 18965 20768 19196 20770
rect 18965 20712 18970 20768
rect 19026 20712 19196 20768
rect 18965 20710 19196 20712
rect 18965 20707 19031 20710
rect 19190 20708 19196 20710
rect 19260 20708 19266 20772
rect 59261 20710 59327 20713
rect 59261 20708 59524 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 28993 20634 29059 20637
rect 31526 20634 32108 20654
rect 59261 20652 59266 20708
rect 59322 20652 59524 20708
rect 86677 20702 86743 20705
rect 59261 20650 59524 20652
rect 86358 20700 86940 20702
rect 59261 20647 59327 20650
rect 86358 20644 86682 20700
rect 86738 20644 86940 20700
rect 86358 20642 86940 20644
rect 28993 20632 32108 20634
rect 28993 20576 28998 20632
rect 29054 20594 32108 20632
rect 29054 20576 31586 20594
rect 28993 20574 31586 20576
rect 28993 20571 29059 20574
rect 83222 20572 83228 20636
rect 83292 20634 83298 20636
rect 86358 20634 86418 20642
rect 86677 20639 86743 20642
rect 83292 20574 86418 20634
rect 83292 20572 83298 20574
rect 0 20498 800 20528
rect 3969 20498 4035 20501
rect 0 20496 4035 20498
rect 0 20440 3974 20496
rect 4030 20440 4035 20496
rect 0 20438 4035 20440
rect 0 20408 800 20438
rect 3969 20435 4035 20438
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 15561 20090 15627 20093
rect 15694 20090 15700 20092
rect 15561 20088 15700 20090
rect 15561 20032 15566 20088
rect 15622 20032 15700 20088
rect 15561 20030 15700 20032
rect 15561 20027 15627 20030
rect 15694 20028 15700 20030
rect 15764 20028 15770 20092
rect 0 19818 800 19848
rect 3877 19818 3943 19821
rect 0 19816 3943 19818
rect 0 19760 3882 19816
rect 3938 19760 3943 19816
rect 0 19758 3943 19760
rect 0 19728 800 19758
rect 3877 19755 3943 19758
rect 59353 19622 59419 19625
rect 59353 19620 59524 19622
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 28901 19546 28967 19549
rect 31526 19546 32108 19566
rect 59353 19564 59358 19620
rect 59414 19564 59524 19620
rect 86677 19614 86743 19617
rect 59353 19562 59524 19564
rect 86358 19612 86940 19614
rect 59353 19559 59419 19562
rect 86358 19556 86682 19612
rect 86738 19556 86940 19612
rect 86358 19554 86940 19556
rect 28901 19544 32108 19546
rect 28901 19488 28906 19544
rect 28962 19506 32108 19544
rect 28962 19488 31586 19506
rect 28901 19486 31586 19488
rect 28901 19483 28967 19486
rect 82854 19484 82860 19548
rect 82924 19546 82930 19548
rect 86358 19546 86418 19554
rect 86677 19551 86743 19554
rect 82924 19486 86418 19546
rect 82924 19484 82930 19486
rect 19149 19412 19215 19413
rect 19149 19410 19196 19412
rect 19104 19408 19196 19410
rect 19104 19352 19154 19408
rect 19104 19350 19196 19352
rect 19149 19348 19196 19350
rect 19260 19348 19266 19412
rect 19149 19347 19215 19348
rect 0 19138 800 19168
rect 3325 19138 3391 19141
rect 0 19136 3391 19138
rect 0 19080 3330 19136
rect 3386 19080 3391 19136
rect 0 19078 3391 19080
rect 0 19048 800 19078
rect 3325 19075 3391 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 4208 18528 4528 18529
rect 0 18458 800 18488
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 3693 18458 3759 18461
rect 0 18456 3759 18458
rect 0 18400 3698 18456
rect 3754 18400 3759 18456
rect 0 18398 3759 18400
rect 0 18368 800 18398
rect 3693 18395 3759 18398
rect 19568 17984 19888 17985
rect 0 17914 800 17944
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4061 17914 4127 17917
rect 0 17912 4127 17914
rect 0 17856 4066 17912
rect 4122 17856 4127 17912
rect 0 17854 4127 17856
rect 0 17824 800 17854
rect 4061 17851 4127 17854
rect 83641 17778 83707 17781
rect 86677 17778 86743 17781
rect 83641 17776 86743 17778
rect 83641 17720 83646 17776
rect 83702 17720 86682 17776
rect 86738 17720 86743 17776
rect 83641 17718 86743 17720
rect 83641 17715 83707 17718
rect 86677 17715 86743 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 86677 17438 86743 17441
rect 86358 17436 86940 17438
rect 59353 17396 59419 17399
rect 58942 17394 59524 17396
rect 4208 17375 4528 17376
rect 28901 17370 28967 17373
rect 31526 17370 32108 17390
rect 28901 17368 32108 17370
rect 28901 17312 28906 17368
rect 28962 17330 32108 17368
rect 28962 17312 31586 17330
rect 28901 17310 31586 17312
rect 28901 17307 28967 17310
rect 53414 17308 53420 17372
rect 53484 17370 53490 17372
rect 58942 17370 59358 17394
rect 53484 17338 59358 17370
rect 59414 17338 59524 17394
rect 86358 17380 86682 17436
rect 86738 17380 86940 17436
rect 86358 17378 86940 17380
rect 53484 17336 59524 17338
rect 53484 17310 59002 17336
rect 59353 17333 59419 17336
rect 53484 17308 53490 17310
rect 83958 17308 83964 17372
rect 84028 17370 84034 17372
rect 86358 17370 86418 17378
rect 86677 17375 86743 17378
rect 84028 17310 86418 17370
rect 84028 17308 84034 17310
rect 0 17234 800 17264
rect 3509 17234 3575 17237
rect 0 17232 3575 17234
rect 0 17176 3514 17232
rect 3570 17176 3575 17232
rect 0 17174 3575 17176
rect 0 17144 800 17174
rect 3509 17171 3575 17174
rect 14181 17098 14247 17101
rect 14958 17098 14964 17100
rect 14181 17096 14964 17098
rect 14181 17040 14186 17096
rect 14242 17040 14964 17096
rect 14181 17038 14964 17040
rect 14181 17035 14247 17038
rect 14958 17036 14964 17038
rect 15028 17036 15034 17100
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 13445 16692 13511 16693
rect 20805 16692 20871 16693
rect 13445 16690 13492 16692
rect 13400 16688 13492 16690
rect 13400 16632 13450 16688
rect 13400 16630 13492 16632
rect 13445 16628 13492 16630
rect 13556 16628 13562 16692
rect 20805 16690 20852 16692
rect 20760 16688 20852 16690
rect 20760 16632 20810 16688
rect 20760 16630 20852 16632
rect 20805 16628 20852 16630
rect 20916 16628 20922 16692
rect 82854 16628 82860 16692
rect 82924 16690 82930 16692
rect 83641 16690 83707 16693
rect 82924 16688 83707 16690
rect 82924 16632 83646 16688
rect 83702 16632 83707 16688
rect 82924 16630 83707 16632
rect 82924 16628 82930 16630
rect 13445 16627 13511 16628
rect 20805 16627 20871 16628
rect 83641 16627 83707 16630
rect 0 16554 800 16584
rect 4061 16554 4127 16557
rect 0 16552 4127 16554
rect 0 16496 4066 16552
rect 4122 16496 4127 16552
rect 0 16494 4127 16496
rect 0 16464 800 16494
rect 4061 16491 4127 16494
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 21265 16010 21331 16013
rect 21398 16010 21404 16012
rect 21265 16008 21404 16010
rect 21265 15952 21270 16008
rect 21326 15952 21404 16008
rect 21265 15950 21404 15952
rect 21265 15947 21331 15950
rect 21398 15948 21404 15950
rect 21468 15948 21474 16012
rect 0 15874 800 15904
rect 3601 15874 3667 15877
rect 0 15872 3667 15874
rect 0 15816 3606 15872
rect 3662 15816 3667 15872
rect 0 15814 3667 15816
rect 0 15784 800 15814
rect 3601 15811 3667 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 53046 15268 53052 15332
rect 53116 15330 53122 15332
rect 59118 15330 59124 15332
rect 53116 15270 59124 15330
rect 53116 15268 53122 15270
rect 59118 15268 59124 15270
rect 59188 15268 59194 15332
rect 4208 15264 4528 15265
rect 0 15194 800 15224
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 4061 15194 4127 15197
rect 0 15192 4127 15194
rect 0 15136 4066 15192
rect 4122 15136 4127 15192
rect 0 15134 4127 15136
rect 0 15104 800 15134
rect 4061 15131 4127 15134
rect 19568 14720 19888 14721
rect 0 14650 800 14680
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 3969 14650 4035 14653
rect 0 14648 4035 14650
rect 0 14592 3974 14648
rect 4030 14592 4035 14648
rect 0 14590 4035 14592
rect 0 14560 800 14590
rect 3969 14587 4035 14590
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 0 13970 800 14000
rect 4061 13970 4127 13973
rect 0 13968 4127 13970
rect 0 13912 4066 13968
rect 4122 13912 4127 13968
rect 0 13910 4127 13912
rect 0 13880 800 13910
rect 4061 13907 4127 13910
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 0 13290 800 13320
rect 3877 13290 3943 13293
rect 0 13288 3943 13290
rect 0 13232 3882 13288
rect 3938 13232 3943 13288
rect 0 13230 3943 13232
rect 0 13200 800 13230
rect 3877 13227 3943 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 31753 13088 31819 13091
rect 31753 13086 32108 13088
rect 31753 13030 31758 13086
rect 31814 13030 32108 13086
rect 59118 13032 59124 13096
rect 59188 13094 59194 13096
rect 59188 13034 59524 13094
rect 59188 13032 59194 13034
rect 31753 13028 32108 13030
rect 31753 13025 31819 13028
rect 4208 13023 4528 13024
rect 86358 13006 86940 13066
rect 83641 12882 83707 12885
rect 86358 12882 86418 13006
rect 83641 12880 86418 12882
rect 83641 12824 83646 12880
rect 83702 12824 86418 12880
rect 83641 12822 86418 12824
rect 83641 12819 83707 12822
rect 0 12610 800 12640
rect 3969 12610 4035 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 0 12520 800 12550
rect 3969 12547 4035 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 0 12066 800 12096
rect 3325 12066 3391 12069
rect 0 12064 3391 12066
rect 0 12008 3330 12064
rect 3386 12008 3391 12064
rect 0 12006 3391 12008
rect 0 11976 800 12006
rect 3325 12003 3391 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 19568 11456 19888 11457
rect 0 11386 800 11416
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 800 11326
rect 3969 11323 4035 11326
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 0 10706 800 10736
rect 3969 10706 4035 10709
rect 0 10704 4035 10706
rect 0 10648 3974 10704
rect 4030 10648 4035 10704
rect 0 10646 4035 10648
rect 0 10616 800 10646
rect 3969 10643 4035 10646
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 0 10026 800 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 800 9966
rect 3969 9963 4035 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 0 9346 800 9376
rect 3509 9346 3575 9349
rect 0 9344 3575 9346
rect 0 9288 3514 9344
rect 3570 9288 3575 9344
rect 0 9286 3575 9288
rect 0 9256 800 9286
rect 3509 9283 3575 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 0 8802 800 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 800 8742
rect 4061 8739 4127 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 19568 8192 19888 8193
rect 0 8122 800 8152
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 3785 8122 3851 8125
rect 0 8120 3851 8122
rect 0 8064 3790 8120
rect 3846 8064 3851 8120
rect 0 8062 3851 8064
rect 0 8032 800 8062
rect 3785 8059 3851 8062
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 0 7442 800 7472
rect 3969 7442 4035 7445
rect 0 7440 4035 7442
rect 0 7384 3974 7440
rect 4030 7384 4035 7440
rect 0 7382 4035 7384
rect 0 7352 800 7382
rect 3969 7379 4035 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 0 6762 800 6792
rect 3969 6762 4035 6765
rect 0 6760 4035 6762
rect 0 6704 3974 6760
rect 4030 6704 4035 6760
rect 0 6702 4035 6704
rect 0 6672 800 6702
rect 3969 6699 4035 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 0 5538 800 5568
rect 3417 5538 3483 5541
rect 0 5536 3483 5538
rect 0 5480 3422 5536
rect 3478 5480 3483 5536
rect 0 5478 3483 5480
rect 0 5448 800 5478
rect 3417 5475 3483 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 19568 4928 19888 4929
rect 0 4858 800 4888
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 800 4798
rect 4061 4795 4127 4798
rect 29913 4858 29979 4861
rect 29913 4856 32138 4858
rect 29913 4800 29918 4856
rect 29974 4800 32138 4856
rect 29913 4798 32138 4800
rect 29913 4795 29979 4798
rect 59494 4725 59554 4848
rect 86358 4846 86940 4906
rect 59494 4720 59603 4725
rect 59494 4664 59542 4720
rect 59598 4664 59603 4720
rect 59494 4662 59603 4664
rect 59537 4659 59603 4662
rect 83917 4722 83983 4725
rect 86358 4722 86418 4846
rect 83917 4720 86418 4722
rect 83917 4664 83922 4720
rect 83978 4664 86418 4720
rect 83917 4662 86418 4664
rect 83917 4659 83983 4662
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 0 4178 800 4208
rect 2957 4178 3023 4181
rect 0 4176 3023 4178
rect 0 4120 2962 4176
rect 3018 4120 3023 4176
rect 0 4118 3023 4120
rect 0 4088 800 4118
rect 2957 4115 3023 4118
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3498 800 3528
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3408 800 3438
rect 4061 3435 4127 3438
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 0 2954 800 2984
rect 3325 2954 3391 2957
rect 0 2952 3391 2954
rect 0 2896 3330 2952
rect 3386 2896 3391 2952
rect 0 2894 3391 2896
rect 0 2864 800 2894
rect 3325 2891 3391 2894
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 0 2274 800 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 800 2214
rect 2865 2211 2931 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 0 1594 800 1624
rect 3233 1594 3299 1597
rect 0 1592 3299 1594
rect 0 1536 3238 1592
rect 3294 1536 3299 1592
rect 0 1534 3299 1536
rect 0 1504 800 1534
rect 3233 1531 3299 1534
rect 0 914 800 944
rect 2773 914 2839 917
rect 0 912 2839 914
rect 0 856 2778 912
rect 2834 856 2839 912
rect 0 854 2839 856
rect 0 824 800 854
rect 2773 851 2839 854
rect 0 370 800 400
rect 3417 370 3483 373
rect 0 368 3483 370
rect 0 312 3422 368
rect 3478 312 3483 368
rect 0 310 3483 312
rect 0 280 800 310
rect 3417 307 3483 310
<< via3 >>
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 65656 47900 65720 47904
rect 65656 47844 65660 47900
rect 65660 47844 65716 47900
rect 65716 47844 65720 47900
rect 65656 47840 65720 47844
rect 65736 47900 65800 47904
rect 65736 47844 65740 47900
rect 65740 47844 65796 47900
rect 65796 47844 65800 47900
rect 65736 47840 65800 47844
rect 65816 47900 65880 47904
rect 65816 47844 65820 47900
rect 65820 47844 65876 47900
rect 65876 47844 65880 47900
rect 65816 47840 65880 47844
rect 65896 47900 65960 47904
rect 65896 47844 65900 47900
rect 65900 47844 65956 47900
rect 65956 47844 65960 47900
rect 65896 47840 65960 47844
rect 96376 47900 96440 47904
rect 96376 47844 96380 47900
rect 96380 47844 96436 47900
rect 96436 47844 96440 47900
rect 96376 47840 96440 47844
rect 96456 47900 96520 47904
rect 96456 47844 96460 47900
rect 96460 47844 96516 47900
rect 96516 47844 96520 47900
rect 96456 47840 96520 47844
rect 96536 47900 96600 47904
rect 96536 47844 96540 47900
rect 96540 47844 96596 47900
rect 96596 47844 96600 47900
rect 96536 47840 96600 47844
rect 96616 47900 96680 47904
rect 96616 47844 96620 47900
rect 96620 47844 96676 47900
rect 96676 47844 96680 47900
rect 96616 47840 96680 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 50296 47356 50360 47360
rect 50296 47300 50300 47356
rect 50300 47300 50356 47356
rect 50356 47300 50360 47356
rect 50296 47296 50360 47300
rect 50376 47356 50440 47360
rect 50376 47300 50380 47356
rect 50380 47300 50436 47356
rect 50436 47300 50440 47356
rect 50376 47296 50440 47300
rect 50456 47356 50520 47360
rect 50456 47300 50460 47356
rect 50460 47300 50516 47356
rect 50516 47300 50520 47356
rect 50456 47296 50520 47300
rect 50536 47356 50600 47360
rect 50536 47300 50540 47356
rect 50540 47300 50596 47356
rect 50596 47300 50600 47356
rect 50536 47296 50600 47300
rect 81016 47356 81080 47360
rect 81016 47300 81020 47356
rect 81020 47300 81076 47356
rect 81076 47300 81080 47356
rect 81016 47296 81080 47300
rect 81096 47356 81160 47360
rect 81096 47300 81100 47356
rect 81100 47300 81156 47356
rect 81156 47300 81160 47356
rect 81096 47296 81160 47300
rect 81176 47356 81240 47360
rect 81176 47300 81180 47356
rect 81180 47300 81236 47356
rect 81236 47300 81240 47356
rect 81176 47296 81240 47300
rect 81256 47356 81320 47360
rect 81256 47300 81260 47356
rect 81260 47300 81316 47356
rect 81316 47300 81320 47356
rect 81256 47296 81320 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 65656 46812 65720 46816
rect 65656 46756 65660 46812
rect 65660 46756 65716 46812
rect 65716 46756 65720 46812
rect 65656 46752 65720 46756
rect 65736 46812 65800 46816
rect 65736 46756 65740 46812
rect 65740 46756 65796 46812
rect 65796 46756 65800 46812
rect 65736 46752 65800 46756
rect 65816 46812 65880 46816
rect 65816 46756 65820 46812
rect 65820 46756 65876 46812
rect 65876 46756 65880 46812
rect 65816 46752 65880 46756
rect 65896 46812 65960 46816
rect 65896 46756 65900 46812
rect 65900 46756 65956 46812
rect 65956 46756 65960 46812
rect 65896 46752 65960 46756
rect 96376 46812 96440 46816
rect 96376 46756 96380 46812
rect 96380 46756 96436 46812
rect 96436 46756 96440 46812
rect 96376 46752 96440 46756
rect 96456 46812 96520 46816
rect 96456 46756 96460 46812
rect 96460 46756 96516 46812
rect 96516 46756 96520 46812
rect 96456 46752 96520 46756
rect 96536 46812 96600 46816
rect 96536 46756 96540 46812
rect 96540 46756 96596 46812
rect 96596 46756 96600 46812
rect 96536 46752 96600 46756
rect 96616 46812 96680 46816
rect 96616 46756 96620 46812
rect 96620 46756 96676 46812
rect 96676 46756 96680 46812
rect 96616 46752 96680 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 50296 46268 50360 46272
rect 50296 46212 50300 46268
rect 50300 46212 50356 46268
rect 50356 46212 50360 46268
rect 50296 46208 50360 46212
rect 50376 46268 50440 46272
rect 50376 46212 50380 46268
rect 50380 46212 50436 46268
rect 50436 46212 50440 46268
rect 50376 46208 50440 46212
rect 50456 46268 50520 46272
rect 50456 46212 50460 46268
rect 50460 46212 50516 46268
rect 50516 46212 50520 46268
rect 50456 46208 50520 46212
rect 50536 46268 50600 46272
rect 50536 46212 50540 46268
rect 50540 46212 50596 46268
rect 50596 46212 50600 46268
rect 50536 46208 50600 46212
rect 81016 46268 81080 46272
rect 81016 46212 81020 46268
rect 81020 46212 81076 46268
rect 81076 46212 81080 46268
rect 81016 46208 81080 46212
rect 81096 46268 81160 46272
rect 81096 46212 81100 46268
rect 81100 46212 81156 46268
rect 81156 46212 81160 46268
rect 81096 46208 81160 46212
rect 81176 46268 81240 46272
rect 81176 46212 81180 46268
rect 81180 46212 81236 46268
rect 81236 46212 81240 46268
rect 81176 46208 81240 46212
rect 81256 46268 81320 46272
rect 81256 46212 81260 46268
rect 81260 46212 81316 46268
rect 81316 46212 81320 46268
rect 81256 46208 81320 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 65656 45724 65720 45728
rect 65656 45668 65660 45724
rect 65660 45668 65716 45724
rect 65716 45668 65720 45724
rect 65656 45664 65720 45668
rect 65736 45724 65800 45728
rect 65736 45668 65740 45724
rect 65740 45668 65796 45724
rect 65796 45668 65800 45724
rect 65736 45664 65800 45668
rect 65816 45724 65880 45728
rect 65816 45668 65820 45724
rect 65820 45668 65876 45724
rect 65876 45668 65880 45724
rect 65816 45664 65880 45668
rect 65896 45724 65960 45728
rect 65896 45668 65900 45724
rect 65900 45668 65956 45724
rect 65956 45668 65960 45724
rect 65896 45664 65960 45668
rect 96376 45724 96440 45728
rect 96376 45668 96380 45724
rect 96380 45668 96436 45724
rect 96436 45668 96440 45724
rect 96376 45664 96440 45668
rect 96456 45724 96520 45728
rect 96456 45668 96460 45724
rect 96460 45668 96516 45724
rect 96516 45668 96520 45724
rect 96456 45664 96520 45668
rect 96536 45724 96600 45728
rect 96536 45668 96540 45724
rect 96540 45668 96596 45724
rect 96596 45668 96600 45724
rect 96536 45664 96600 45668
rect 96616 45724 96680 45728
rect 96616 45668 96620 45724
rect 96620 45668 96676 45724
rect 96676 45668 96680 45724
rect 96616 45664 96680 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 50296 45180 50360 45184
rect 50296 45124 50300 45180
rect 50300 45124 50356 45180
rect 50356 45124 50360 45180
rect 50296 45120 50360 45124
rect 50376 45180 50440 45184
rect 50376 45124 50380 45180
rect 50380 45124 50436 45180
rect 50436 45124 50440 45180
rect 50376 45120 50440 45124
rect 50456 45180 50520 45184
rect 50456 45124 50460 45180
rect 50460 45124 50516 45180
rect 50516 45124 50520 45180
rect 50456 45120 50520 45124
rect 50536 45180 50600 45184
rect 50536 45124 50540 45180
rect 50540 45124 50596 45180
rect 50596 45124 50600 45180
rect 50536 45120 50600 45124
rect 81016 45180 81080 45184
rect 81016 45124 81020 45180
rect 81020 45124 81076 45180
rect 81076 45124 81080 45180
rect 81016 45120 81080 45124
rect 81096 45180 81160 45184
rect 81096 45124 81100 45180
rect 81100 45124 81156 45180
rect 81156 45124 81160 45180
rect 81096 45120 81160 45124
rect 81176 45180 81240 45184
rect 81176 45124 81180 45180
rect 81180 45124 81236 45180
rect 81236 45124 81240 45180
rect 81176 45120 81240 45124
rect 81256 45180 81320 45184
rect 81256 45124 81260 45180
rect 81260 45124 81316 45180
rect 81316 45124 81320 45180
rect 81256 45120 81320 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 65656 44636 65720 44640
rect 65656 44580 65660 44636
rect 65660 44580 65716 44636
rect 65716 44580 65720 44636
rect 65656 44576 65720 44580
rect 65736 44636 65800 44640
rect 65736 44580 65740 44636
rect 65740 44580 65796 44636
rect 65796 44580 65800 44636
rect 65736 44576 65800 44580
rect 65816 44636 65880 44640
rect 65816 44580 65820 44636
rect 65820 44580 65876 44636
rect 65876 44580 65880 44636
rect 65816 44576 65880 44580
rect 65896 44636 65960 44640
rect 65896 44580 65900 44636
rect 65900 44580 65956 44636
rect 65956 44580 65960 44636
rect 65896 44576 65960 44580
rect 96376 44636 96440 44640
rect 96376 44580 96380 44636
rect 96380 44580 96436 44636
rect 96436 44580 96440 44636
rect 96376 44576 96440 44580
rect 96456 44636 96520 44640
rect 96456 44580 96460 44636
rect 96460 44580 96516 44636
rect 96516 44580 96520 44636
rect 96456 44576 96520 44580
rect 96536 44636 96600 44640
rect 96536 44580 96540 44636
rect 96540 44580 96596 44636
rect 96596 44580 96600 44636
rect 96536 44576 96600 44580
rect 96616 44636 96680 44640
rect 96616 44580 96620 44636
rect 96620 44580 96676 44636
rect 96676 44580 96680 44636
rect 96616 44576 96680 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 81016 44092 81080 44096
rect 81016 44036 81020 44092
rect 81020 44036 81076 44092
rect 81076 44036 81080 44092
rect 81016 44032 81080 44036
rect 81096 44092 81160 44096
rect 81096 44036 81100 44092
rect 81100 44036 81156 44092
rect 81156 44036 81160 44092
rect 81096 44032 81160 44036
rect 81176 44092 81240 44096
rect 81176 44036 81180 44092
rect 81180 44036 81236 44092
rect 81236 44036 81240 44092
rect 81176 44032 81240 44036
rect 81256 44092 81320 44096
rect 81256 44036 81260 44092
rect 81260 44036 81316 44092
rect 81316 44036 81320 44092
rect 81256 44032 81320 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 65656 43548 65720 43552
rect 65656 43492 65660 43548
rect 65660 43492 65716 43548
rect 65716 43492 65720 43548
rect 65656 43488 65720 43492
rect 65736 43548 65800 43552
rect 65736 43492 65740 43548
rect 65740 43492 65796 43548
rect 65796 43492 65800 43548
rect 65736 43488 65800 43492
rect 65816 43548 65880 43552
rect 65816 43492 65820 43548
rect 65820 43492 65876 43548
rect 65876 43492 65880 43548
rect 65816 43488 65880 43492
rect 65896 43548 65960 43552
rect 65896 43492 65900 43548
rect 65900 43492 65956 43548
rect 65956 43492 65960 43548
rect 65896 43488 65960 43492
rect 96376 43548 96440 43552
rect 96376 43492 96380 43548
rect 96380 43492 96436 43548
rect 96436 43492 96440 43548
rect 96376 43488 96440 43492
rect 96456 43548 96520 43552
rect 96456 43492 96460 43548
rect 96460 43492 96516 43548
rect 96516 43492 96520 43548
rect 96456 43488 96520 43492
rect 96536 43548 96600 43552
rect 96536 43492 96540 43548
rect 96540 43492 96596 43548
rect 96596 43492 96600 43548
rect 96536 43488 96600 43492
rect 96616 43548 96680 43552
rect 96616 43492 96620 43548
rect 96620 43492 96676 43548
rect 96676 43492 96680 43548
rect 96616 43488 96680 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 81016 43004 81080 43008
rect 81016 42948 81020 43004
rect 81020 42948 81076 43004
rect 81076 42948 81080 43004
rect 81016 42944 81080 42948
rect 81096 43004 81160 43008
rect 81096 42948 81100 43004
rect 81100 42948 81156 43004
rect 81156 42948 81160 43004
rect 81096 42944 81160 42948
rect 81176 43004 81240 43008
rect 81176 42948 81180 43004
rect 81180 42948 81236 43004
rect 81236 42948 81240 43004
rect 81176 42944 81240 42948
rect 81256 43004 81320 43008
rect 81256 42948 81260 43004
rect 81260 42948 81316 43004
rect 81316 42948 81320 43004
rect 81256 42944 81320 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 65656 42460 65720 42464
rect 65656 42404 65660 42460
rect 65660 42404 65716 42460
rect 65716 42404 65720 42460
rect 65656 42400 65720 42404
rect 65736 42460 65800 42464
rect 65736 42404 65740 42460
rect 65740 42404 65796 42460
rect 65796 42404 65800 42460
rect 65736 42400 65800 42404
rect 65816 42460 65880 42464
rect 65816 42404 65820 42460
rect 65820 42404 65876 42460
rect 65876 42404 65880 42460
rect 65816 42400 65880 42404
rect 65896 42460 65960 42464
rect 65896 42404 65900 42460
rect 65900 42404 65956 42460
rect 65956 42404 65960 42460
rect 65896 42400 65960 42404
rect 96376 42460 96440 42464
rect 96376 42404 96380 42460
rect 96380 42404 96436 42460
rect 96436 42404 96440 42460
rect 96376 42400 96440 42404
rect 96456 42460 96520 42464
rect 96456 42404 96460 42460
rect 96460 42404 96516 42460
rect 96516 42404 96520 42460
rect 96456 42400 96520 42404
rect 96536 42460 96600 42464
rect 96536 42404 96540 42460
rect 96540 42404 96596 42460
rect 96596 42404 96600 42460
rect 96536 42400 96600 42404
rect 96616 42460 96680 42464
rect 96616 42404 96620 42460
rect 96620 42404 96676 42460
rect 96676 42404 96680 42460
rect 96616 42400 96680 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 81016 41916 81080 41920
rect 81016 41860 81020 41916
rect 81020 41860 81076 41916
rect 81076 41860 81080 41916
rect 81016 41856 81080 41860
rect 81096 41916 81160 41920
rect 81096 41860 81100 41916
rect 81100 41860 81156 41916
rect 81156 41860 81160 41916
rect 81096 41856 81160 41860
rect 81176 41916 81240 41920
rect 81176 41860 81180 41916
rect 81180 41860 81236 41916
rect 81236 41860 81240 41916
rect 81176 41856 81240 41860
rect 81256 41916 81320 41920
rect 81256 41860 81260 41916
rect 81260 41860 81316 41916
rect 81316 41860 81320 41916
rect 81256 41856 81320 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 65656 41372 65720 41376
rect 65656 41316 65660 41372
rect 65660 41316 65716 41372
rect 65716 41316 65720 41372
rect 65656 41312 65720 41316
rect 65736 41372 65800 41376
rect 65736 41316 65740 41372
rect 65740 41316 65796 41372
rect 65796 41316 65800 41372
rect 65736 41312 65800 41316
rect 65816 41372 65880 41376
rect 65816 41316 65820 41372
rect 65820 41316 65876 41372
rect 65876 41316 65880 41372
rect 65816 41312 65880 41316
rect 65896 41372 65960 41376
rect 65896 41316 65900 41372
rect 65900 41316 65956 41372
rect 65956 41316 65960 41372
rect 65896 41312 65960 41316
rect 96376 41372 96440 41376
rect 96376 41316 96380 41372
rect 96380 41316 96436 41372
rect 96436 41316 96440 41372
rect 96376 41312 96440 41316
rect 96456 41372 96520 41376
rect 96456 41316 96460 41372
rect 96460 41316 96516 41372
rect 96516 41316 96520 41372
rect 96456 41312 96520 41316
rect 96536 41372 96600 41376
rect 96536 41316 96540 41372
rect 96540 41316 96596 41372
rect 96596 41316 96600 41372
rect 96536 41312 96600 41316
rect 96616 41372 96680 41376
rect 96616 41316 96620 41372
rect 96620 41316 96676 41372
rect 96676 41316 96680 41372
rect 96616 41312 96680 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 81016 40828 81080 40832
rect 81016 40772 81020 40828
rect 81020 40772 81076 40828
rect 81076 40772 81080 40828
rect 81016 40768 81080 40772
rect 81096 40828 81160 40832
rect 81096 40772 81100 40828
rect 81100 40772 81156 40828
rect 81156 40772 81160 40828
rect 81096 40768 81160 40772
rect 81176 40828 81240 40832
rect 81176 40772 81180 40828
rect 81180 40772 81236 40828
rect 81236 40772 81240 40828
rect 81176 40768 81240 40772
rect 81256 40828 81320 40832
rect 81256 40772 81260 40828
rect 81260 40772 81316 40828
rect 81316 40772 81320 40828
rect 81256 40768 81320 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 65656 40284 65720 40288
rect 65656 40228 65660 40284
rect 65660 40228 65716 40284
rect 65716 40228 65720 40284
rect 65656 40224 65720 40228
rect 65736 40284 65800 40288
rect 65736 40228 65740 40284
rect 65740 40228 65796 40284
rect 65796 40228 65800 40284
rect 65736 40224 65800 40228
rect 65816 40284 65880 40288
rect 65816 40228 65820 40284
rect 65820 40228 65876 40284
rect 65876 40228 65880 40284
rect 65816 40224 65880 40228
rect 65896 40284 65960 40288
rect 65896 40228 65900 40284
rect 65900 40228 65956 40284
rect 65956 40228 65960 40284
rect 65896 40224 65960 40228
rect 96376 40284 96440 40288
rect 96376 40228 96380 40284
rect 96380 40228 96436 40284
rect 96436 40228 96440 40284
rect 96376 40224 96440 40228
rect 96456 40284 96520 40288
rect 96456 40228 96460 40284
rect 96460 40228 96516 40284
rect 96516 40228 96520 40284
rect 96456 40224 96520 40228
rect 96536 40284 96600 40288
rect 96536 40228 96540 40284
rect 96540 40228 96596 40284
rect 96596 40228 96600 40284
rect 96536 40224 96600 40228
rect 96616 40284 96680 40288
rect 96616 40228 96620 40284
rect 96620 40228 96676 40284
rect 96676 40228 96680 40284
rect 96616 40224 96680 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 81016 39740 81080 39744
rect 81016 39684 81020 39740
rect 81020 39684 81076 39740
rect 81076 39684 81080 39740
rect 81016 39680 81080 39684
rect 81096 39740 81160 39744
rect 81096 39684 81100 39740
rect 81100 39684 81156 39740
rect 81156 39684 81160 39740
rect 81096 39680 81160 39684
rect 81176 39740 81240 39744
rect 81176 39684 81180 39740
rect 81180 39684 81236 39740
rect 81236 39684 81240 39740
rect 81176 39680 81240 39684
rect 81256 39740 81320 39744
rect 81256 39684 81260 39740
rect 81260 39684 81316 39740
rect 81316 39684 81320 39740
rect 81256 39680 81320 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 65656 39196 65720 39200
rect 65656 39140 65660 39196
rect 65660 39140 65716 39196
rect 65716 39140 65720 39196
rect 65656 39136 65720 39140
rect 65736 39196 65800 39200
rect 65736 39140 65740 39196
rect 65740 39140 65796 39196
rect 65796 39140 65800 39196
rect 65736 39136 65800 39140
rect 65816 39196 65880 39200
rect 65816 39140 65820 39196
rect 65820 39140 65876 39196
rect 65876 39140 65880 39196
rect 65816 39136 65880 39140
rect 65896 39196 65960 39200
rect 65896 39140 65900 39196
rect 65900 39140 65956 39196
rect 65956 39140 65960 39196
rect 65896 39136 65960 39140
rect 96376 39196 96440 39200
rect 96376 39140 96380 39196
rect 96380 39140 96436 39196
rect 96436 39140 96440 39196
rect 96376 39136 96440 39140
rect 96456 39196 96520 39200
rect 96456 39140 96460 39196
rect 96460 39140 96516 39196
rect 96516 39140 96520 39196
rect 96456 39136 96520 39140
rect 96536 39196 96600 39200
rect 96536 39140 96540 39196
rect 96540 39140 96596 39196
rect 96596 39140 96600 39196
rect 96536 39136 96600 39140
rect 96616 39196 96680 39200
rect 96616 39140 96620 39196
rect 96620 39140 96676 39196
rect 96676 39140 96680 39196
rect 96616 39136 96680 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 81016 38652 81080 38656
rect 81016 38596 81020 38652
rect 81020 38596 81076 38652
rect 81076 38596 81080 38652
rect 81016 38592 81080 38596
rect 81096 38652 81160 38656
rect 81096 38596 81100 38652
rect 81100 38596 81156 38652
rect 81156 38596 81160 38652
rect 81096 38592 81160 38596
rect 81176 38652 81240 38656
rect 81176 38596 81180 38652
rect 81180 38596 81236 38652
rect 81236 38596 81240 38652
rect 81176 38592 81240 38596
rect 81256 38652 81320 38656
rect 81256 38596 81260 38652
rect 81260 38596 81316 38652
rect 81316 38596 81320 38652
rect 81256 38592 81320 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 65656 38108 65720 38112
rect 65656 38052 65660 38108
rect 65660 38052 65716 38108
rect 65716 38052 65720 38108
rect 65656 38048 65720 38052
rect 65736 38108 65800 38112
rect 65736 38052 65740 38108
rect 65740 38052 65796 38108
rect 65796 38052 65800 38108
rect 65736 38048 65800 38052
rect 65816 38108 65880 38112
rect 65816 38052 65820 38108
rect 65820 38052 65876 38108
rect 65876 38052 65880 38108
rect 65816 38048 65880 38052
rect 65896 38108 65960 38112
rect 65896 38052 65900 38108
rect 65900 38052 65956 38108
rect 65956 38052 65960 38108
rect 65896 38048 65960 38052
rect 96376 38108 96440 38112
rect 96376 38052 96380 38108
rect 96380 38052 96436 38108
rect 96436 38052 96440 38108
rect 96376 38048 96440 38052
rect 96456 38108 96520 38112
rect 96456 38052 96460 38108
rect 96460 38052 96516 38108
rect 96516 38052 96520 38108
rect 96456 38048 96520 38052
rect 96536 38108 96600 38112
rect 96536 38052 96540 38108
rect 96540 38052 96596 38108
rect 96596 38052 96600 38108
rect 96536 38048 96600 38052
rect 96616 38108 96680 38112
rect 96616 38052 96620 38108
rect 96620 38052 96676 38108
rect 96676 38052 96680 38108
rect 96616 38048 96680 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 81016 37564 81080 37568
rect 81016 37508 81020 37564
rect 81020 37508 81076 37564
rect 81076 37508 81080 37564
rect 81016 37504 81080 37508
rect 81096 37564 81160 37568
rect 81096 37508 81100 37564
rect 81100 37508 81156 37564
rect 81156 37508 81160 37564
rect 81096 37504 81160 37508
rect 81176 37564 81240 37568
rect 81176 37508 81180 37564
rect 81180 37508 81236 37564
rect 81236 37508 81240 37564
rect 81176 37504 81240 37508
rect 81256 37564 81320 37568
rect 81256 37508 81260 37564
rect 81260 37508 81316 37564
rect 81316 37508 81320 37564
rect 81256 37504 81320 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 65656 37020 65720 37024
rect 65656 36964 65660 37020
rect 65660 36964 65716 37020
rect 65716 36964 65720 37020
rect 65656 36960 65720 36964
rect 65736 37020 65800 37024
rect 65736 36964 65740 37020
rect 65740 36964 65796 37020
rect 65796 36964 65800 37020
rect 65736 36960 65800 36964
rect 65816 37020 65880 37024
rect 65816 36964 65820 37020
rect 65820 36964 65876 37020
rect 65876 36964 65880 37020
rect 65816 36960 65880 36964
rect 65896 37020 65960 37024
rect 65896 36964 65900 37020
rect 65900 36964 65956 37020
rect 65956 36964 65960 37020
rect 65896 36960 65960 36964
rect 96376 37020 96440 37024
rect 96376 36964 96380 37020
rect 96380 36964 96436 37020
rect 96436 36964 96440 37020
rect 96376 36960 96440 36964
rect 96456 37020 96520 37024
rect 96456 36964 96460 37020
rect 96460 36964 96516 37020
rect 96516 36964 96520 37020
rect 96456 36960 96520 36964
rect 96536 37020 96600 37024
rect 96536 36964 96540 37020
rect 96540 36964 96596 37020
rect 96596 36964 96600 37020
rect 96536 36960 96600 36964
rect 96616 37020 96680 37024
rect 96616 36964 96620 37020
rect 96620 36964 96676 37020
rect 96676 36964 96680 37020
rect 96616 36960 96680 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 81016 36476 81080 36480
rect 81016 36420 81020 36476
rect 81020 36420 81076 36476
rect 81076 36420 81080 36476
rect 81016 36416 81080 36420
rect 81096 36476 81160 36480
rect 81096 36420 81100 36476
rect 81100 36420 81156 36476
rect 81156 36420 81160 36476
rect 81096 36416 81160 36420
rect 81176 36476 81240 36480
rect 81176 36420 81180 36476
rect 81180 36420 81236 36476
rect 81236 36420 81240 36476
rect 81176 36416 81240 36420
rect 81256 36476 81320 36480
rect 81256 36420 81260 36476
rect 81260 36420 81316 36476
rect 81316 36420 81320 36476
rect 81256 36416 81320 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 65656 35932 65720 35936
rect 65656 35876 65660 35932
rect 65660 35876 65716 35932
rect 65716 35876 65720 35932
rect 65656 35872 65720 35876
rect 65736 35932 65800 35936
rect 65736 35876 65740 35932
rect 65740 35876 65796 35932
rect 65796 35876 65800 35932
rect 65736 35872 65800 35876
rect 65816 35932 65880 35936
rect 65816 35876 65820 35932
rect 65820 35876 65876 35932
rect 65876 35876 65880 35932
rect 65816 35872 65880 35876
rect 65896 35932 65960 35936
rect 65896 35876 65900 35932
rect 65900 35876 65956 35932
rect 65956 35876 65960 35932
rect 65896 35872 65960 35876
rect 96376 35932 96440 35936
rect 96376 35876 96380 35932
rect 96380 35876 96436 35932
rect 96436 35876 96440 35932
rect 96376 35872 96440 35876
rect 96456 35932 96520 35936
rect 96456 35876 96460 35932
rect 96460 35876 96516 35932
rect 96516 35876 96520 35932
rect 96456 35872 96520 35876
rect 96536 35932 96600 35936
rect 96536 35876 96540 35932
rect 96540 35876 96596 35932
rect 96596 35876 96600 35932
rect 96536 35872 96600 35876
rect 96616 35932 96680 35936
rect 96616 35876 96620 35932
rect 96620 35876 96676 35932
rect 96676 35876 96680 35932
rect 96616 35872 96680 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 81016 35388 81080 35392
rect 81016 35332 81020 35388
rect 81020 35332 81076 35388
rect 81076 35332 81080 35388
rect 81016 35328 81080 35332
rect 81096 35388 81160 35392
rect 81096 35332 81100 35388
rect 81100 35332 81156 35388
rect 81156 35332 81160 35388
rect 81096 35328 81160 35332
rect 81176 35388 81240 35392
rect 81176 35332 81180 35388
rect 81180 35332 81236 35388
rect 81236 35332 81240 35388
rect 81176 35328 81240 35332
rect 81256 35388 81320 35392
rect 81256 35332 81260 35388
rect 81260 35332 81316 35388
rect 81316 35332 81320 35388
rect 81256 35328 81320 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 65656 34844 65720 34848
rect 65656 34788 65660 34844
rect 65660 34788 65716 34844
rect 65716 34788 65720 34844
rect 65656 34784 65720 34788
rect 65736 34844 65800 34848
rect 65736 34788 65740 34844
rect 65740 34788 65796 34844
rect 65796 34788 65800 34844
rect 65736 34784 65800 34788
rect 65816 34844 65880 34848
rect 65816 34788 65820 34844
rect 65820 34788 65876 34844
rect 65876 34788 65880 34844
rect 65816 34784 65880 34788
rect 65896 34844 65960 34848
rect 65896 34788 65900 34844
rect 65900 34788 65956 34844
rect 65956 34788 65960 34844
rect 65896 34784 65960 34788
rect 96376 34844 96440 34848
rect 96376 34788 96380 34844
rect 96380 34788 96436 34844
rect 96436 34788 96440 34844
rect 96376 34784 96440 34788
rect 96456 34844 96520 34848
rect 96456 34788 96460 34844
rect 96460 34788 96516 34844
rect 96516 34788 96520 34844
rect 96456 34784 96520 34788
rect 96536 34844 96600 34848
rect 96536 34788 96540 34844
rect 96540 34788 96596 34844
rect 96596 34788 96600 34844
rect 96536 34784 96600 34788
rect 96616 34844 96680 34848
rect 96616 34788 96620 34844
rect 96620 34788 96676 34844
rect 96676 34788 96680 34844
rect 96616 34784 96680 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 81016 34300 81080 34304
rect 81016 34244 81020 34300
rect 81020 34244 81076 34300
rect 81076 34244 81080 34300
rect 81016 34240 81080 34244
rect 81096 34300 81160 34304
rect 81096 34244 81100 34300
rect 81100 34244 81156 34300
rect 81156 34244 81160 34300
rect 81096 34240 81160 34244
rect 81176 34300 81240 34304
rect 81176 34244 81180 34300
rect 81180 34244 81236 34300
rect 81236 34244 81240 34300
rect 81176 34240 81240 34244
rect 81256 34300 81320 34304
rect 81256 34244 81260 34300
rect 81260 34244 81316 34300
rect 81316 34244 81320 34300
rect 81256 34240 81320 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 65656 33756 65720 33760
rect 65656 33700 65660 33756
rect 65660 33700 65716 33756
rect 65716 33700 65720 33756
rect 65656 33696 65720 33700
rect 65736 33756 65800 33760
rect 65736 33700 65740 33756
rect 65740 33700 65796 33756
rect 65796 33700 65800 33756
rect 65736 33696 65800 33700
rect 65816 33756 65880 33760
rect 65816 33700 65820 33756
rect 65820 33700 65876 33756
rect 65876 33700 65880 33756
rect 65816 33696 65880 33700
rect 65896 33756 65960 33760
rect 65896 33700 65900 33756
rect 65900 33700 65956 33756
rect 65956 33700 65960 33756
rect 65896 33696 65960 33700
rect 96376 33756 96440 33760
rect 96376 33700 96380 33756
rect 96380 33700 96436 33756
rect 96436 33700 96440 33756
rect 96376 33696 96440 33700
rect 96456 33756 96520 33760
rect 96456 33700 96460 33756
rect 96460 33700 96516 33756
rect 96516 33700 96520 33756
rect 96456 33696 96520 33700
rect 96536 33756 96600 33760
rect 96536 33700 96540 33756
rect 96540 33700 96596 33756
rect 96596 33700 96600 33756
rect 96536 33696 96600 33700
rect 96616 33756 96680 33760
rect 96616 33700 96620 33756
rect 96620 33700 96676 33756
rect 96676 33700 96680 33756
rect 96616 33696 96680 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 50296 33212 50360 33216
rect 50296 33156 50300 33212
rect 50300 33156 50356 33212
rect 50356 33156 50360 33212
rect 50296 33152 50360 33156
rect 50376 33212 50440 33216
rect 50376 33156 50380 33212
rect 50380 33156 50436 33212
rect 50436 33156 50440 33212
rect 50376 33152 50440 33156
rect 50456 33212 50520 33216
rect 50456 33156 50460 33212
rect 50460 33156 50516 33212
rect 50516 33156 50520 33212
rect 50456 33152 50520 33156
rect 50536 33212 50600 33216
rect 50536 33156 50540 33212
rect 50540 33156 50596 33212
rect 50596 33156 50600 33212
rect 50536 33152 50600 33156
rect 81016 33212 81080 33216
rect 81016 33156 81020 33212
rect 81020 33156 81076 33212
rect 81076 33156 81080 33212
rect 81016 33152 81080 33156
rect 81096 33212 81160 33216
rect 81096 33156 81100 33212
rect 81100 33156 81156 33212
rect 81156 33156 81160 33212
rect 81096 33152 81160 33156
rect 81176 33212 81240 33216
rect 81176 33156 81180 33212
rect 81180 33156 81236 33212
rect 81236 33156 81240 33212
rect 81176 33152 81240 33156
rect 81256 33212 81320 33216
rect 81256 33156 81260 33212
rect 81260 33156 81316 33212
rect 81316 33156 81320 33212
rect 81256 33152 81320 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 65656 32668 65720 32672
rect 65656 32612 65660 32668
rect 65660 32612 65716 32668
rect 65716 32612 65720 32668
rect 65656 32608 65720 32612
rect 65736 32668 65800 32672
rect 65736 32612 65740 32668
rect 65740 32612 65796 32668
rect 65796 32612 65800 32668
rect 65736 32608 65800 32612
rect 65816 32668 65880 32672
rect 65816 32612 65820 32668
rect 65820 32612 65876 32668
rect 65876 32612 65880 32668
rect 65816 32608 65880 32612
rect 65896 32668 65960 32672
rect 65896 32612 65900 32668
rect 65900 32612 65956 32668
rect 65956 32612 65960 32668
rect 65896 32608 65960 32612
rect 96376 32668 96440 32672
rect 96376 32612 96380 32668
rect 96380 32612 96436 32668
rect 96436 32612 96440 32668
rect 96376 32608 96440 32612
rect 96456 32668 96520 32672
rect 96456 32612 96460 32668
rect 96460 32612 96516 32668
rect 96516 32612 96520 32668
rect 96456 32608 96520 32612
rect 96536 32668 96600 32672
rect 96536 32612 96540 32668
rect 96540 32612 96596 32668
rect 96596 32612 96600 32668
rect 96536 32608 96600 32612
rect 96616 32668 96680 32672
rect 96616 32612 96620 32668
rect 96620 32612 96676 32668
rect 96676 32612 96680 32668
rect 96616 32608 96680 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 50296 32124 50360 32128
rect 50296 32068 50300 32124
rect 50300 32068 50356 32124
rect 50356 32068 50360 32124
rect 50296 32064 50360 32068
rect 50376 32124 50440 32128
rect 50376 32068 50380 32124
rect 50380 32068 50436 32124
rect 50436 32068 50440 32124
rect 50376 32064 50440 32068
rect 50456 32124 50520 32128
rect 50456 32068 50460 32124
rect 50460 32068 50516 32124
rect 50516 32068 50520 32124
rect 50456 32064 50520 32068
rect 50536 32124 50600 32128
rect 50536 32068 50540 32124
rect 50540 32068 50596 32124
rect 50596 32068 50600 32124
rect 50536 32064 50600 32068
rect 81016 32124 81080 32128
rect 81016 32068 81020 32124
rect 81020 32068 81076 32124
rect 81076 32068 81080 32124
rect 81016 32064 81080 32068
rect 81096 32124 81160 32128
rect 81096 32068 81100 32124
rect 81100 32068 81156 32124
rect 81156 32068 81160 32124
rect 81096 32064 81160 32068
rect 81176 32124 81240 32128
rect 81176 32068 81180 32124
rect 81180 32068 81236 32124
rect 81236 32068 81240 32124
rect 81176 32064 81240 32068
rect 81256 32124 81320 32128
rect 81256 32068 81260 32124
rect 81260 32068 81316 32124
rect 81316 32068 81320 32124
rect 81256 32064 81320 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 65656 31580 65720 31584
rect 65656 31524 65660 31580
rect 65660 31524 65716 31580
rect 65716 31524 65720 31580
rect 65656 31520 65720 31524
rect 65736 31580 65800 31584
rect 65736 31524 65740 31580
rect 65740 31524 65796 31580
rect 65796 31524 65800 31580
rect 65736 31520 65800 31524
rect 65816 31580 65880 31584
rect 65816 31524 65820 31580
rect 65820 31524 65876 31580
rect 65876 31524 65880 31580
rect 65816 31520 65880 31524
rect 65896 31580 65960 31584
rect 65896 31524 65900 31580
rect 65900 31524 65956 31580
rect 65956 31524 65960 31580
rect 65896 31520 65960 31524
rect 96376 31580 96440 31584
rect 96376 31524 96380 31580
rect 96380 31524 96436 31580
rect 96436 31524 96440 31580
rect 96376 31520 96440 31524
rect 96456 31580 96520 31584
rect 96456 31524 96460 31580
rect 96460 31524 96516 31580
rect 96516 31524 96520 31580
rect 96456 31520 96520 31524
rect 96536 31580 96600 31584
rect 96536 31524 96540 31580
rect 96540 31524 96596 31580
rect 96596 31524 96600 31580
rect 96536 31520 96600 31524
rect 96616 31580 96680 31584
rect 96616 31524 96620 31580
rect 96620 31524 96676 31580
rect 96676 31524 96680 31580
rect 96616 31520 96680 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 50296 31036 50360 31040
rect 50296 30980 50300 31036
rect 50300 30980 50356 31036
rect 50356 30980 50360 31036
rect 50296 30976 50360 30980
rect 50376 31036 50440 31040
rect 50376 30980 50380 31036
rect 50380 30980 50436 31036
rect 50436 30980 50440 31036
rect 50376 30976 50440 30980
rect 50456 31036 50520 31040
rect 50456 30980 50460 31036
rect 50460 30980 50516 31036
rect 50516 30980 50520 31036
rect 50456 30976 50520 30980
rect 50536 31036 50600 31040
rect 50536 30980 50540 31036
rect 50540 30980 50596 31036
rect 50596 30980 50600 31036
rect 50536 30976 50600 30980
rect 81016 31036 81080 31040
rect 81016 30980 81020 31036
rect 81020 30980 81076 31036
rect 81076 30980 81080 31036
rect 81016 30976 81080 30980
rect 81096 31036 81160 31040
rect 81096 30980 81100 31036
rect 81100 30980 81156 31036
rect 81156 30980 81160 31036
rect 81096 30976 81160 30980
rect 81176 31036 81240 31040
rect 81176 30980 81180 31036
rect 81180 30980 81236 31036
rect 81236 30980 81240 31036
rect 81176 30976 81240 30980
rect 81256 31036 81320 31040
rect 81256 30980 81260 31036
rect 81260 30980 81316 31036
rect 81316 30980 81320 31036
rect 81256 30976 81320 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 65656 30492 65720 30496
rect 65656 30436 65660 30492
rect 65660 30436 65716 30492
rect 65716 30436 65720 30492
rect 65656 30432 65720 30436
rect 65736 30492 65800 30496
rect 65736 30436 65740 30492
rect 65740 30436 65796 30492
rect 65796 30436 65800 30492
rect 65736 30432 65800 30436
rect 65816 30492 65880 30496
rect 65816 30436 65820 30492
rect 65820 30436 65876 30492
rect 65876 30436 65880 30492
rect 65816 30432 65880 30436
rect 65896 30492 65960 30496
rect 65896 30436 65900 30492
rect 65900 30436 65956 30492
rect 65956 30436 65960 30492
rect 65896 30432 65960 30436
rect 96376 30492 96440 30496
rect 96376 30436 96380 30492
rect 96380 30436 96436 30492
rect 96436 30436 96440 30492
rect 96376 30432 96440 30436
rect 96456 30492 96520 30496
rect 96456 30436 96460 30492
rect 96460 30436 96516 30492
rect 96516 30436 96520 30492
rect 96456 30432 96520 30436
rect 96536 30492 96600 30496
rect 96536 30436 96540 30492
rect 96540 30436 96596 30492
rect 96596 30436 96600 30492
rect 96536 30432 96600 30436
rect 96616 30492 96680 30496
rect 96616 30436 96620 30492
rect 96620 30436 96676 30492
rect 96676 30436 96680 30492
rect 96616 30432 96680 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 50296 29948 50360 29952
rect 50296 29892 50300 29948
rect 50300 29892 50356 29948
rect 50356 29892 50360 29948
rect 50296 29888 50360 29892
rect 50376 29948 50440 29952
rect 50376 29892 50380 29948
rect 50380 29892 50436 29948
rect 50436 29892 50440 29948
rect 50376 29888 50440 29892
rect 50456 29948 50520 29952
rect 50456 29892 50460 29948
rect 50460 29892 50516 29948
rect 50516 29892 50520 29948
rect 50456 29888 50520 29892
rect 50536 29948 50600 29952
rect 50536 29892 50540 29948
rect 50540 29892 50596 29948
rect 50596 29892 50600 29948
rect 50536 29888 50600 29892
rect 81016 29948 81080 29952
rect 81016 29892 81020 29948
rect 81020 29892 81076 29948
rect 81076 29892 81080 29948
rect 81016 29888 81080 29892
rect 81096 29948 81160 29952
rect 81096 29892 81100 29948
rect 81100 29892 81156 29948
rect 81156 29892 81160 29948
rect 81096 29888 81160 29892
rect 81176 29948 81240 29952
rect 81176 29892 81180 29948
rect 81180 29892 81236 29948
rect 81236 29892 81240 29948
rect 81176 29888 81240 29892
rect 81256 29948 81320 29952
rect 81256 29892 81260 29948
rect 81260 29892 81316 29948
rect 81316 29892 81320 29948
rect 81256 29888 81320 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 65656 29404 65720 29408
rect 65656 29348 65660 29404
rect 65660 29348 65716 29404
rect 65716 29348 65720 29404
rect 65656 29344 65720 29348
rect 65736 29404 65800 29408
rect 65736 29348 65740 29404
rect 65740 29348 65796 29404
rect 65796 29348 65800 29404
rect 65736 29344 65800 29348
rect 65816 29404 65880 29408
rect 65816 29348 65820 29404
rect 65820 29348 65876 29404
rect 65876 29348 65880 29404
rect 65816 29344 65880 29348
rect 65896 29404 65960 29408
rect 65896 29348 65900 29404
rect 65900 29348 65956 29404
rect 65956 29348 65960 29404
rect 65896 29344 65960 29348
rect 96376 29404 96440 29408
rect 96376 29348 96380 29404
rect 96380 29348 96436 29404
rect 96436 29348 96440 29404
rect 96376 29344 96440 29348
rect 96456 29404 96520 29408
rect 96456 29348 96460 29404
rect 96460 29348 96516 29404
rect 96516 29348 96520 29404
rect 96456 29344 96520 29348
rect 96536 29404 96600 29408
rect 96536 29348 96540 29404
rect 96540 29348 96596 29404
rect 96596 29348 96600 29404
rect 96536 29344 96600 29348
rect 96616 29404 96680 29408
rect 96616 29348 96620 29404
rect 96620 29348 96676 29404
rect 96676 29348 96680 29404
rect 96616 29344 96680 29348
rect 59124 29064 59188 29068
rect 59124 29008 59174 29064
rect 59174 29008 59188 29064
rect 59124 29004 59188 29008
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 18460 26208 18524 26212
rect 18460 26152 18474 26208
rect 18474 26152 18524 26208
rect 18460 26148 18524 26152
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 82860 25468 82924 25532
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 57468 24924 57532 24988
rect 83596 24924 83660 24988
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 26924 24032 26988 24036
rect 26924 23976 26938 24032
rect 26938 23976 26988 24032
rect 26924 23972 26988 23976
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 56548 23836 56612 23900
rect 82860 23836 82924 23900
rect 12756 23488 12820 23492
rect 12756 23432 12770 23488
rect 12770 23432 12820 23488
rect 12756 23428 12820 23432
rect 14964 23428 15028 23492
rect 18828 23488 18892 23492
rect 18828 23432 18842 23488
rect 18842 23432 18892 23488
rect 18828 23428 18892 23432
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 56916 22884 56980 22948
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 14596 22808 14660 22812
rect 14596 22752 14610 22808
rect 14610 22752 14660 22808
rect 14596 22748 14660 22752
rect 82860 22748 82924 22812
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 82860 21660 82924 21724
rect 25452 21448 25516 21452
rect 25452 21392 25466 21448
rect 25466 21392 25516 21448
rect 25452 21388 25516 21392
rect 57836 21388 57900 21452
rect 14228 21252 14292 21316
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 19196 20708 19260 20772
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 83228 20572 83292 20636
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 15700 20028 15764 20092
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 82860 19484 82924 19548
rect 19196 19408 19260 19412
rect 19196 19352 19210 19408
rect 19210 19352 19260 19408
rect 19196 19348 19260 19352
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 53420 17308 53484 17372
rect 83964 17308 84028 17372
rect 14964 17036 15028 17100
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 13492 16688 13556 16692
rect 13492 16632 13506 16688
rect 13506 16632 13556 16688
rect 13492 16628 13556 16632
rect 20852 16688 20916 16692
rect 20852 16632 20866 16688
rect 20866 16632 20916 16688
rect 20852 16628 20916 16632
rect 82860 16628 82924 16692
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 21404 15948 21468 16012
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 53052 15268 53116 15332
rect 59124 15268 59188 15332
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 59124 13032 59188 13096
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
<< metal4 >>
rect 4208 47904 4528 47920
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43014 4528 43488
rect 4208 42778 4250 43014
rect 4486 42778 4528 43014
rect 4208 42694 4528 42778
rect 4208 42464 4250 42694
rect 4486 42464 4528 42694
rect 4208 42400 4216 42464
rect 4280 42400 4296 42458
rect 4360 42400 4376 42458
rect 4440 42400 4456 42458
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 19568 47360 19888 47920
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 34928 47904 35248 47920
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43014 35248 43488
rect 34928 42778 34970 43014
rect 35206 42778 35248 43014
rect 34928 42694 35248 42778
rect 34928 42464 34970 42694
rect 35206 42464 35248 42694
rect 34928 42400 34936 42464
rect 35000 42400 35016 42458
rect 35080 42400 35096 42458
rect 35160 42400 35176 42458
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29153 35248 29344
rect 50288 47360 50608 47920
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 46272 50608 47296
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 45184 50608 46208
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 44096 50608 45120
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33216 50608 34240
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 32128 50608 33152
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 31040 50608 32064
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 29952 50608 30976
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29153 50608 29888
rect 65648 47904 65968 47920
rect 65648 47840 65656 47904
rect 65720 47840 65736 47904
rect 65800 47840 65816 47904
rect 65880 47840 65896 47904
rect 65960 47840 65968 47904
rect 65648 46816 65968 47840
rect 65648 46752 65656 46816
rect 65720 46752 65736 46816
rect 65800 46752 65816 46816
rect 65880 46752 65896 46816
rect 65960 46752 65968 46816
rect 65648 45728 65968 46752
rect 65648 45664 65656 45728
rect 65720 45664 65736 45728
rect 65800 45664 65816 45728
rect 65880 45664 65896 45728
rect 65960 45664 65968 45728
rect 65648 44640 65968 45664
rect 65648 44576 65656 44640
rect 65720 44576 65736 44640
rect 65800 44576 65816 44640
rect 65880 44576 65896 44640
rect 65960 44576 65968 44640
rect 65648 43552 65968 44576
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43014 65968 43488
rect 65648 42778 65690 43014
rect 65926 42778 65968 43014
rect 65648 42694 65968 42778
rect 65648 42464 65690 42694
rect 65926 42464 65968 42694
rect 65648 42400 65656 42464
rect 65720 42400 65736 42458
rect 65800 42400 65816 42458
rect 65880 42400 65896 42458
rect 65960 42400 65968 42464
rect 65648 41376 65968 42400
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 40288 65968 41312
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 39200 65968 40224
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 38112 65968 39136
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 37024 65968 38048
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 35936 65968 36960
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 34848 65968 35872
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 33760 65968 34784
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 32672 65968 33696
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 31584 65968 32608
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 30496 65968 31520
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 29408 65968 30432
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 29153 65968 29344
rect 81008 47360 81328 47920
rect 81008 47296 81016 47360
rect 81080 47296 81096 47360
rect 81160 47296 81176 47360
rect 81240 47296 81256 47360
rect 81320 47296 81328 47360
rect 81008 46272 81328 47296
rect 81008 46208 81016 46272
rect 81080 46208 81096 46272
rect 81160 46208 81176 46272
rect 81240 46208 81256 46272
rect 81320 46208 81328 46272
rect 81008 45184 81328 46208
rect 81008 45120 81016 45184
rect 81080 45120 81096 45184
rect 81160 45120 81176 45184
rect 81240 45120 81256 45184
rect 81320 45120 81328 45184
rect 81008 44096 81328 45120
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 43008 81328 44032
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 41920 81328 42944
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 40832 81328 41856
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 39744 81328 40768
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 38656 81328 39680
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 37568 81328 38592
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 36480 81328 37504
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 35392 81328 36416
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 34304 81328 35328
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 33216 81328 34240
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 32128 81328 33152
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 31040 81328 32064
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 29952 81328 30976
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 29153 81328 29888
rect 96368 47904 96688 47920
rect 96368 47840 96376 47904
rect 96440 47840 96456 47904
rect 96520 47840 96536 47904
rect 96600 47840 96616 47904
rect 96680 47840 96688 47904
rect 96368 46816 96688 47840
rect 96368 46752 96376 46816
rect 96440 46752 96456 46816
rect 96520 46752 96536 46816
rect 96600 46752 96616 46816
rect 96680 46752 96688 46816
rect 96368 45728 96688 46752
rect 96368 45664 96376 45728
rect 96440 45664 96456 45728
rect 96520 45664 96536 45728
rect 96600 45664 96616 45728
rect 96680 45664 96688 45728
rect 96368 44640 96688 45664
rect 96368 44576 96376 44640
rect 96440 44576 96456 44640
rect 96520 44576 96536 44640
rect 96600 44576 96616 44640
rect 96680 44576 96688 44640
rect 96368 43552 96688 44576
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43014 96688 43488
rect 96368 42778 96410 43014
rect 96646 42778 96688 43014
rect 96368 42694 96688 42778
rect 96368 42464 96410 42694
rect 96646 42464 96688 42694
rect 96368 42400 96376 42464
rect 96440 42400 96456 42458
rect 96520 42400 96536 42458
rect 96600 42400 96616 42458
rect 96680 42400 96688 42464
rect 96368 41376 96688 42400
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 40288 96688 41312
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 39200 96688 40224
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 38112 96688 39136
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 37024 96688 38048
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 35936 96688 36960
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 34848 96688 35872
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 33760 96688 34784
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 32672 96688 33696
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 31584 96688 32608
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 30496 96688 31520
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 29408 96688 30432
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 29153 96688 29344
rect 59123 29068 59189 29069
rect 59123 29004 59124 29068
rect 59188 29004 59189 29068
rect 59123 29003 59189 29004
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25014 19888 25536
rect 19568 24778 19610 25014
rect 19846 24778 19888 25014
rect 57467 24988 57533 24989
rect 57467 24924 57468 24988
rect 57532 24924 57533 24988
rect 57467 24923 57533 24924
rect 19568 24694 19888 24778
rect 19568 24512 19610 24694
rect 19846 24512 19888 24694
rect 19568 24448 19576 24512
rect 19640 24448 19656 24458
rect 19720 24448 19736 24458
rect 19800 24448 19816 24458
rect 19880 24448 19888 24512
rect 12755 23492 12821 23493
rect 12755 23428 12756 23492
rect 12820 23428 12821 23492
rect 12755 23427 12821 23428
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 12758 22218 12818 23427
rect 18827 23492 18893 23493
rect 18827 23428 18828 23492
rect 18892 23428 18893 23492
rect 18827 23427 18893 23428
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 14227 21316 14293 21317
rect 14227 21252 14228 21316
rect 14292 21252 14293 21316
rect 14227 21251 14293 21252
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 14230 14738 14290 21251
rect 18830 18818 18890 23427
rect 19568 23424 19888 24448
rect 26923 24036 26989 24037
rect 26923 23972 26924 24036
rect 26988 23972 26989 24036
rect 26923 23971 26989 23972
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 26926 18138 26986 23971
rect 56547 23900 56613 23901
rect 56547 23836 56548 23900
rect 56612 23836 56613 23900
rect 56547 23835 56613 23836
rect 56550 22218 56610 23835
rect 56915 22948 56981 22949
rect 56915 22884 56916 22948
rect 56980 22884 56981 22948
rect 56915 22883 56981 22884
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 14963 17100 15029 17101
rect 14963 17036 14964 17100
rect 15028 17036 15029 17100
rect 14963 17035 15029 17036
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 14966 12018 15026 17035
rect 19568 16896 19888 17920
rect 53419 17372 53485 17373
rect 53419 17308 53420 17372
rect 53484 17308 53485 17372
rect 53419 17307 53485 17308
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 20851 16692 20917 16693
rect 20851 16628 20852 16692
rect 20916 16628 20917 16692
rect 20851 16627 20917 16628
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 20854 13378 20914 16627
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7014 4528 7584
rect 4208 6778 4250 7014
rect 4486 6778 4528 7014
rect 4208 6694 4528 6778
rect 4208 6560 4250 6694
rect 4486 6560 4528 6694
rect 4208 6496 4216 6560
rect 4520 6496 4528 6560
rect 4208 6458 4250 6496
rect 4486 6458 4528 6496
rect 4208 5472 4528 6458
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 33734 11250 33794 15862
rect 34470 14738 34530 15862
rect 53051 15332 53117 15333
rect 53051 15268 53052 15332
rect 53116 15268 53117 15332
rect 53051 15267 53117 15268
rect 53054 14058 53114 15267
rect 53422 13378 53482 17307
rect 56918 14738 56978 22883
rect 57470 18138 57530 24923
rect 59126 15333 59186 29003
rect 82862 25533 82922 26062
rect 82859 25532 82925 25533
rect 82859 25468 82860 25532
rect 82924 25468 82925 25532
rect 82859 25467 82925 25468
rect 83595 24988 83661 24989
rect 83595 24924 83596 24988
rect 83660 24924 83661 24988
rect 83595 24923 83661 24924
rect 82859 23900 82925 23901
rect 82859 23836 82860 23900
rect 82924 23836 82925 23900
rect 82859 23835 82925 23836
rect 82862 23578 82922 23835
rect 82859 21724 82925 21725
rect 82859 21660 82860 21724
rect 82924 21660 82925 21724
rect 82859 21659 82925 21660
rect 82862 20858 82922 21659
rect 83227 20636 83293 20637
rect 83227 20572 83228 20636
rect 83292 20572 83293 20636
rect 83227 20571 83293 20572
rect 82862 19549 82922 19942
rect 82859 19548 82925 19549
rect 82859 19484 82860 19548
rect 82924 19484 82925 19548
rect 83230 19498 83290 20571
rect 82859 19483 82925 19484
rect 83598 18818 83658 24923
rect 83963 17372 84029 17373
rect 83963 17308 83964 17372
rect 84028 17308 84029 17372
rect 83963 17307 84029 17308
rect 59123 15332 59189 15333
rect 59123 15268 59124 15332
rect 59188 15268 59189 15332
rect 59123 15267 59189 15268
rect 34102 11250 34162 11782
rect 35390 11338 35450 13142
rect 59126 13097 59186 15267
rect 59123 13096 59189 13097
rect 59123 13032 59124 13096
rect 59188 13032 59189 13096
rect 59123 13031 59189 13032
rect 83966 12018 84026 17307
rect 33734 11190 34162 11250
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
<< via4 >>
rect 4250 42778 4486 43014
rect 4250 42464 4486 42694
rect 4250 42458 4280 42464
rect 4280 42458 4296 42464
rect 4296 42458 4360 42464
rect 4360 42458 4376 42464
rect 4376 42458 4440 42464
rect 4440 42458 4456 42464
rect 4456 42458 4486 42464
rect 34970 42778 35206 43014
rect 34970 42464 35206 42694
rect 34970 42458 35000 42464
rect 35000 42458 35016 42464
rect 35016 42458 35080 42464
rect 35080 42458 35096 42464
rect 35096 42458 35160 42464
rect 35160 42458 35176 42464
rect 35176 42458 35206 42464
rect 65690 42778 65926 43014
rect 65690 42464 65926 42694
rect 65690 42458 65720 42464
rect 65720 42458 65736 42464
rect 65736 42458 65800 42464
rect 65800 42458 65816 42464
rect 65816 42458 65880 42464
rect 65880 42458 65896 42464
rect 65896 42458 65926 42464
rect 96410 42778 96646 43014
rect 96410 42464 96646 42694
rect 96410 42458 96440 42464
rect 96440 42458 96456 42464
rect 96456 42458 96520 42464
rect 96520 42458 96536 42464
rect 96536 42458 96600 42464
rect 96600 42458 96616 42464
rect 96616 42458 96646 42464
rect 18374 26212 18610 26298
rect 18374 26148 18460 26212
rect 18460 26148 18524 26212
rect 18524 26148 18610 26212
rect 18374 26062 18610 26148
rect 19610 24778 19846 25014
rect 19610 24512 19846 24694
rect 19610 24458 19640 24512
rect 19640 24458 19656 24512
rect 19656 24458 19720 24512
rect 19720 24458 19736 24512
rect 19736 24458 19800 24512
rect 19800 24458 19816 24512
rect 19816 24458 19846 24512
rect 14878 23492 15114 23578
rect 14878 23428 14964 23492
rect 14964 23428 15028 23492
rect 15028 23428 15114 23492
rect 14878 23342 15114 23428
rect 14510 22812 14746 22898
rect 14510 22748 14596 22812
rect 14596 22748 14660 22812
rect 14660 22748 14746 22812
rect 14510 22662 14746 22748
rect 12670 21982 12906 22218
rect 13406 16692 13642 16778
rect 13406 16628 13492 16692
rect 13492 16628 13556 16692
rect 13556 16628 13642 16692
rect 13406 16542 13642 16628
rect 15614 20092 15850 20178
rect 15614 20028 15700 20092
rect 15700 20028 15764 20092
rect 15764 20028 15850 20092
rect 15614 19942 15850 20028
rect 25366 21452 25602 21538
rect 25366 21388 25452 21452
rect 25452 21388 25516 21452
rect 25516 21388 25602 21452
rect 25366 21302 25602 21388
rect 19110 20772 19346 20858
rect 19110 20708 19196 20772
rect 19196 20708 19260 20772
rect 19260 20708 19346 20772
rect 19110 20622 19346 20708
rect 19110 19412 19346 19498
rect 19110 19348 19196 19412
rect 19196 19348 19260 19412
rect 19260 19348 19346 19412
rect 19110 19262 19346 19348
rect 18742 18582 18978 18818
rect 56462 21982 56698 22218
rect 14142 14502 14378 14738
rect 26838 17902 27074 18138
rect 21318 16012 21554 16098
rect 21318 15948 21404 16012
rect 21404 15948 21468 16012
rect 21468 15948 21554 16012
rect 21318 15862 21554 15948
rect 33646 15862 33882 16098
rect 34382 15862 34618 16098
rect 20766 13142 21002 13378
rect 14878 11782 15114 12018
rect 4250 6778 4486 7014
rect 4250 6560 4486 6694
rect 4250 6496 4280 6560
rect 4280 6496 4296 6560
rect 4296 6496 4360 6560
rect 4360 6496 4376 6560
rect 4376 6496 4440 6560
rect 4440 6496 4456 6560
rect 4456 6496 4486 6560
rect 4250 6458 4486 6496
rect 34382 14502 34618 14738
rect 52966 13822 53202 14058
rect 57750 21452 57986 21538
rect 57750 21388 57836 21452
rect 57836 21388 57900 21452
rect 57900 21388 57986 21452
rect 57750 21302 57986 21388
rect 57382 17902 57618 18138
rect 82774 26062 83010 26298
rect 82774 23342 83010 23578
rect 82774 22812 83010 22898
rect 82774 22748 82860 22812
rect 82860 22748 82924 22812
rect 82924 22748 83010 22812
rect 82774 22662 83010 22748
rect 82774 20622 83010 20858
rect 82774 19942 83010 20178
rect 83142 19262 83378 19498
rect 83510 18582 83746 18818
rect 82774 16692 83010 16778
rect 82774 16628 82860 16692
rect 82860 16628 82924 16692
rect 82924 16628 83010 16692
rect 82774 16542 83010 16628
rect 56830 14502 57066 14738
rect 35302 13142 35538 13378
rect 53334 13142 53570 13378
rect 34014 11782 34250 12018
rect 83878 11782 84114 12018
rect 35302 11102 35538 11338
<< metal5 >>
rect 4208 43036 4528 43038
rect 34928 43036 35248 43038
rect 65648 43036 65968 43038
rect 96368 43036 96688 43038
rect 1104 43014 108008 43036
rect 1104 42778 4250 43014
rect 4486 42778 34970 43014
rect 35206 42778 65690 43014
rect 65926 42778 96410 43014
rect 96646 42778 108008 43014
rect 1104 42694 108008 42778
rect 1104 42458 4250 42694
rect 4486 42458 34970 42694
rect 35206 42458 65690 42694
rect 65926 42458 96410 42694
rect 96646 42458 108008 42694
rect 1104 42436 108008 42458
rect 4208 42434 4528 42436
rect 34928 42434 35248 42436
rect 65648 42434 65968 42436
rect 96368 42434 96688 42436
rect 18332 26298 83052 26340
rect 18332 26062 18374 26298
rect 18610 26062 82774 26298
rect 83010 26062 83052 26298
rect 18332 26020 83052 26062
rect 19568 25036 19888 25038
rect 1104 25014 108008 25036
rect 1104 24778 19610 25014
rect 19846 24778 108008 25014
rect 1104 24694 108008 24778
rect 1104 24458 19610 24694
rect 19846 24458 108008 24694
rect 1104 24436 108008 24458
rect 19568 24434 19888 24436
rect 14836 23578 83052 23620
rect 14836 23342 14878 23578
rect 15114 23342 82774 23578
rect 83010 23342 83052 23578
rect 14836 23300 83052 23342
rect 14468 22898 83052 22940
rect 14468 22662 14510 22898
rect 14746 22662 82774 22898
rect 83010 22662 83052 22898
rect 14468 22620 83052 22662
rect 12628 22218 56740 22260
rect 12628 21982 12670 22218
rect 12906 21982 56462 22218
rect 56698 21982 56740 22218
rect 12628 21940 56740 21982
rect 25324 21538 58028 21580
rect 25324 21302 25366 21538
rect 25602 21302 57750 21538
rect 57986 21302 58028 21538
rect 25324 21260 58028 21302
rect 19068 20858 83052 20900
rect 19068 20622 19110 20858
rect 19346 20622 82774 20858
rect 83010 20622 83052 20858
rect 19068 20580 83052 20622
rect 15572 20178 83052 20220
rect 15572 19942 15614 20178
rect 15850 19942 82774 20178
rect 83010 19942 83052 20178
rect 15572 19900 83052 19942
rect 19068 19498 83420 19540
rect 19068 19262 19110 19498
rect 19346 19262 83142 19498
rect 83378 19262 83420 19498
rect 19068 19220 83420 19262
rect 18700 18818 83788 18860
rect 18700 18582 18742 18818
rect 18978 18582 83510 18818
rect 83746 18582 83788 18818
rect 18700 18540 83788 18582
rect 26796 18138 57660 18180
rect 26796 17902 26838 18138
rect 27074 17902 57382 18138
rect 57618 17902 57660 18138
rect 26796 17860 57660 17902
rect 13364 16778 83052 16820
rect 13364 16542 13406 16778
rect 13642 16542 82774 16778
rect 83010 16542 83052 16778
rect 13364 16500 83052 16542
rect 21276 16098 33924 16140
rect 21276 15862 21318 16098
rect 21554 15862 33646 16098
rect 33882 15862 33924 16098
rect 21276 15820 33924 15862
rect 34340 16098 38524 16140
rect 34340 15862 34382 16098
rect 34618 15862 38524 16098
rect 34340 15820 38524 15862
rect 38204 14780 38524 15820
rect 14100 14738 34660 14780
rect 14100 14502 14142 14738
rect 14378 14502 34382 14738
rect 34618 14502 34660 14738
rect 14100 14460 34660 14502
rect 38204 14738 57108 14780
rect 38204 14502 56830 14738
rect 57066 14502 57108 14738
rect 38204 14460 57108 14502
rect 38204 14058 53244 14100
rect 38204 13822 52966 14058
rect 53202 13822 53244 14058
rect 38204 13780 53244 13822
rect 38204 13420 38524 13780
rect 20724 13378 35580 13420
rect 20724 13142 20766 13378
rect 21002 13142 35302 13378
rect 35538 13142 35580 13378
rect 20724 13100 35580 13142
rect 38020 13100 38524 13420
rect 39124 13378 53612 13420
rect 39124 13142 53334 13378
rect 53570 13142 53612 13378
rect 39124 13100 53612 13142
rect 38020 12060 38340 13100
rect 39124 12740 39444 13100
rect 14836 12018 33372 12060
rect 14836 11782 14878 12018
rect 15114 11782 33372 12018
rect 14836 11740 33372 11782
rect 33972 12018 38340 12060
rect 33972 11782 34014 12018
rect 34250 11782 38340 12018
rect 33972 11740 38340 11782
rect 38756 12420 39444 12740
rect 33052 10020 33372 11740
rect 38756 11380 39076 12420
rect 35260 11338 39076 11380
rect 35260 11102 35302 11338
rect 35538 11102 39076 11338
rect 35260 11060 39076 11102
rect 39492 12018 84156 12060
rect 39492 11782 83878 12018
rect 84114 11782 84156 12018
rect 39492 11740 84156 11782
rect 39492 10020 39812 11740
rect 33052 9700 39812 10020
rect 4208 7036 4528 7038
rect 1104 7014 108008 7036
rect 1104 6778 4250 7014
rect 4486 6778 108008 7014
rect 1104 6694 108008 6778
rect 1104 6458 4250 6694
rect 4486 6458 108008 6694
rect 1104 6436 108008 6458
rect 4208 6434 4528 6436
use sky130_fd_sc_hd__fill_1  FILLER_1_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2852 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607194113
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607194113
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607194113
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607194113
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1607194113
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__D $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1483_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2944 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1607194113
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1607194113
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607194113
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__CLK
timestamp 1607194113
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1607194113
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607194113
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1607194113
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607194113
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1607194113
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607194113
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1607194113
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1607194113
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607194113
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1607194113
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607194113
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1607194113
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607194113
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607194113
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1607194113
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1607194113
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1607194113
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607194113
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1607194113
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607194113
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1607194113
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1607194113
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1607194113
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607194113
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607194113
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607194113
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1607194113
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1607194113
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1607194113
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1607194113
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1607194113
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1607194113
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607194113
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1607194113
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1607194113
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1607194113
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1607194113
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607194113
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1607194113
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1607194113
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1607194113
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607194113
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607194113
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607194113
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607194113
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607194113
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607194113
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607194113
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607194113
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607194113
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607194113
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1607194113
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607194113
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1607194113
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607194113
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1607194113
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607194113
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1607194113
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607194113
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1607194113
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1607194113
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1607194113
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1607194113
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1607194113
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607194113
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1607194113
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1607194113
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607194113
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607194113
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1484_
timestamp 1607194113
transform 1 0 3588 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1607194113
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5704 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__CLK
timestamp 1607194113
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__D
timestamp 1607194113
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1607194113
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1607194113
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607194113
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1607194113
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1607194113
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1607194113
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1607194113
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1607194113
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607194113
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1607194113
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1607194113
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1607194113
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1607194113
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1607194113
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607194113
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1607194113
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1607194113
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1607194113
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607194113
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607194113
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607194113
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607194113
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607194113
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607194113
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1607194113
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1607194113
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1607194113
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1607194113
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607194113
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1485_
timestamp 1607194113
transform 1 0 9660 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_114
timestamp 1607194113
transform 1 0 11592 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__CLK
timestamp 1607194113
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_138
timestamp 1607194113
transform 1 0 13800 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_126
timestamp 1607194113
transform 1 0 12696 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1607194113
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1607194113
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607194113
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1607194113
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1607194113
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1607194113
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607194113
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1607194113
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607194113
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1607194113
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1607194113
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607194113
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607194113
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1607194113
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1607194113
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1607194113
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1607194113
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1607194113
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607194113
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1607194113
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1607194113
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1607194113
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1607194113
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1607194113
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607194113
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1607194113
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1607194113
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1607194113
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1607194113
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607194113
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607194113
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1607194113
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1607194113
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1607194113
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp 1607194113
transform 1 0 2484 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607194113
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607194113
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607194113
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607194113
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607194113
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_21
timestamp 1607194113
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1607194113
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607194113
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607194113
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1486_
timestamp 1607194113
transform 1 0 3128 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_7_55
timestamp 1607194113
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1607194113
transform 1 0 5060 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1607194113
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1607194113
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__CLK
timestamp 1607194113
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1607194113
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1607194113
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1607194113
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607194113
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1607194113
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1607194113
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1607194113
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1607194113
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607194113
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1607194113
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1607194113
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1607194113
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1607194113
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1607194113
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1607194113
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607194113
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1607194113
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1607194113
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1607194113
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607194113
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1607194113
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1607194113
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1607194113
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1607194113
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1607194113
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1607194113
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1607194113
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607194113
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1607194113
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1607194113
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1607194113
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607194113
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1607194113
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1607194113
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1607194113
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607194113
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607194113
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607194113
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607194113
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607194113
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607194113
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1607194113
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1607194113
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1607194113
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1607194113
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:5.inst.g_clkdly15_2.dly $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1607194113
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1607194113
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607194113
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1607194113
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1607194113
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__CLK
timestamp 1607194113
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1343_
timestamp 1607194113
transform 1 0 12236 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1607194113
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1607194113
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_140
timestamp 1607194113
transform 1 0 13984 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607194113
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1607194113
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1607194113
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1607194113
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1607194113
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1607194113
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607194113
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1607194113
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1607194113
transform 1 0 2484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607194113
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607194113
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1487_
timestamp 1607194113
transform 1 0 2576 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_37
timestamp 1607194113
transform 1 0 4508 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__CLK
timestamp 1607194113
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_49
timestamp 1607194113
transform 1 0 5612 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_70
timestamp 1607194113
transform 1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1607194113
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607194113
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1342_
timestamp 1607194113
transform 1 0 7820 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1607194113
transform 1 0 9752 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__CLK
timestamp 1607194113
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1607194113
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp 1607194113
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:6.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_131
timestamp 1607194113
transform 1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1607194113
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__CLK
timestamp 1607194113
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607194113
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1335_
timestamp 1607194113
transform 1 0 13616 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_155
timestamp 1607194113
transform 1 0 15364 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_167
timestamp 1607194113
transform 1 0 16468 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1607194113
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1607194113
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1607194113
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607194113
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1607194113
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1607194113
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1607194113
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607194113
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607194113
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607194113
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607194113
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607194113
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1341_
timestamp 1607194113
transform 1 0 4048 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1607194113
transform 1 0 5980 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1607194113
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1607194113
transform 1 0 7084 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:4.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1607194113
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1607194113
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607194113
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1607194113
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1607194113
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1607194113
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1607194113
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1607194113
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607194113
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1607194113
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1607194113
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1607194113
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1607194113
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1607194113
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607194113
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1607194113
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1607194113
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607194113
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607194113
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1607194113
transform 1 0 2576 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1607194113
transform 1 0 4508 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__CLK
timestamp 1607194113
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_49
timestamp 1607194113
transform 1 0 5612 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1607194113
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1607194113
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607194113
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__CLK
timestamp 1607194113
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1334_
timestamp 1607194113
transform 1 0 8464 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1607194113
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_101
timestamp 1607194113
transform 1 0 10396 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1607194113
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1607194113
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1607194113
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607194113
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1340_
timestamp 1607194113
transform 1 0 12788 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_158
timestamp 1607194113
transform 1 0 15640 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_146
timestamp 1607194113
transform 1 0 14536 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_170
timestamp 1607194113
transform 1 0 16744 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1607194113
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1607194113
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1607194113
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607194113
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_208
timestamp 1607194113
transform 1 0 20240 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:3.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 20792 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_223
timestamp 1607194113
transform 1 0 21620 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607194113
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607194113
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607194113
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1607194113
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607194113
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607194113
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1607194113
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1333_
timestamp 1607194113
transform 1 0 4968 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_12_75
timestamp 1607194113
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_63
timestamp 1607194113
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__CLK
timestamp 1607194113
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1607194113
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1607194113
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1607194113
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607194113
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1607194113
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1607194113
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1607194113
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1607194113
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1607194113
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607194113
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_178
timestamp 1607194113
transform 1 0 17480 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1607194113
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1444_
timestamp 1607194113
transform 1 0 17756 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1607194113
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1607194113
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1607194113
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607194113
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_223
timestamp 1607194113
transform 1 0 21620 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1339_
timestamp 1607194113
transform 1 0 21896 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607194113
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607194113
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1607194113
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607194113
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607194113
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607194113
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607194113
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607194113
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1607194113
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1607194113
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607194113
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1607194113
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1607194113
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1607194113
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1607194113
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1607194113
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_76
timestamp 1607194113
transform 1 0 8096 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607194113
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6808 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _1164_
timestamp 1607194113
transform 1 0 7544 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1607194113
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1607194113
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_88
timestamp 1607194113
transform 1 0 9200 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607194113
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_117
timestamp 1607194113
transform 1 0 11868 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1607194113
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1607194113
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_100
timestamp 1607194113
transform 1 0 10304 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_123
timestamp 1607194113
transform 1 0 12420 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1607194113
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1607194113
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1607194113
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607194113
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1445_
timestamp 1607194113
transform 1 0 12696 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1332_
timestamp 1607194113
transform 1 0 13708 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1607194113
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1607194113
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1607194113
transform 1 0 15640 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__CLK
timestamp 1607194113
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607194113
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1607194113
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1607194113
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_170
timestamp 1607194113
transform 1 0 16744 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1607194113
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1607194113
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B2
timestamp 1607194113
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607194113
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1167_
timestamp 1607194113
transform 1 0 18032 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_14_211
timestamp 1607194113
transform 1 0 20516 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1607194113
transform 1 0 19964 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_218
timestamp 1607194113
transform 1 0 21160 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_212
timestamp 1607194113
transform 1 0 20608 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_200
timestamp 1607194113
transform 1 0 19504 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 19688 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607194113
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1338_
timestamp 1607194113
transform 1 0 20884 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_13_228
timestamp 1607194113
transform 1 0 22080 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:2.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 21252 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1607194113
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607194113
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607194113
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1489_
timestamp 1607194113
transform 1 0 2576 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1607194113
transform 1 0 4508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__CLK
timestamp 1607194113
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_49
timestamp 1607194113
transform 1 0 5612 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1607194113
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607194113
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1447_
timestamp 1607194113
transform 1 0 7360 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_89
timestamp 1607194113
transform 1 0 9292 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1607194113
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1607194113
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_101
timestamp 1607194113
transform 1 0 10396 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1607194113
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1607194113
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607194113
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1166_
timestamp 1607194113
transform 1 0 13524 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1607194113
transform 1 0 14812 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_173
timestamp 1607194113
transform 1 0 17020 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_161
timestamp 1607194113
transform 1 0 15916 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1607194113
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1607194113
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1607194113
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607194113
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1607194113
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__CLK
timestamp 1607194113
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1330_
timestamp 1607194113
transform 1 0 20608 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_231
timestamp 1607194113
transform 1 0 22356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607194113
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607194113
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607194113
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607194113
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607194113
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607194113
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_48
timestamp 1607194113
transform 1 0 5520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_44
timestamp 1607194113
transform 1 0 5152 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1446_
timestamp 1607194113
transform 1 0 5612 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_70
timestamp 1607194113
transform 1 0 7544 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__CLK
timestamp 1607194113
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1607194113
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1607194113
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_82
timestamp 1607194113
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607194113
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1607194113
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1607194113
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1607194113
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1162_
timestamp 1607194113
transform 1 0 13156 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_16_154
timestamp 1607194113
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_147
timestamp 1607194113
transform 1 0 14628 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A2
timestamp 1607194113
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607194113
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_167
timestamp 1607194113
transform 1 0 16468 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_160
timestamp 1607194113
transform 1 0 15824 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1607194113
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15916 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_191
timestamp 1607194113
transform 1 0 18676 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_179
timestamp 1607194113
transform 1 0 17572 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1607194113
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1607194113
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_203
timestamp 1607194113
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607194113
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1607194113
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1607194113
transform 1 0 2484 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607194113
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607194113
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1490_
timestamp 1607194113
transform 1 0 2576 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1607194113
transform 1 0 4508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__CLK
timestamp 1607194113
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1607194113
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_74
timestamp 1607194113
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1607194113
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607194113
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8188 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_96
timestamp 1607194113
transform 1 0 9936 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_84
timestamp 1607194113
transform 1 0 8832 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_108
timestamp 1607194113
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1607194113
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607194113
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1448_
timestamp 1607194113
transform 1 0 12420 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1607194113
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1607194113
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__CLK
timestamp 1607194113
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1607194113
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_168
timestamp 1607194113
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1161_
timestamp 1607194113
transform 1 0 16836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__B2
timestamp 1607194113
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607194113
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1168_
timestamp 1607194113
transform 1 0 18032 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_17_212
timestamp 1607194113
transform 1 0 20608 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_200
timestamp 1607194113
transform 1 0 19504 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:1.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 20976 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1607194113
transform 1 0 21804 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607194113
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607194113
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607194113
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607194113
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607194113
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607194113
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_56
timestamp 1607194113
transform 1 0 6256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1607194113
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_71
timestamp 1607194113
transform 1 0 7636 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0976_
timestamp 1607194113
transform 1 0 6992 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1607194113
transform 1 0 10212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1607194113
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1607194113
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1607194113
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607194113
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_107
timestamp 1607194113
transform 1 0 10948 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0983_
timestamp 1607194113
transform 1 0 10304 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0960_
timestamp 1607194113
transform 1 0 11684 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_134
timestamp 1607194113
transform 1 0 13432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_122
timestamp 1607194113
transform 1 0 12328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1607194113
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1607194113
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_146
timestamp 1607194113
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607194113
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_174
timestamp 1607194113
transform 1 0 17112 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_166
timestamp 1607194113
transform 1 0 16376 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1443_
timestamp 1607194113
transform 1 0 17204 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_196
timestamp 1607194113
transform 1 0 19136 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1607194113
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1607194113
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_208
timestamp 1607194113
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607194113
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_233
timestamp 1607194113
transform 1 0 22540 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_227
timestamp 1607194113
transform 1 0 21988 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607194113
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607194113
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp 1607194113
transform 1 0 2484 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607194113
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607194113
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607194113
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1491_
timestamp 1607194113
transform 1 0 2576 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607194113
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607194113
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1607194113
transform 1 0 4508 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__CLK
timestamp 1607194113
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607194113
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1607194113
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1607194113
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_49
timestamp 1607194113
transform 1 0 5612 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1607194113
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_71
timestamp 1607194113
transform 1 0 7636 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_74
timestamp 1607194113
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1607194113
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1607194113
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607194113
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8188 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6624 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0975_
timestamp 1607194113
transform 1 0 8188 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1607194113
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_86
timestamp 1607194113
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_88
timestamp 1607194113
transform 1 0 9200 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B
timestamp 1607194113
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__C
timestamp 1607194113
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607194113
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1002_
timestamp 1607194113
transform 1 0 9752 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_20_115
timestamp 1607194113
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_103
timestamp 1607194113
transform 1 0 10580 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1607194113
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1607194113
transform 1 0 10304 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B
timestamp 1607194113
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0968_
timestamp 1607194113
transform 1 0 10396 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1607194113
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1607194113
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1607194113
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607194113
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1607194113
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1607194113
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1607194113
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1607194113
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A
timestamp 1607194113
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607194113
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1607194113
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_166
timestamp 1607194113
transform 1 0 16376 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_172
timestamp 1607194113
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_160
timestamp 1607194113
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1169_
timestamp 1607194113
transform 1 0 17020 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_20_189
timestamp 1607194113
transform 1 0 18492 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1607194113
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1607194113
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1607194113
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B1
timestamp 1607194113
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607194113
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1607194113
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1607194113
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1607194113
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1607194113
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607194113
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1607194113
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1607194113
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1329_
timestamp 1607194113
transform 1 0 21620 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1607194113
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607194113
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607194113
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1492_
timestamp 1607194113
transform 1 0 2576 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1607194113
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__CLK
timestamp 1607194113
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__D
timestamp 1607194113
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1607194113
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1607194113
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_72
timestamp 1607194113
transform 1 0 7728 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1607194113
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1607194113
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A
timestamp 1607194113
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607194113
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1607194113
transform 1 0 7360 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_91
timestamp 1607194113
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__C
timestamp 1607194113
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0990_
timestamp 1607194113
transform 1 0 8464 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1607194113
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_106
timestamp 1607194113
transform 1 0 10856 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk_i
timestamp 1607194113
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_128
timestamp 1607194113
transform 1 0 12880 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1607194113
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607194113
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1607194113
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_156
timestamp 1607194113
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B1
timestamp 1607194113
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1170_
timestamp 1607194113
transform 1 0 13984 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_21_168
timestamp 1607194113
transform 1 0 16560 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1607194113
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1607194113
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1607194113
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607194113
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1607194113
transform 1 0 20608 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1607194113
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__CLK
timestamp 1607194113
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1337_
timestamp 1607194113
transform 1 0 20884 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607194113
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607194113
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607194113
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607194113
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607194113
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607194113
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1607194113
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1607194113
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_76
timestamp 1607194113
transform 1 0 8096 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_68
timestamp 1607194113
transform 1 0 7360 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0956_
timestamp 1607194113
transform 1 0 8188 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1607194113
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1607194113
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607194113
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_117
timestamp 1607194113
transform 1 0 11868 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1607194113
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1607194113
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1441_
timestamp 1607194113
transform 1 0 12696 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1607194113
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1607194113
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607194113
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1442_
timestamp 1607194113
transform 1 0 16376 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_187
timestamp 1607194113
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__CLK
timestamp 1607194113
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1607194113
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1607194113
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607194113
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_226
timestamp 1607194113
transform 1 0 21896 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly_A
timestamp 1607194113
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 1607194113
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607194113
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607194113
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1493_
timestamp 1607194113
transform 1 0 2668 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__CLK
timestamp 1607194113
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__D
timestamp 1607194113
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_52
timestamp 1607194113
transform 1 0 5888 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1607194113
transform 1 0 4784 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1607194113
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1607194113
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1607194113
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607194113
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1607194113
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1607194113
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1607194113
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1607194113
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1607194113
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__CLK
timestamp 1607194113
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607194113
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1328_
timestamp 1607194113
transform 1 0 13524 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1607194113
transform 1 0 15272 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1607194113
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_166
timestamp 1607194113
transform 1 0 16376 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1607194113
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1607194113
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1607194113
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607194113
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1607194113
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1607194113
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1607194113
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607194113
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607194113
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607194113
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1607194113
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607194113
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607194113
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1607194113
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__B1
timestamp 1607194113
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6440 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1607194113
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1607194113
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1607194113
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607194113
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1607194113
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1607194113
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1607194113
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1607194113
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1607194113
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607194113
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1607194113
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1607194113
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1607194113
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1607194113
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1607194113
transform 1 0 21160 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607194113
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1607194113
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_232
timestamp 1607194113
transform 1 0 22448 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_220
timestamp 1607194113
transform 1 0 21344 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1607194113
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607194113
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607194113
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1494_
timestamp 1607194113
transform 1 0 2576 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1607194113
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__CLK
timestamp 1607194113
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__D
timestamp 1607194113
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607194113
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1607194113
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1607194113
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607194113
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1367_
timestamp 1607194113
transform 1 0 7176 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_96
timestamp 1607194113
transform 1 0 9936 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1607194113
transform 1 0 9108 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__CLK
timestamp 1607194113
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A
timestamp 1607194113
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1281_
timestamp 1607194113
transform 1 0 9660 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_108
timestamp 1607194113
transform 1 0 11040 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1607194113
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1607194113
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__CLK
timestamp 1607194113
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607194113
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1336_
timestamp 1607194113
transform 1 0 12972 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_150
timestamp 1607194113
transform 1 0 14904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__D
timestamp 1607194113
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1607194113
transform 1 0 17112 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_162
timestamp 1607194113
transform 1 0 16008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1607194113
transform 1 0 19136 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1607194113
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1607194113
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607194113
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1607194113
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1408_
timestamp 1607194113
transform 1 0 19596 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_222
timestamp 1607194113
transform 1 0 21528 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__CLK
timestamp 1607194113
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_15
timestamp 1607194113
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607194113
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607194113
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607194113
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607194113
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607194113
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1495_
timestamp 1607194113
transform 1 0 2576 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1607194113
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607194113
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607194113
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__CLK
timestamp 1607194113
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__D
timestamp 1607194113
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607194113
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1607194113
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1607194113
transform 1 0 6256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607194113
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B1
timestamp 1607194113
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_78
timestamp 1607194113
transform 1 0 8280 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607194113
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1366_
timestamp 1607194113
transform 1 0 6992 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1287_
timestamp 1607194113
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1607194113
transform 1 0 9384 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1607194113
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1607194113
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1607194113
transform 1 0 8924 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__CLK
timestamp 1607194113
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607194113
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1607194113
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1607194113
transform 1 0 10488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1607194113
transform 1 0 11868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1607194113
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_123
timestamp 1607194113
transform 1 0 12420 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_137
timestamp 1607194113
transform 1 0 13708 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1607194113
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1607194113
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_i
timestamp 1607194113
transform 1 0 13156 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607194113
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0967_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13432 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_4  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12420 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1607194113
transform 1 0 15364 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1607194113
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1607194113
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__C1
timestamp 1607194113
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B1
timestamp 1607194113
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607194113
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_167
timestamp 1607194113
transform 1 0 16468 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_178
timestamp 1607194113
transform 1 0 17480 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1607194113
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1607194113
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1607194113
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1607194113
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B1
timestamp 1607194113
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607194113
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1407_
timestamp 1607194113
transform 1 0 19136 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1222_
timestamp 1607194113
transform 1 0 18584 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_217
timestamp 1607194113
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1607194113
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1607194113
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__CLK
timestamp 1607194113
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A2_N
timestamp 1607194113
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B2
timestamp 1607194113
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607194113
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1607194113
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1607194113
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1607194113
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607194113
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607194113
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1607194113
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1607194113
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607194113
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1607194113
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1607194113
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_78
timestamp 1607194113
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1607194113
transform 1 0 7728 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1607194113
transform 1 0 7360 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1607194113
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1607194113
transform 1 0 7820 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1607194113
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1607194113
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607194113
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1607194113
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1607194113
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1607194113
transform 1 0 13616 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_133
timestamp 1607194113
transform 1 0 13340 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1607194113
transform 1 0 12972 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_i_A
timestamp 1607194113
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1607194113
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1607194113
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_144
timestamp 1607194113
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_140
timestamp 1607194113
transform 1 0 13984 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607194113
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1607194113
transform 1 0 14076 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_178
timestamp 1607194113
transform 1 0 17480 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1607194113
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_186
timestamp 1607194113
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B1
timestamp 1607194113
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1223_
timestamp 1607194113
transform 1 0 18492 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1607194113
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1607194113
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1607194113
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A2_N
timestamp 1607194113
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B2
timestamp 1607194113
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607194113
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1607194113
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_232
timestamp 1607194113
transform 1 0 22448 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_220
timestamp 1607194113
transform 1 0 21344 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1607194113
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1607194113
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607194113
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1496_
timestamp 1607194113
transform 1 0 2576 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1607194113
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__CLK
timestamp 1607194113
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__D
timestamp 1607194113
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1607194113
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1607194113
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1607194113
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1607194113
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607194113
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_96
timestamp 1607194113
transform 1 0 9936 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_92
timestamp 1607194113
transform 1 0 9568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_86
timestamp 1607194113
transform 1 0 9016 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk_i
timestamp 1607194113
transform 1 0 9660 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_108
timestamp 1607194113
transform 1 0 11040 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_135
timestamp 1607194113
transform 1 0 13524 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1607194113
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1607194113
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607194113
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_157
timestamp 1607194113
transform 1 0 15548 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_145
timestamp 1607194113
transform 1 0 14444 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_141
timestamp 1607194113
transform 1 0 14076 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1607194113
transform 1 0 14168 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1607194113
transform 1 0 16652 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_190
timestamp 1607194113
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1607194113
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1607194113
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607194113
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0953_
timestamp 1607194113
transform 1 0 18676 0 1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_29_209
timestamp 1607194113
transform 1 0 20332 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B2
timestamp 1607194113
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B1
timestamp 1607194113
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_233
timestamp 1607194113
transform 1 0 22540 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_221
timestamp 1607194113
transform 1 0 21436 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607194113
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607194113
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607194113
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1607194113
transform 1 0 4600 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_32
timestamp 1607194113
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607194113
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607194113
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1365_
timestamp 1607194113
transform 1 0 4692 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__CLK
timestamp 1607194113
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1607194113
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_60
timestamp 1607194113
transform 1 0 6624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_84
timestamp 1607194113
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607194113
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1363_
timestamp 1607194113
transform 1 0 9660 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_30_114
timestamp 1607194113
transform 1 0 11592 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__CLK
timestamp 1607194113
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1607194113
transform 1 0 11408 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1364_
timestamp 1607194113
transform 1 0 12144 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_30_154
timestamp 1607194113
transform 1 0 15272 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1607194113
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_139
timestamp 1607194113
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607194113
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_162
timestamp 1607194113
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__B1
timestamp 1607194113
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1320_
timestamp 1607194113
transform 1 0 16284 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_189
timestamp 1607194113
transform 1 0 18492 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_181
timestamp 1607194113
transform 1 0 17756 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0965_
timestamp 1607194113
transform 1 0 18768 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1607194113
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1607194113
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1607194113
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A2
timestamp 1607194113
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607194113
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1607194113
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1607194113
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607194113
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607194113
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1607194113
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1607194113
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1607194113
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1607194113
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_73
timestamp 1607194113
transform 1 0 7820 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_67
timestamp 1607194113
transform 1 0 7268 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1607194113
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__B1
timestamp 1607194113
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607194113
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1294_
timestamp 1607194113
transform 1 0 8096 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1607194113
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_92
timestamp 1607194113
transform 1 0 9568 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1607194113
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_105
timestamp 1607194113
transform 1 0 10764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A
timestamp 1607194113
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1607194113
transform 1 0 10304 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_133
timestamp 1607194113
transform 1 0 13340 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_127
timestamp 1607194113
transform 1 0 12788 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1607194113
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1607194113
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A
timestamp 1607194113
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607194113
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1607194113
transform 1 0 12880 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_157
timestamp 1607194113
transform 1 0 15548 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_145
timestamp 1607194113
transform 1 0 14444 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_175
timestamp 1607194113
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1607194113
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1607194113
transform 1 0 16836 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1607194113
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1607194113
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607194113
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1607194113
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1607194113
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1607194113
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1607194113
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607194113
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607194113
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_32
timestamp 1607194113
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1607194113
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607194113
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1607194113
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__B1
timestamp 1607194113
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1290_
timestamp 1607194113
transform 1 0 5152 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_72
timestamp 1607194113
transform 1 0 7728 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_60
timestamp 1607194113
transform 1 0 6624 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1607194113
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1607194113
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607194113
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_105
timestamp 1607194113
transform 1 0 10764 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B1
timestamp 1607194113
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1292_
timestamp 1607194113
transform 1 0 11224 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_138
timestamp 1607194113
transform 1 0 13800 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_126
timestamp 1607194113
transform 1 0 12696 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1607194113
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1607194113
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607194113
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1607194113
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607194113
transform 1 0 16560 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1607194113
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1607194113
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1607194113
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_199
timestamp 1607194113
transform 1 0 19412 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_i_A
timestamp 1607194113
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_i
timestamp 1607194113
transform 1 0 20148 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607194113
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__B1
timestamp 1607194113
transform 1 0 21252 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1318_
timestamp 1607194113
transform 1 0 21436 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607194113
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607194113
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1607194113
transform 1 0 2484 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607194113
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607194113
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607194113
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1498_
timestamp 1607194113
transform 1 0 2576 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1607194113
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607194113
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1607194113
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__CLK
timestamp 1607194113
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__D
timestamp 1607194113
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607194113
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1607194113
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1607194113
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1607194113
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1607194113
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1607194113
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1607194113
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_66
timestamp 1607194113
transform 1 0 7176 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607194113
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1607194113
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1283_
timestamp 1607194113
transform 1 0 8096 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1607194113
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1607194113
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_92
timestamp 1607194113
transform 1 0 9568 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_80
timestamp 1607194113
transform 1 0 8464 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607194113
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1607194113
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1607194113
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1607194113
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_107
timestamp 1607194113
transform 1 0 10948 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_100
timestamp 1607194113
transform 1 0 10304 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1289_
timestamp 1607194113
transform 1 0 10580 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1607194113
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1607194113
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1607194113
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607194113
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1607194113
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1607194113
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_143
timestamp 1607194113
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp 1607194113
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607194113
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0974_
timestamp 1607194113
transform 1 0 14720 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1607194113
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1607194113
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1607194113
transform 1 0 16652 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__C1
timestamp 1607194113
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B1
timestamp 1607194113
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1607194113
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_189
timestamp 1607194113
transform 1 0 18492 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1607194113
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1607194113
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607194113
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1607194113
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1607194113
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1607194113
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_213
timestamp 1607194113
transform 1 0 20700 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_201
timestamp 1607194113
transform 1 0 19596 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607194113
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1607194113
transform 1 0 21804 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607194113
transform 1 0 21988 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1317_
timestamp 1607194113
transform 1 0 22540 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_15
timestamp 1607194113
transform 1 0 2484 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1607194113
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607194113
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1362_
timestamp 1607194113
transform 1 0 2760 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_35_39
timestamp 1607194113
transform 1 0 4692 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__CLK
timestamp 1607194113
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_53
timestamp 1607194113
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_47
timestamp 1607194113
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1296_
timestamp 1607194113
transform 1 0 5612 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_70
timestamp 1607194113
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_62
timestamp 1607194113
transform 1 0 6808 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607194113
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1361_
timestamp 1607194113
transform 1 0 7728 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1607194113
transform 1 0 9660 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1607194113
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_117
timestamp 1607194113
transform 1 0 11868 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_105
timestamp 1607194113
transform 1 0 10764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1607194113
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607194113
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1403_
timestamp 1607194113
transform 1 0 12420 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1607194113
transform 1 0 15272 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_142
timestamp 1607194113
transform 1 0 14168 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1607194113
transform 1 0 15640 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_173
timestamp 1607194113
transform 1 0 17020 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_161
timestamp 1607194113
transform 1 0 15916 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1607194113
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1607194113
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1607194113
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607194113
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1607194113
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1607194113
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1607194113
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1607194113
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607194113
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607194113
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_37
timestamp 1607194113
transform 1 0 4508 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1607194113
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1607194113
transform 1 0 4324 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607194113
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 1607194113
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_57
timestamp 1607194113
transform 1 0 6348 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_49
timestamp 1607194113
transform 1 0 5612 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_78
timestamp 1607194113
transform 1 0 8280 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B1
timestamp 1607194113
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1299_
timestamp 1607194113
transform 1 0 6808 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1607194113
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_90
timestamp 1607194113
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607194113
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_109
timestamp 1607194113
transform 1 0 11132 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1607194113
transform 1 0 10764 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B1
timestamp 1607194113
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1229_
timestamp 1607194113
transform 1 0 11408 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_132
timestamp 1607194113
transform 1 0 13248 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A2_N
timestamp 1607194113
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B2
timestamp 1607194113
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1607194113
transform 1 0 13616 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_154
timestamp 1607194113
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1607194113
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1607194113
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607194113
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1607194113
transform 1 0 15548 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_173
timestamp 1607194113
transform 1 0 17020 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_161
timestamp 1607194113
transform 1 0 15916 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_181
timestamp 1607194113
transform 1 0 17756 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A1
timestamp 1607194113
transform 1 0 17940 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__B1
timestamp 1607194113
transform 1 0 18124 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _0981_
timestamp 1607194113
transform 1 0 18308 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1607194113
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1607194113
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_204
timestamp 1607194113
transform 1 0 19872 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607194113
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1607194113
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1607194113
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B1
timestamp 1607194113
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607194113
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1297_
timestamp 1607194113
transform 1 0 2668 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_33
timestamp 1607194113
transform 1 0 4140 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1607194113
transform 1 0 6348 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_45
timestamp 1607194113
transform 1 0 5244 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_74
timestamp 1607194113
transform 1 0 7912 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1607194113
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607194113
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_97
timestamp 1607194113
transform 1 0 10028 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_85
timestamp 1607194113
transform 1 0 8924 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A
timestamp 1607194113
transform 1 0 8740 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1607194113
transform 1 0 8464 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_109
timestamp 1607194113
transform 1 0 11132 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1607194113
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1607194113
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1607194113
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607194113
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0995_
timestamp 1607194113
transform 1 0 13708 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_37_154
timestamp 1607194113
transform 1 0 15272 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_178
timestamp 1607194113
transform 1 0 17480 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_166
timestamp 1607194113
transform 1 0 16376 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1607194113
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B1
timestamp 1607194113
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607194113
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0989_
timestamp 1607194113
transform 1 0 18216 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_37_214
timestamp 1607194113
transform 1 0 20792 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_203
timestamp 1607194113
transform 1 0 19780 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1607194113
transform 1 0 20516 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_226
timestamp 1607194113
transform 1 0 21896 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607194113
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607194113
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607194113
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_32
timestamp 1607194113
transform 1 0 4048 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607194113
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__B1
timestamp 1607194113
transform 1 0 4140 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607194113
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1301_
timestamp 1607194113
transform 1 0 4324 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_38_51
timestamp 1607194113
transform 1 0 5796 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_75
timestamp 1607194113
transform 1 0 8004 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_63
timestamp 1607194113
transform 1 0 6900 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1607194113
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1607194113
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_87
timestamp 1607194113
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607194113
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_117
timestamp 1607194113
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1607194113
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_125
timestamp 1607194113
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B1
timestamp 1607194113
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0992_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12972 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1607194113
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_150
timestamp 1607194113
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_142
timestamp 1607194113
transform 1 0 14168 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607194113
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_178
timestamp 1607194113
transform 1 0 17480 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1607194113
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_196
timestamp 1607194113
transform 1 0 19136 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_184
timestamp 1607194113
transform 1 0 18032 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1607194113
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1607194113
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_208
timestamp 1607194113
transform 1 0 20240 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607194113
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_227
timestamp 1607194113
transform 1 0 21988 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1607194113
transform 1 0 22540 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1607194113
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607194113
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607194113
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1607194113
transform 1 0 4140 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_27
timestamp 1607194113
transform 1 0 3588 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1360_
timestamp 1607194113
transform 1 0 4232 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_39_55
timestamp 1607194113
transform 1 0 6164 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1607194113
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_79
timestamp 1607194113
transform 1 0 8372 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_67
timestamp 1607194113
transform 1 0 7268 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1607194113
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607194113
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1607194113
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_91
timestamp 1607194113
transform 1 0 9476 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_115
timestamp 1607194113
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_103
timestamp 1607194113
transform 1 0 10580 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_136
timestamp 1607194113
transform 1 0 13616 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_130
timestamp 1607194113
transform 1 0 13064 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_123
timestamp 1607194113
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1607194113
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A1
timestamp 1607194113
transform 1 0 13708 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1607194113
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607194113
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1607194113
transform 1 0 12788 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_156
timestamp 1607194113
transform 1 0 15456 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__a2111o_4  _1001_
timestamp 1607194113
transform 1 0 13892 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_39_168
timestamp 1607194113
transform 1 0 16560 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_190
timestamp 1607194113
transform 1 0 18584 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_184
timestamp 1607194113
transform 1 0 18032 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1607194113
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1607194113
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607194113
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1007_
timestamp 1607194113
transform 1 0 18860 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_39_212
timestamp 1607194113
transform 1 0 20608 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_200
timestamp 1607194113
transform 1 0 19504 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_224
timestamp 1607194113
transform 1 0 21712 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1607194113
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1607194113
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1607194113
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1607194113
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607194113
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1607194113
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1607194113
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1607194113
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1607194113
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_292
timestamp 1607194113
transform 1 0 27968 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1607194113
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1607194113
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607194113
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_301
timestamp 1607194113
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1607194113
transform 1 0 28060 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_300
timestamp 1607194113
transform 1 0 28704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1607194113
transform -1 0 29256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607194113
transform -1 0 29256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1607194113
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1607194113
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1607194113
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1607194113
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1607194113
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607194113
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_300
timestamp 1607194113
transform 1 0 28704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607194113
transform -1 0 29256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1607194113
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1607194113
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1607194113
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607194113
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1607194113
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1607194113
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1607194113
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1607194113
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1607194113
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1607194113
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607194113
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_300
timestamp 1607194113
transform 1 0 28704 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_301
timestamp 1607194113
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_293
timestamp 1607194113
transform 1 0 28060 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607194113
transform -1 0 29256 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607194113
transform -1 0 29256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1607194113
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607194113
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_269
timestamp 1607194113
transform 1 0 25852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1607194113
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__CLK
timestamp 1607194113
transform 1 0 26036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__D
timestamp 1607194113
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1346_
timestamp 1607194113
transform 1 0 26404 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_5_302
timestamp 1607194113
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_294
timestamp 1607194113
transform 1 0 28152 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607194113
transform -1 0 29256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1607194113
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1607194113
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1607194113
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607194113
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1607194113
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1607194113
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1607194113
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1607194113
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_288
timestamp 1607194113
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1607194113
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607194113
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_301
timestamp 1607194113
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_293
timestamp 1607194113
transform 1 0 28060 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_300
timestamp 1607194113
transform 1 0 28704 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607194113
transform -1 0 29256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607194113
transform -1 0 29256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1607194113
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1607194113
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1607194113
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_288
timestamp 1607194113
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1607194113
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607194113
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_300
timestamp 1607194113
transform 1 0 28704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607194113
transform -1 0 29256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1607194113
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607194113
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1607194113
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1607194113
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1607194113
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_301
timestamp 1607194113
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_293
timestamp 1607194113
transform 1 0 28060 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607194113
transform -1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp 1607194113
transform 1 0 23276 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_235
timestamp 1607194113
transform 1 0 22724 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1607194113
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1607194113
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__CLK
timestamp 1607194113
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607194113
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1331_
timestamp 1607194113
transform 1 0 23644 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_264
timestamp 1607194113
transform 1 0 25392 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1607194113
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_288
timestamp 1607194113
transform 1 0 27600 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_276
timestamp 1607194113
transform 1 0 26496 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_288
timestamp 1607194113
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1607194113
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607194113
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_300
timestamp 1607194113
transform 1 0 28704 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_300
timestamp 1607194113
transform 1 0 28704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607194113
transform -1 0 29256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607194113
transform -1 0 29256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_245
timestamp 1607194113
transform 1 0 23644 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_269
timestamp 1607194113
transform 1 0 25852 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_257
timestamp 1607194113
transform 1 0 24748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_288
timestamp 1607194113
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1607194113
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607194113
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_300
timestamp 1607194113
transform 1 0 28704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607194113
transform -1 0 29256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_246
timestamp 1607194113
transform 1 0 23736 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_234
timestamp 1607194113
transform 1 0 22632 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1607194113
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1607194113
transform 1 0 23184 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607194113
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_270
timestamp 1607194113
transform 1 0 25944 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_258
timestamp 1607194113
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1607194113
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1607194113
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1607194113
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607194113
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1347_
timestamp 1607194113
transform 1 0 26496 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_14_295
timestamp 1607194113
transform 1 0 28244 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_301
timestamp 1607194113
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_293
timestamp 1607194113
transform 1 0 28060 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607194113
transform -1 0 29256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607194113
transform -1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1607194113
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1607194113
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607194113
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_265
timestamp 1607194113
transform 1 0 25484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_257
timestamp 1607194113
transform 1 0 24748 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__CLK
timestamp 1607194113
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1348_
timestamp 1607194113
transform 1 0 25760 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_287
timestamp 1607194113
transform 1 0 27508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_299
timestamp 1607194113
transform 1 0 28612 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607194113
transform -1 0 29256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1607194113
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1607194113
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1607194113
transform 1 0 22908 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1607194113
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1607194113
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607194113
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_257
timestamp 1607194113
transform 1 0 24748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1607194113
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__CLK
timestamp 1607194113
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1349_
timestamp 1607194113
transform 1 0 25208 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1607194113
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_288
timestamp 1607194113
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1607194113
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607194113
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_301
timestamp 1607194113
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_293
timestamp 1607194113
transform 1 0 28060 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_300
timestamp 1607194113
transform 1 0 28704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607194113
transform -1 0 29256 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607194113
transform -1 0 29256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1607194113
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1607194113
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_i_A
timestamp 1607194113
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_i
timestamp 1607194113
transform 1 0 22816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1607194113
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_288
timestamp 1607194113
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1607194113
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607194113
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_300
timestamp 1607194113
transform 1 0 28704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607194113
transform -1 0 29256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_251
timestamp 1607194113
transform 1 0 24196 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_245
timestamp 1607194113
transform 1 0 23644 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1607194113
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607194113
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1449_
timestamp 1607194113
transform 1 0 24472 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_19_285
timestamp 1607194113
transform 1 0 27324 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_273
timestamp 1607194113
transform 1 0 26220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_297
timestamp 1607194113
transform 1 0 28428 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607194113
transform -1 0 29256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1607194113
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_242
timestamp 1607194113
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_234
timestamp 1607194113
transform 1 0 22632 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_244
timestamp 1607194113
transform 1 0 23552 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__CLK
timestamp 1607194113
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607194113
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_263
timestamp 1607194113
transform 1 0 25300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_257
timestamp 1607194113
transform 1 0 24748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_272
timestamp 1607194113
transform 1 0 26128 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1607194113
transform 1 0 25760 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_256
timestamp 1607194113
transform 1 0 24656 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__B1
timestamp 1607194113
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1305_
timestamp 1607194113
transform 1 0 25576 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_282
timestamp 1607194113
transform 1 0 27048 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607194113
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1358_
timestamp 1607194113
transform 1 0 26496 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1607194113
transform 1 0 27784 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_301
timestamp 1607194113
transform 1 0 28796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_293
timestamp 1607194113
transform 1 0 28060 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_295
timestamp 1607194113
transform 1 0 28244 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607194113
transform -1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607194113
transform -1 0 29256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_250
timestamp 1607194113
transform 1 0 24104 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_238
timestamp 1607194113
transform 1 0 23000 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_262
timestamp 1607194113
transform 1 0 25208 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_288
timestamp 1607194113
transform 1 0 27600 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1607194113
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1607194113
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607194113
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_300
timestamp 1607194113
transform 1 0 28704 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607194113
transform -1 0 29256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1607194113
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607194113
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1607194113
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1607194113
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1607194113
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_301
timestamp 1607194113
transform 1 0 28796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_293
timestamp 1607194113
transform 1 0 28060 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607194113
transform -1 0 29256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_248
timestamp 1607194113
transform 1 0 23920 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_244
timestamp 1607194113
transform 1 0 23552 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B1
timestamp 1607194113
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1307_
timestamp 1607194113
transform 1 0 24196 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_267
timestamp 1607194113
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_291
timestamp 1607194113
transform 1 0 27876 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_279
timestamp 1607194113
transform 1 0 26772 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607194113
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 1607194113
transform 1 0 26496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607194113
transform -1 0 29256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_251
timestamp 1607194113
transform 1 0 24196 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_242
timestamp 1607194113
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_234
timestamp 1607194113
transform 1 0 22632 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1607194113
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607194113
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1159_
timestamp 1607194113
transform 1 0 23828 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__CLK
timestamp 1607194113
transform 1 0 24748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1357_
timestamp 1607194113
transform 1 0 24932 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_290
timestamp 1607194113
transform 1 0 27784 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_278
timestamp 1607194113
transform 1 0 26680 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_302
timestamp 1607194113
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607194113
transform -1 0 29256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_248
timestamp 1607194113
transform 1 0 23920 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_239
timestamp 1607194113
transform 1 0 23092 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk_i
timestamp 1607194113
transform 1 0 23644 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_272
timestamp 1607194113
transform 1 0 26128 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_260
timestamp 1607194113
transform 1 0 25024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607194113
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607194113
transform 1 0 26496 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_26_295
timestamp 1607194113
transform 1 0 28244 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607194113
transform -1 0 29256 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_244
timestamp 1607194113
transform 1 0 23552 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1607194113
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_241
timestamp 1607194113
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607194113
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_268
timestamp 1607194113
transform 1 0 25760 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_256
timestamp 1607194113
transform 1 0 24656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp 1607194113
transform 1 0 25852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1607194113
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1607194113
transform 1 0 27600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1607194113
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1607194113
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_291
timestamp 1607194113
transform 1 0 27876 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__B1
timestamp 1607194113
transform 1 0 26220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607194113
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1311_
timestamp 1607194113
transform 1 0 26404 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1607194113
transform 1 0 27968 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_295
timestamp 1607194113
transform 1 0 28244 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607194113
transform -1 0 29256 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607194113
transform -1 0 29256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_245
timestamp 1607194113
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_241
timestamp 1607194113
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607194113
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_253
timestamp 1607194113
transform 1 0 24380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__CLK
timestamp 1607194113
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1355_
timestamp 1607194113
transform 1 0 24840 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_29_289
timestamp 1607194113
transform 1 0 27692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_277
timestamp 1607194113
transform 1 0 26588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_301
timestamp 1607194113
transform 1 0 28796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607194113
transform -1 0 29256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_247
timestamp 1607194113
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_239
timestamp 1607194113
transform 1 0 23092 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B1
timestamp 1607194113
transform 1 0 24012 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1313_
timestamp 1607194113
transform 1 0 24196 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_267
timestamp 1607194113
transform 1 0 25668 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_292
timestamp 1607194113
transform 1 0 27968 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B1
timestamp 1607194113
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607194113
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1316_
timestamp 1607194113
transform 1 0 26496 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1607194113
transform 1 0 28704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607194113
transform -1 0 29256 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1607194113
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607194113
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_263
timestamp 1607194113
transform 1 0 25300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_257
timestamp 1607194113
transform 1 0 24748 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1607194113
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607194113
transform 1 0 25576 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_31_285
timestamp 1607194113
transform 1 0 27324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_297
timestamp 1607194113
transform 1 0 28428 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607194113
transform -1 0 29256 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_249
timestamp 1607194113
transform 1 0 24012 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1607194113
transform 1 0 22908 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_262
timestamp 1607194113
transform 1 0 25208 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_257
timestamp 1607194113
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1310_
timestamp 1607194113
transform 1 0 24840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_291
timestamp 1607194113
transform 1 0 27876 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_279
timestamp 1607194113
transform 1 0 26772 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1607194113
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607194113
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1607194113
transform 1 0 26496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607194113
transform -1 0 29256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_251
timestamp 1607194113
transform 1 0 24196 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1607194113
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1607194113
transform 1 0 24012 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607194113
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1607194113
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_271
timestamp 1607194113
transform 1 0 26036 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_263
timestamp 1607194113
transform 1 0 25300 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_289
timestamp 1607194113
transform 1 0 27692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_277
timestamp 1607194113
transform 1 0 26588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1607194113
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_301
timestamp 1607194113
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607194113
transform -1 0 29256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_245
timestamp 1607194113
transform 1 0 23644 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_248
timestamp 1607194113
transform 1 0 23920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__CLK
timestamp 1607194113
transform 1 0 23736 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1607194113
transform 1 0 24196 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607194113
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_272
timestamp 1607194113
transform 1 0 26128 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_272
timestamp 1607194113
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_260
timestamp 1607194113
transform 1 0 25024 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607194113
transform 1 0 24380 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_35_284
timestamp 1607194113
transform 1 0 27232 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_288
timestamp 1607194113
transform 1 0 27600 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1607194113
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607194113
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_302
timestamp 1607194113
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_296
timestamp 1607194113
transform 1 0 28336 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_300
timestamp 1607194113
transform 1 0 28704 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607194113
transform -1 0 29256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607194113
transform -1 0 29256 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_239
timestamp 1607194113
transform 1 0 23092 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__CLK
timestamp 1607194113
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1406_
timestamp 1607194113
transform 1 0 23828 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_36_266
timestamp 1607194113
transform 1 0 25576 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_288
timestamp 1607194113
transform 1 0 27600 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1607194113
transform 1 0 26496 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1607194113
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607194113
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_300
timestamp 1607194113
transform 1 0 28704 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607194113
transform -1 0 29256 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1607194113
transform 1 0 23644 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1607194113
transform 1 0 23000 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B1
timestamp 1607194113
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607194113
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1322_
timestamp 1607194113
transform 1 0 23736 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_37_262
timestamp 1607194113
transform 1 0 25208 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1321_
timestamp 1607194113
transform 1 0 25944 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_285
timestamp 1607194113
transform 1 0 27324 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_273
timestamp 1607194113
transform 1 0 26220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_297
timestamp 1607194113
transform 1 0 28428 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607194113
transform -1 0 29256 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1607194113
transform 1 0 23000 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1607194113
transform 1 0 22816 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__B1
timestamp 1607194113
transform 1 0 23368 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1324_
timestamp 1607194113
transform 1 0 23552 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_38_272
timestamp 1607194113
transform 1 0 26128 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_260
timestamp 1607194113
transform 1 0 25024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_291
timestamp 1607194113
transform 1 0 27876 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_279
timestamp 1607194113
transform 1 0 26772 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607194113
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1607194113
transform 1 0 26496 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607194113
transform -1 0 29256 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_245
timestamp 1607194113
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_236
timestamp 1607194113
transform 1 0 22816 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__CLK
timestamp 1607194113
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607194113
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1350_
timestamp 1607194113
transform 1 0 24104 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1607194113
transform 1 0 25852 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1607194113
transform 1 0 26956 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_301
timestamp 1607194113
transform 1 0 28796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_293
timestamp 1607194113
transform 1 0 28060 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607194113
transform -1 0 29256 0 1 23392
box -38 -48 314 592
use delayline_9_hd  inst_tdelay_line
timestamp 1607276172
transform 1 0 31280 0 1 4016
box 800 800 22236 22385
use delayline_9_hd  inst_idelay_line
timestamp 1607276172
transform 1 0 58696 0 1 4016
box 800 800 22236 22385
use delayline_9_hd  inst_rdelay_line
timestamp 1607276172
transform 1 0 86020 0 1 4016
box 800 800 22236 22385
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1607194113
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1607194113
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607194113
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_32
timestamp 1607194113
transform 1 0 4048 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1607194113
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607194113
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_58
timestamp 1607194113
transform 1 0 6440 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__B1
timestamp 1607194113
transform 1 0 4784 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1303_
timestamp 1607194113
transform 1 0 4968 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_70
timestamp 1607194113
transform 1 0 7544 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1607194113
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1607194113
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_82
timestamp 1607194113
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607194113
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_105
timestamp 1607194113
transform 1 0 10764 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__CLK
timestamp 1607194113
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1402_
timestamp 1607194113
transform 1 0 11224 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1607194113
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1607194113
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1607194113
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607194113
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_178
timestamp 1607194113
transform 1 0 17480 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1607194113
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_192
timestamp 1607194113
transform 1 0 18768 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_184
timestamp 1607194113
transform 1 0 18032 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1005_
timestamp 1607194113
transform 1 0 18124 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1607194113
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_212
timestamp 1607194113
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_204
timestamp 1607194113
transform 1 0 19872 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607194113
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_227
timestamp 1607194113
transform 1 0 21988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1607194113
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1607194113
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1607194113
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1607194113
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607194113
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607194113
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1607194113
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1607194113
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_39
timestamp 1607194113
transform 1 0 4692 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1607194113
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607194113
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_48
timestamp 1607194113
transform 1 0 5520 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_44
timestamp 1607194113
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_55
timestamp 1607194113
transform 1 0 6164 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C
timestamp 1607194113
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1607194113
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1359_
timestamp 1607194113
transform 1 0 5612 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1011_
timestamp 1607194113
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_42_70
timestamp 1607194113
transform 1 0 7544 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_79
timestamp 1607194113
transform 1 0 8372 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_67
timestamp 1607194113
transform 1 0 7268 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1607194113
transform 1 0 7360 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1607194113
transform 1 0 7084 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607194113
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1607194113
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1607194113
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_90
timestamp 1607194113
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_82
timestamp 1607194113
transform 1 0 8648 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_91
timestamp 1607194113
transform 1 0 9476 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607194113
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_115
timestamp 1607194113
transform 1 0 11684 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_103
timestamp 1607194113
transform 1 0 10580 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B1
timestamp 1607194113
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1230_
timestamp 1607194113
transform 1 0 10948 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_42_127
timestamp 1607194113
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_123
timestamp 1607194113
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1607194113
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A2_N
timestamp 1607194113
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B2
timestamp 1607194113
transform 1 0 12420 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1607194113
transform 1 0 12604 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607194113
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1607194113
transform 1 0 12972 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0950_
timestamp 1607194113
transform 1 0 13156 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_135
timestamp 1607194113
transform 1 0 13524 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _0998_
timestamp 1607194113
transform 1 0 12788 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_42_147
timestamp 1607194113
transform 1 0 14628 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_152
timestamp 1607194113
transform 1 0 15088 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_140
timestamp 1607194113
transform 1 0 13984 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607194113
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1020_
timestamp 1607194113
transform 1 0 15272 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1607194113
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_176
timestamp 1607194113
transform 1 0 17296 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_164
timestamp 1607194113
transform 1 0 16192 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_192
timestamp 1607194113
transform 1 0 18768 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1607194113
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_182
timestamp 1607194113
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B1
timestamp 1607194113
transform 1 0 18032 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607194113
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 18952 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1009_
timestamp 1607194113
transform 1 0 18216 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_42_215
timestamp 1607194113
transform 1 0 20884 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_211
timestamp 1607194113
transform 1 0 20516 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_203
timestamp 1607194113
transform 1 0 19780 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_211
timestamp 1607194113
transform 1 0 20516 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_207
timestamp 1607194113
transform 1 0 20148 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_199
timestamp 1607194113
transform 1 0 19412 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607194113
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1607194113
transform 1 0 20240 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1607194113
transform 1 0 21436 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_223
timestamp 1607194113
transform 1 0 21620 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B2
timestamp 1607194113
transform 1 0 21528 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0972_
timestamp 1607194113
transform 1 0 21712 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1607194113
transform 1 0 2484 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1607194113
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607194113
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1500_
timestamp 1607194113
transform 1 0 2576 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_43_37
timestamp 1607194113
transform 1 0 4508 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__CLK
timestamp 1607194113
transform 1 0 4324 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_49
timestamp 1607194113
transform 1 0 5612 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1607194113
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1607194113
transform 1 0 7912 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607194113
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0680_
timestamp 1607194113
transform 1 0 8096 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_92
timestamp 1607194113
transform 1 0 9568 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_80
timestamp 1607194113
transform 1 0 8464 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_116
timestamp 1607194113
transform 1 0 11776 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_104
timestamp 1607194113
transform 1 0 10672 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1607194113
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1607194113
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607194113
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_155
timestamp 1607194113
transform 1 0 15364 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_43_147
timestamp 1607194113
transform 1 0 14628 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1607194113
transform 1 0 14904 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1607194113
transform 1 0 15088 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_178
timestamp 1607194113
transform 1 0 17480 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_166
timestamp 1607194113
transform 1 0 16376 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1607194113
transform 1 0 15916 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1607194113
transform 1 0 16100 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1607194113
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_184
timestamp 1607194113
transform 1 0 18032 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_182
timestamp 1607194113
transform 1 0 17848 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1607194113
transform 1 0 18308 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607194113
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1017_
timestamp 1607194113
transform 1 0 18492 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1607194113
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1607194113
transform 1 0 22448 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1607194113
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1607194113
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1607194113
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607194113
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1607194113
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607194113
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1022_
timestamp 1607194113
transform 1 0 4048 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_45
timestamp 1607194113
transform 1 0 5244 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1607194113
transform 1 0 6440 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__C
timestamp 1607194113
transform 1 0 5060 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B
timestamp 1607194113
transform 1 0 6256 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1607194113
transform 1 0 4876 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1004_
timestamp 1607194113
transform 1 0 5612 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_44_72
timestamp 1607194113
transform 1 0 7728 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_60
timestamp 1607194113
transform 1 0 6624 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1607194113
transform 1 0 8004 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0667_
timestamp 1607194113
transform 1 0 8188 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_98
timestamp 1607194113
transform 1 0 10120 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_89
timestamp 1607194113
transform 1 0 9292 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_81
timestamp 1607194113
transform 1 0 8556 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1607194113
transform 1 0 9936 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607194113
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1607194113
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_108
timestamp 1607194113
transform 1 0 11040 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0949_
timestamp 1607194113
transform 1 0 10672 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_132
timestamp 1607194113
transform 1 0 13248 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_120
timestamp 1607194113
transform 1 0 12144 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1607194113
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1607194113
transform 1 0 15088 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1607194113
transform 1 0 14352 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607194113
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_172
timestamp 1607194113
transform 1 0 16928 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_166
timestamp 1607194113
transform 1 0 16376 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1607194113
transform 1 0 17020 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0957_
timestamp 1607194113
transform 1 0 17204 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_44_182
timestamp 1607194113
transform 1 0 17848 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1021_
timestamp 1607194113
transform 1 0 18584 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1607194113
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_211
timestamp 1607194113
transform 1 0 20516 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_199
timestamp 1607194113
transform 1 0 19412 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607194113
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_227
timestamp 1607194113
transform 1 0 21988 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B2
timestamp 1607194113
transform 1 0 22540 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1607194113
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1607194113
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607194113
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_27
timestamp 1607194113
transform 1 0 3588 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1607194113
transform 1 0 4600 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B
timestamp 1607194113
transform 1 0 4416 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1012_
timestamp 1607194113
transform 1 0 3772 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_45_52
timestamp 1607194113
transform 1 0 5888 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_40
timestamp 1607194113
transform 1 0 4784 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1607194113
transform 1 0 7452 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_62
timestamp 1607194113
transform 1 0 6808 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_60
timestamp 1607194113
transform 1 0 6624 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1607194113
transform 1 0 6992 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__C
timestamp 1607194113
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1607194113
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607194113
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8188 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1607194113
transform 1 0 7176 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_94
timestamp 1607194113
transform 1 0 9752 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_86
timestamp 1607194113
transform 1 0 9016 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0948_
timestamp 1607194113
transform 1 0 9844 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_45_116
timestamp 1607194113
transform 1 0 11776 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_104
timestamp 1607194113
transform 1 0 10672 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_135
timestamp 1607194113
transform 1 0 13524 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1607194113
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607194113
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_141
timestamp 1607194113
transform 1 0 14076 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 14168 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1607194113
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_159
timestamp 1607194113
transform 1 0 15732 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1607194113
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1607194113
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607194113
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1607194113
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_232
timestamp 1607194113
transform 1 0 22448 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_220
timestamp 1607194113
transform 1 0 21344 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1607194113
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1607194113
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607194113
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1607194113
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1607194113
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607194113
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_56
timestamp 1607194113
transform 1 0 6256 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1607194113
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_67
timestamp 1607194113
transform 1 0 7268 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_62
timestamp 1607194113
transform 1 0 6808 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B
timestamp 1607194113
transform 1 0 7820 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1607194113
transform 1 0 6900 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _0669_
timestamp 1607194113
transform 1 0 8004 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_46_84
timestamp 1607194113
transform 1 0 8832 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607194113
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1003_
timestamp 1607194113
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_46_114
timestamp 1607194113
transform 1 0 11592 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_102
timestamp 1607194113
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1607194113
transform 1 0 11224 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_128
timestamp 1607194113
transform 1 0 12880 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_122
timestamp 1607194113
transform 1 0 12328 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13616 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1607194113
transform 1 0 12512 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_145
timestamp 1607194113
transform 1 0 14444 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607194113
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0941_
timestamp 1607194113
transform 1 0 15272 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_46_173
timestamp 1607194113
transform 1 0 17020 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_161
timestamp 1607194113
transform 1 0 15916 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_185
timestamp 1607194113
transform 1 0 18124 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A1
timestamp 1607194113
transform 1 0 18216 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1000_
timestamp 1607194113
transform 1 0 18400 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1607194113
transform 1 0 20884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1607194113
transform 1 0 20700 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1607194113
transform 1 0 20332 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A3
timestamp 1607194113
transform 1 0 20148 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B1
timestamp 1607194113
transform 1 0 19964 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607194113
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_227
timestamp 1607194113
transform 1 0 21988 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0670_
timestamp 1607194113
transform 1 0 22540 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_15
timestamp 1607194113
transform 1 0 2484 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1607194113
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607194113
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1501_
timestamp 1607194113
transform 1 0 2576 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_47_37
timestamp 1607194113
transform 1 0 4508 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__CLK
timestamp 1607194113
transform 1 0 4324 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_49
timestamp 1607194113
transform 1 0 5612 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1607194113
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1607194113
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607194113
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0679_
timestamp 1607194113
transform 1 0 8096 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_92
timestamp 1607194113
transform 1 0 9568 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_80
timestamp 1607194113
transform 1 0 8464 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__C
timestamp 1607194113
transform 1 0 9752 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0907_
timestamp 1607194113
transform 1 0 9936 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_117
timestamp 1607194113
transform 1 0 11868 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_105
timestamp 1607194113
transform 1 0 10764 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_135
timestamp 1607194113
transform 1 0 13524 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1607194113
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_121
timestamp 1607194113
transform 1 0 12236 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607194113
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_153
timestamp 1607194113
transform 1 0 15180 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_141
timestamp 1607194113
transform 1 0 14076 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__D
timestamp 1607194113
transform 1 0 14996 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0999_
timestamp 1607194113
transform 1 0 14168 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_47_168
timestamp 1607194113
transform 1 0 16560 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1158_
timestamp 1607194113
transform 1 0 15732 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_184
timestamp 1607194113
transform 1 0 18032 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_180
timestamp 1607194113
transform 1 0 17664 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A1
timestamp 1607194113
transform 1 0 18400 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607194113
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0994_
timestamp 1607194113
transform 1 0 18584 0 1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_47_211
timestamp 1607194113
transform 1 0 20516 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A3
timestamp 1607194113
transform 1 0 20332 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B1
timestamp 1607194113
transform 1 0 20148 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0977_
timestamp 1607194113
transform 1 0 20884 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_47_224
timestamp 1607194113
transform 1 0 21712 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1607194113
transform 1 0 21528 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_15
timestamp 1607194113
transform 1 0 2484 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1607194113
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1607194113
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1607194113
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607194113
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607194113
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1503_
timestamp 1607194113
transform 1 0 2760 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1607194113
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_38
timestamp 1607194113
transform 1 0 4600 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1607194113
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__CLK
timestamp 1607194113
transform 1 0 4508 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1607194113
transform 1 0 4416 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607194113
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1607194113
transform 1 0 4048 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_59
timestamp 1607194113
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_51
timestamp 1607194113
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_50
timestamp 1607194113
transform 1 0 5704 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_74
timestamp 1607194113
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1607194113
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_74
timestamp 1607194113
transform 1 0 7912 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_62
timestamp 1607194113
transform 1 0 6808 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1607194113
transform 1 0 8004 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607194113
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1607194113
transform 1 0 8188 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_98
timestamp 1607194113
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_86
timestamp 1607194113
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1607194113
transform 1 0 10028 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1607194113
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607194113
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0905_
timestamp 1607194113
transform 1 0 9660 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_110
timestamp 1607194113
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_114
timestamp 1607194113
transform 1 0 11592 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_109
timestamp 1607194113
transform 1 0 11132 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0908_
timestamp 1607194113
transform 1 0 11224 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_132
timestamp 1607194113
transform 1 0 13248 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_134
timestamp 1607194113
transform 1 0 13432 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_126
timestamp 1607194113
transform 1 0 12696 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1607194113
transform 1 0 13064 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607194113
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0993_
timestamp 1607194113
transform 1 0 13616 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1607194113
transform 1 0 12420 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_49_144
timestamp 1607194113
transform 1 0 14352 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_147
timestamp 1607194113
transform 1 0 14628 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__D
timestamp 1607194113
transform 1 0 14444 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1607194113
transform 1 0 14444 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0682_
timestamp 1607194113
transform 1 0 14628 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_48_154
timestamp 1607194113
transform 1 0 15272 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__C
timestamp 1607194113
transform 1 0 14996 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1607194113
transform 1 0 15364 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607194113
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1219_
timestamp 1607194113
transform 1 0 15548 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_49_156
timestamp 1607194113
transform 1 0 15456 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_168
timestamp 1607194113
transform 1 0 16560 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1607194113
transform 1 0 17480 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1607194113
transform 1 0 16376 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_196
timestamp 1607194113
transform 1 0 19136 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1607194113
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_180
timestamp 1607194113
transform 1 0 17664 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_190
timestamp 1607194113
transform 1 0 18584 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607194113
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_204
timestamp 1607194113
transform 1 0 19872 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1607194113
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_202
timestamp 1607194113
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1607194113
transform 1 0 21068 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_i
timestamp 1607194113
transform 1 0 20148 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607194113
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0970_
timestamp 1607194113
transform 1 0 20424 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_49_233
timestamp 1607194113
transform 1 0 22540 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_221
timestamp 1607194113
transform 1 0 21436 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1607194113
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_i_A
timestamp 1607194113
transform 1 0 21252 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1607194113
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1607194113
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607194113
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_38
timestamp 1607194113
transform 1 0 4600 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_32
timestamp 1607194113
transform 1 0 4048 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1607194113
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607194113
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1497_
timestamp 1607194113
transform 1 0 4692 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__CLK
timestamp 1607194113
transform 1 0 6440 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_72
timestamp 1607194113
transform 1 0 7728 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_60
timestamp 1607194113
transform 1 0 6624 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_84
timestamp 1607194113
transform 1 0 8832 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__CLK
timestamp 1607194113
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607194113
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1376_
timestamp 1607194113
transform 1 0 9660 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_112
timestamp 1607194113
transform 1 0 11408 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_136
timestamp 1607194113
transform 1 0 13616 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_124
timestamp 1607194113
transform 1 0 12512 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_158
timestamp 1607194113
transform 1 0 15640 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_152
timestamp 1607194113
transform 1 0 15088 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_148
timestamp 1607194113
transform 1 0 14720 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607194113
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1025_
timestamp 1607194113
transform 1 0 15272 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_170
timestamp 1607194113
transform 1 0 16744 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_191
timestamp 1607194113
transform 1 0 18676 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1607194113
transform 1 0 17848 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1607194113
transform 1 0 19228 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0962_
timestamp 1607194113
transform 1 0 18032 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1607194113
transform 1 0 20884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_206
timestamp 1607194113
transform 1 0 20056 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607194113
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0984_
timestamp 1607194113
transform 1 0 19412 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1607194113
transform 1 0 21988 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_15
timestamp 1607194113
transform 1 0 2484 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1607194113
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607194113
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1499_
timestamp 1607194113
transform 1 0 2576 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1607194113
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__CLK
timestamp 1607194113
transform 1 0 4508 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__D
timestamp 1607194113
transform 1 0 4324 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_59
timestamp 1607194113
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_51
timestamp 1607194113
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_75
timestamp 1607194113
transform 1 0 8004 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_70
timestamp 1607194113
transform 1 0 7544 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_62
timestamp 1607194113
transform 1 0 6808 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk_i
timestamp 1607194113
transform 1 0 7728 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607194113
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_87
timestamp 1607194113
transform 1 0 9108 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A3
timestamp 1607194113
transform 1 0 9844 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1271_
timestamp 1607194113
transform 1 0 10028 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1607194113
transform 1 0 11960 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__B1
timestamp 1607194113
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A2
timestamp 1607194113
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_135
timestamp 1607194113
transform 1 0 13524 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1607194113
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607194113
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_155
timestamp 1607194113
transform 1 0 15364 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_147
timestamp 1607194113
transform 1 0 14628 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1607194113
transform 1 0 15456 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_171
timestamp 1607194113
transform 1 0 16836 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_159
timestamp 1607194113
transform 1 0 15732 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_196
timestamp 1607194113
transform 1 0 19136 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1607194113
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607194113
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_207
timestamp 1607194113
transform 1 0 20148 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_202
timestamp 1607194113
transform 1 0 19688 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0961_
timestamp 1607194113
transform 1 0 19780 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_233
timestamp 1607194113
transform 1 0 22540 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_219
timestamp 1607194113
transform 1 0 21252 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1607194113
transform 1 0 22356 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 21528 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1607194113
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1607194113
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607194113
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_32
timestamp 1607194113
transform 1 0 4048 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1607194113
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607194113
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_40
timestamp 1607194113
transform 1 0 4784 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1505_
timestamp 1607194113
transform 1 0 4876 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_52_74
timestamp 1607194113
transform 1 0 7912 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_62
timestamp 1607194113
transform 1 0 6808 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__CLK
timestamp 1607194113
transform 1 0 6624 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_93
timestamp 1607194113
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_86
timestamp 1607194113
transform 1 0 9016 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607194113
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_105
timestamp 1607194113
transform 1 0 10764 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A3
timestamp 1607194113
transform 1 0 10948 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1272_
timestamp 1607194113
transform 1 0 11132 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_52_130
timestamp 1607194113
transform 1 0 13064 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B1
timestamp 1607194113
transform 1 0 12880 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A2
timestamp 1607194113
transform 1 0 12696 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_154
timestamp 1607194113
transform 1 0 15272 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_150
timestamp 1607194113
transform 1 0 14904 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_142
timestamp 1607194113
transform 1 0 14168 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607194113
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_166
timestamp 1607194113
transform 1 0 16376 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__CLK
timestamp 1607194113
transform 1 0 16468 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1372_
timestamp 1607194113
transform 1 0 16652 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_52_196
timestamp 1607194113
transform 1 0 19136 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1607194113
transform 1 0 18400 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1607194113
transform 1 0 20884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_211
timestamp 1607194113
transform 1 0 20516 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_203
timestamp 1607194113
transform 1 0 19780 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607194113
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1607194113
transform 1 0 19412 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1607194113
transform 1 0 21988 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1607194113
transform 1 0 2484 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1607194113
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607194113
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1506_
timestamp 1607194113
transform 1 0 2852 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__CLK
timestamp 1607194113
transform 1 0 4600 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_52
timestamp 1607194113
transform 1 0 5888 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_40
timestamp 1607194113
transform 1 0 4784 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_74
timestamp 1607194113
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1607194113
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_60
timestamp 1607194113
transform 1 0 6624 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607194113
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_98
timestamp 1607194113
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_86
timestamp 1607194113
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_114
timestamp 1607194113
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_110
timestamp 1607194113
transform 1 0 11224 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_i_A
timestamp 1607194113
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_i
timestamp 1607194113
transform 1 0 11684 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_135
timestamp 1607194113
transform 1 0 13524 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1607194113
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_120
timestamp 1607194113
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607194113
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_155
timestamp 1607194113
transform 1 0 15364 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_147
timestamp 1607194113
transform 1 0 14628 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1233_
timestamp 1607194113
transform 1 0 15548 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_53_176
timestamp 1607194113
transform 1 0 17296 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_164
timestamp 1607194113
transform 1 0 16192 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1607194113
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1607194113
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1607194113
transform 1 0 17848 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607194113
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1607194113
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_232
timestamp 1607194113
transform 1 0 22448 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_220
timestamp 1607194113
transform 1 0 21344 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1607194113
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1607194113
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607194113
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1607194113
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1607194113
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607194113
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1607194113
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1607194113
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1607194113
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1607194113
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_80
timestamp 1607194113
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607194113
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1607194113
transform 1 0 10764 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1375_
timestamp 1607194113
transform 1 0 10948 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_54_138
timestamp 1607194113
transform 1 0 13800 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_126
timestamp 1607194113
transform 1 0 12696 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_154
timestamp 1607194113
transform 1 0 15272 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_150
timestamp 1607194113
transform 1 0 14904 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607194113
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_162
timestamp 1607194113
transform 1 0 16008 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A2
timestamp 1607194113
transform 1 0 16192 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A3
timestamp 1607194113
transform 1 0 16376 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1275_
timestamp 1607194113
transform 1 0 16560 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_54_187
timestamp 1607194113
transform 1 0 18308 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B1
timestamp 1607194113
transform 1 0 18124 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_215
timestamp 1607194113
transform 1 0 20884 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_206
timestamp 1607194113
transform 1 0 20056 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607194113
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1013_
timestamp 1607194113
transform 1 0 19412 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1607194113
transform 1 0 21988 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1607194113
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1607194113
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1607194113
transform 1 0 2484 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1607194113
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607194113
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607194113
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1504_
timestamp 1607194113
transform 1 0 2852 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1607194113
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1607194113
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__CLK
timestamp 1607194113
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607194113
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1607194113
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1607194113
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_52
timestamp 1607194113
transform 1 0 5888 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_40
timestamp 1607194113
transform 1 0 4784 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_74
timestamp 1607194113
transform 1 0 7912 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_68
timestamp 1607194113
transform 1 0 7360 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1607194113
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_60
timestamp 1607194113
transform 1 0 6624 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607194113
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0934_
timestamp 1607194113
transform 1 0 8004 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0926_
timestamp 1607194113
transform 1 0 7912 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_56_86
timestamp 1607194113
transform 1 0 9016 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_85
timestamp 1607194113
transform 1 0 8924 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B
timestamp 1607194113
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B
timestamp 1607194113
transform 1 0 8740 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607194113
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0936_
timestamp 1607194113
transform 1 0 9660 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0932_
timestamp 1607194113
transform 1 0 9476 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_56_116
timestamp 1607194113
transform 1 0 11776 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_104
timestamp 1607194113
transform 1 0 10672 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_114
timestamp 1607194113
transform 1 0 11592 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_102
timestamp 1607194113
transform 1 0 10488 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B
timestamp 1607194113
transform 1 0 10488 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B
timestamp 1607194113
transform 1 0 10304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_128
timestamp 1607194113
transform 1 0 12880 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_135
timestamp 1607194113
transform 1 0 13524 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1607194113
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607194113
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_148
timestamp 1607194113
transform 1 0 14720 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_140
timestamp 1607194113
transform 1 0 13984 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_155
timestamp 1607194113
transform 1 0 15364 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_147
timestamp 1607194113
transform 1 0 14628 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__CLK
timestamp 1607194113
transform 1 0 14996 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607194113
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1518_
timestamp 1607194113
transform 1 0 15272 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0867_
timestamp 1607194113
transform 1 0 15640 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_173
timestamp 1607194113
transform 1 0 17020 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_173
timestamp 1607194113
transform 1 0 17020 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_162
timestamp 1607194113
transform 1 0 16008 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1607194113
transform 1 0 16744 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_196
timestamp 1607194113
transform 1 0 19136 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_184
timestamp 1607194113
transform 1 0 18032 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_193
timestamp 1607194113
transform 1 0 18860 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_184
timestamp 1607194113
transform 1 0 18032 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_181
timestamp 1607194113
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A
timestamp 1607194113
transform 1 0 17572 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607194113
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1607194113
transform 1 0 18584 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1607194113
transform 1 0 17756 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_213
timestamp 1607194113
transform 1 0 20700 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_205
timestamp 1607194113
transform 1 0 19964 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_200
timestamp 1607194113
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_201
timestamp 1607194113
transform 1 0 19596 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607194113
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1240_
timestamp 1607194113
transform 1 0 20884 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1235_
timestamp 1607194113
transform 1 0 19596 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _1006_
timestamp 1607194113
transform 1 0 19780 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_231
timestamp 1607194113
transform 1 0 22356 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_219
timestamp 1607194113
transform 1 0 21252 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1607194113
transform 1 0 21804 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__B1
timestamp 1607194113
transform 1 0 21620 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A1_N
timestamp 1607194113
transform 1 0 21436 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A2_N
timestamp 1607194113
transform 1 0 21252 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_15
timestamp 1607194113
transform 1 0 2484 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1607194113
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607194113
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1507_
timestamp 1607194113
transform 1 0 2576 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1607194113
transform 1 0 4508 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__CLK
timestamp 1607194113
transform 1 0 4324 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_49
timestamp 1607194113
transform 1 0 5612 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_72
timestamp 1607194113
transform 1 0 7728 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_62
timestamp 1607194113
transform 1 0 6808 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607194113
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1607194113
transform 1 0 7360 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1607194113
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_80
timestamp 1607194113
transform 1 0 8464 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B
timestamp 1607194113
transform 1 0 9568 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0928_
timestamp 1607194113
transform 1 0 8740 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1607194113
transform 1 0 11960 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_106
timestamp 1607194113
transform 1 0 10856 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_135
timestamp 1607194113
transform 1 0 13524 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1607194113
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607194113
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_156
timestamp 1607194113
transform 1 0 15456 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_147
timestamp 1607194113
transform 1 0 14628 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1607194113
transform 1 0 14996 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1607194113
transform 1 0 15180 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_177
timestamp 1607194113
transform 1 0 17388 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1607194113
transform 1 0 17204 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1023_
timestamp 1607194113
transform 1 0 16560 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_57_195
timestamp 1607194113
transform 1 0 19044 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1607194113
transform 1 0 18860 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1607194113
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607194113
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0674_
timestamp 1607194113
transform 1 0 18032 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_207
timestamp 1607194113
transform 1 0 20148 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_203
timestamp 1607194113
transform 1 0 19780 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1607194113
transform 1 0 19872 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_231
timestamp 1607194113
transform 1 0 22356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_219
timestamp 1607194113
transform 1 0 21252 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1607194113
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1607194113
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607194113
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_32
timestamp 1607194113
transform 1 0 4048 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1607194113
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1607194113
transform 1 0 4324 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607194113
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1607194113
transform 1 0 4508 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_52
timestamp 1607194113
transform 1 0 5888 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_40
timestamp 1607194113
transform 1 0 4784 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0895_
timestamp 1607194113
transform 1 0 5520 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_76
timestamp 1607194113
transform 1 0 8096 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_64
timestamp 1607194113
transform 1 0 6992 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1607194113
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_88
timestamp 1607194113
transform 1 0 9200 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk_i
timestamp 1607194113
transform 1 0 9292 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607194113
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_105
timestamp 1607194113
transform 1 0 10764 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__CLK
timestamp 1607194113
transform 1 0 11500 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1519_
timestamp 1607194113
transform 1 0 11684 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_58_134
timestamp 1607194113
transform 1 0 13432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_154
timestamp 1607194113
transform 1 0 15272 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_152
timestamp 1607194113
transform 1 0 15088 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_146
timestamp 1607194113
transform 1 0 14536 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607194113
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1326_
timestamp 1607194113
transform 1 0 15548 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_170
timestamp 1607194113
transform 1 0 16744 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__B
timestamp 1607194113
transform 1 0 16560 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A
timestamp 1607194113
transform 1 0 16376 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_196
timestamp 1607194113
transform 1 0 19136 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp 1607194113
transform 1 0 18952 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 17848 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_215
timestamp 1607194113
transform 1 0 20884 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_58_208
timestamp 1607194113
transform 1 0 20240 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607194113
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_228
timestamp 1607194113
transform 1 0 22080 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_223
timestamp 1607194113
transform 1 0 21620 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0924_
timestamp 1607194113
transform 1 0 21712 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1607194113
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607194113
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607194113
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_35
timestamp 1607194113
transform 1 0 4324 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_27
timestamp 1607194113
transform 1 0 3588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0921_
timestamp 1607194113
transform 1 0 4600 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_59_49
timestamp 1607194113
transform 1 0 5612 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1607194113
transform 1 0 5428 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_69
timestamp 1607194113
transform 1 0 7452 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_62
timestamp 1607194113
transform 1 0 6808 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607194113
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0938_
timestamp 1607194113
transform 1 0 8188 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0861_
timestamp 1607194113
transform 1 0 7084 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1607194113
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1607194113
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1607194113
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_133
timestamp 1607194113
transform 1 0 13340 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_129
timestamp 1607194113
transform 1 0 12972 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_123
timestamp 1607194113
transform 1 0 12420 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607194113
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1607194113
transform 1 0 13064 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_145
timestamp 1607194113
transform 1 0 14444 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__B1
timestamp 1607194113
transform 1 0 14996 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1325_
timestamp 1607194113
transform 1 0 15180 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_177
timestamp 1607194113
transform 1 0 17388 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_165
timestamp 1607194113
transform 1 0 16284 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1607194113
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1607194113
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607194113
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0937_
timestamp 1607194113
transform 1 0 20240 0 1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_59_230
timestamp 1607194113
transform 1 0 22264 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B2
timestamp 1607194113
transform 1 0 22080 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A2
timestamp 1607194113
transform 1 0 21896 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1
timestamp 1607194113
transform 1 0 21712 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1607194113
transform 1 0 21528 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607194113
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607194113
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607194113
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_36
timestamp 1607194113
transform 1 0 4416 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1607194113
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607194113
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607194113
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0899_
timestamp 1607194113
transform 1 0 4508 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_60_48
timestamp 1607194113
transform 1 0 5520 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1607194113
transform 1 0 5336 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0912_
timestamp 1607194113
transform 1 0 6072 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_75
timestamp 1607194113
transform 1 0 8004 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_63
timestamp 1607194113
transform 1 0 6900 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1607194113
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_91
timestamp 1607194113
transform 1 0 9476 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_87
timestamp 1607194113
transform 1 0 9108 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607194113
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1607194113
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1607194113
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_137
timestamp 1607194113
transform 1 0 13708 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_129
timestamp 1607194113
transform 1 0 12972 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_154
timestamp 1607194113
transform 1 0 15272 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_152
timestamp 1607194113
transform 1 0 15088 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_144
timestamp 1607194113
transform 1 0 14352 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A
timestamp 1607194113
transform 1 0 13892 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607194113
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1607194113
transform 1 0 14076 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_172
timestamp 1607194113
transform 1 0 16928 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_166
timestamp 1607194113
transform 1 0 16376 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1607194113
transform 1 0 17388 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0665_
timestamp 1607194113
transform 1 0 17020 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_191
timestamp 1607194113
transform 1 0 18676 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_179
timestamp 1607194113
transform 1 0 17572 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_211
timestamp 1607194113
transform 1 0 20516 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_203
timestamp 1607194113
transform 1 0 19780 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607194113
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1607194113
transform 1 0 20884 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1607194113
transform 1 0 22540 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1607194113
transform 1 0 21436 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1607194113
transform 1 0 21252 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1607194113
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607194113
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_15
timestamp 1607194113
transform 1 0 2484 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607194113
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607194113
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607194113
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1508_
timestamp 1607194113
transform 1 0 2576 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1607194113
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1607194113
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_37
timestamp 1607194113
transform 1 0 4508 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__CLK
timestamp 1607194113
transform 1 0 4324 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1607194113
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_54
timestamp 1607194113
transform 1 0 6072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_44
timestamp 1607194113
transform 1 0 5152 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_54
timestamp 1607194113
transform 1 0 6072 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1607194113
transform 1 0 5888 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0914_
timestamp 1607194113
transform 1 0 5244 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0901_
timestamp 1607194113
transform 1 0 5060 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_78
timestamp 1607194113
transform 1 0 8280 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1607194113
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_78
timestamp 1607194113
transform 1 0 8280 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_74
timestamp 1607194113
transform 1 0 7912 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1607194113
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_60
timestamp 1607194113
transform 1 0 6624 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1607194113
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1502_
timestamp 1607194113
transform 1 0 8372 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1607194113
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_90
timestamp 1607194113
transform 1 0 9384 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__CLK
timestamp 1607194113
transform 1 0 10120 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1607194113
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1607194113
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1607194113
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_112
timestamp 1607194113
transform 1 0 11408 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_100
timestamp 1607194113
transform 1 0 10304 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1607194113
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_131
timestamp 1607194113
transform 1 0 13156 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_123
timestamp 1607194113
transform 1 0 12420 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_120
timestamp 1607194113
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1607194113
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13340 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_62_149
timestamp 1607194113
transform 1 0 14812 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1607194113
transform 1 0 14076 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_146
timestamp 1607194113
transform 1 0 14536 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1607194113
transform 1 0 14996 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B1
timestamp 1607194113
transform 1 0 15088 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1607194113
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0916_
timestamp 1607194113
transform 1 0 15272 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _0909_
timestamp 1607194113
transform 1 0 15272 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_168
timestamp 1607194113
transform 1 0 16560 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_170
timestamp 1607194113
transform 1 0 16744 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_i_A
timestamp 1607194113
transform 1 0 17388 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 1607194113
transform 1 0 16376 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A2
timestamp 1607194113
transform 1 0 16560 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1607194113
transform 1 0 16376 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_i
timestamp 1607194113
transform 1 0 17112 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_191
timestamp 1607194113
transform 1 0 18676 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_179
timestamp 1607194113
transform 1 0 17572 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1607194113
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1607194113
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 1607194113
transform 1 0 17848 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1607194113
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_206
timestamp 1607194113
transform 1 0 20056 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_199
timestamp 1607194113
transform 1 0 19412 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_213
timestamp 1607194113
transform 1 0 20700 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_208
timestamp 1607194113
transform 1 0 20240 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1607194113
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0920_
timestamp 1607194113
transform 1 0 20884 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1607194113
transform 1 0 19688 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1607194113
transform 1 0 20332 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1607194113
transform 1 0 22540 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_227
timestamp 1607194113
transform 1 0 21988 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B1
timestamp 1607194113
transform 1 0 22356 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A2
timestamp 1607194113
transform 1 0 22172 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1607194113
transform 1 0 21804 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1607194113
transform 1 0 21436 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1607194113
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607194113
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607194113
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_27
timestamp 1607194113
transform 1 0 3588 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B1
timestamp 1607194113
transform 1 0 3680 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1258_
timestamp 1607194113
transform 1 0 3864 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_63_52
timestamp 1607194113
transform 1 0 5888 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A2_N
timestamp 1607194113
transform 1 0 5704 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B2
timestamp 1607194113
transform 1 0 5520 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A1_N
timestamp 1607194113
transform 1 0 5336 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_74
timestamp 1607194113
transform 1 0 7912 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1607194113
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_60
timestamp 1607194113
transform 1 0 6624 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1607194113
transform 1 0 8188 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1607194113
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0911_
timestamp 1607194113
transform 1 0 8372 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_63_97
timestamp 1607194113
transform 1 0 10028 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A2
timestamp 1607194113
transform 1 0 9844 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1607194113
transform 1 0 9660 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_109
timestamp 1607194113
transform 1 0 11132 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1607194113
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1607194113
transform 1 0 12236 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1607194113
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0910_
timestamp 1607194113
transform 1 0 13524 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_63_156
timestamp 1607194113
transform 1 0 15456 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_148
timestamp 1607194113
transform 1 0 14720 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_170
timestamp 1607194113
transform 1 0 16744 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B
timestamp 1607194113
transform 1 0 16560 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1607194113
transform 1 0 16376 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0915_
timestamp 1607194113
transform 1 0 15732 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1607194113
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1607194113
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_182
timestamp 1607194113
transform 1 0 17848 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1607194113
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_208
timestamp 1607194113
transform 1 0 20240 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _0898_
timestamp 1607194113
transform 1 0 20792 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1607194113
transform 1 0 22448 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1607194113
transform 1 0 22264 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1607194113
transform 1 0 22080 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1607194113
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1607194113
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607194113
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_32
timestamp 1607194113
transform 1 0 4048 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1607194113
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1607194113
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1385_
timestamp 1607194113
transform 1 0 4140 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_54
timestamp 1607194113
transform 1 0 6072 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1607194113
transform 1 0 5888 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_78
timestamp 1607194113
transform 1 0 8280 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_66
timestamp 1607194113
transform 1 0 7176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1607194113
transform 1 0 9384 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1607194113
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0913_
timestamp 1607194113
transform 1 0 9660 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_64_111
timestamp 1607194113
transform 1 0 11316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1607194113
transform 1 0 11132 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1607194113
transform 1 0 10948 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_135
timestamp 1607194113
transform 1 0 13524 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_123
timestamp 1607194113
transform 1 0 12420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_147
timestamp 1607194113
transform 1 0 14628 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1607194113
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0903_
timestamp 1607194113
transform 1 0 15272 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_64_175
timestamp 1607194113
transform 1 0 17204 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_163
timestamp 1607194113
transform 1 0 16100 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B
timestamp 1607194113
transform 1 0 15916 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1607194113
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_199
timestamp 1607194113
transform 1 0 19412 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk_i
timestamp 1607194113
transform 1 0 20516 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1607194113
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0900_
timestamp 1607194113
transform 1 0 20884 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A2
timestamp 1607194113
transform 1 0 22540 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1607194113
transform 1 0 22356 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1607194113
transform 1 0 22172 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_19
timestamp 1607194113
transform 1 0 2852 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_15
timestamp 1607194113
transform 1 0 2484 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607194113
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607194113
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1_N
timestamp 1607194113
transform 1 0 4600 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B1
timestamp 1607194113
transform 1 0 2944 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1257_
timestamp 1607194113
transform 1 0 3128 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_65_52
timestamp 1607194113
transform 1 0 5888 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_48
timestamp 1607194113
transform 1 0 5520 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_44
timestamp 1607194113
transform 1 0 5152 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A2_N
timestamp 1607194113
transform 1 0 4968 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B2
timestamp 1607194113
transform 1 0 4784 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1607194113
transform 1 0 5612 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_74
timestamp 1607194113
transform 1 0 7912 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_62
timestamp 1607194113
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_60
timestamp 1607194113
transform 1 0 6624 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1607194113
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_86
timestamp 1607194113
transform 1 0 9016 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B1
timestamp 1607194113
transform 1 0 9292 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1195_
timestamp 1607194113
transform 1 0 9476 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_109
timestamp 1607194113
transform 1 0 11132 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A1_N
timestamp 1607194113
transform 1 0 10948 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_138
timestamp 1607194113
transform 1 0 13800 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_126
timestamp 1607194113
transform 1 0 12696 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_121
timestamp 1607194113
transform 1 0 12236 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1607194113
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1607194113
transform 1 0 12420 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_150
timestamp 1607194113
transform 1 0 14904 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_170
timestamp 1607194113
transform 1 0 16744 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_162
timestamp 1607194113
transform 1 0 16008 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A
timestamp 1607194113
transform 1 0 16560 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1255_
timestamp 1607194113
transform 1 0 16192 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1607194113
transform 1 0 19136 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1607194113
transform 1 0 18032 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_182
timestamp 1607194113
transform 1 0 17848 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1607194113
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_208
timestamp 1607194113
transform 1 0 20240 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B1
timestamp 1607194113
transform 1 0 20424 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1254_
timestamp 1607194113
transform 1 0 20608 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_230
timestamp 1607194113
transform 1 0 22264 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A1_N
timestamp 1607194113
transform 1 0 22080 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1607194113
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1607194113
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607194113
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1607194113
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1607194113
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1607194113
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1607194113
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1607194113
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1607194113
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_93
timestamp 1607194113
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_80
timestamp 1607194113
transform 1 0 8464 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1607194113
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1426_
timestamp 1607194113
transform 1 0 10764 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_138
timestamp 1607194113
transform 1 0 13800 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_126
timestamp 1607194113
transform 1 0 12696 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_150
timestamp 1607194113
transform 1 0 14904 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B1
timestamp 1607194113
transform 1 0 14996 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1607194113
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1256_
timestamp 1607194113
transform 1 0 15272 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_172
timestamp 1607194113
transform 1 0 16928 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B2
timestamp 1607194113
transform 1 0 16744 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1607194113
transform 1 0 17480 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_195
timestamp 1607194113
transform 1 0 19044 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_183
timestamp 1607194113
transform 1 0 17940 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1607194113
transform 1 0 17756 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_215
timestamp 1607194113
transform 1 0 20884 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_213
timestamp 1607194113
transform 1 0 20700 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_207
timestamp 1607194113
transform 1 0 20148 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1607194113
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__CLK
timestamp 1607194113
transform 1 0 21252 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1388_
timestamp 1607194113
transform 1 0 21436 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_67_19
timestamp 1607194113
transform 1 0 2852 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_15
timestamp 1607194113
transform 1 0 2484 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1607194113
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607194113
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__CLK
timestamp 1607194113
transform 1 0 4692 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1386_
timestamp 1607194113
transform 1 0 2944 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_67_53
timestamp 1607194113
transform 1 0 5980 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_41
timestamp 1607194113
transform 1 0 4876 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_74
timestamp 1607194113
transform 1 0 7912 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1607194113
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__B1
timestamp 1607194113
transform 1 0 8096 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1607194113
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1194_
timestamp 1607194113
transform 1 0 8280 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_96
timestamp 1607194113
transform 1 0 9936 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1_N
timestamp 1607194113
transform 1 0 9752 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_108
timestamp 1607194113
transform 1 0 11040 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_135
timestamp 1607194113
transform 1 0 13524 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_123
timestamp 1607194113
transform 1 0 12420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_120
timestamp 1607194113
transform 1 0 12144 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk_i
timestamp 1607194113
transform 1 0 13800 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1607194113
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_147
timestamp 1607194113
transform 1 0 14628 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_141
timestamp 1607194113
transform 1 0 14076 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__B1
timestamp 1607194113
transform 1 0 14720 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1193_
timestamp 1607194113
transform 1 0 14904 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_67_178
timestamp 1607194113
transform 1 0 17480 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_166
timestamp 1607194113
transform 1 0 16376 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1607194113
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1607194113
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1607194113
transform 1 0 17848 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1607194113
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1607194113
transform 1 0 20240 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_232
timestamp 1607194113
transform 1 0 22448 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_220
timestamp 1607194113
transform 1 0 21344 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1607194113
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1607194113
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1607194113
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1607194113
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607194113
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607194113
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1607194113
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1607194113
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_36
timestamp 1607194113
transform 1 0 4416 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_32
timestamp 1607194113
transform 1 0 4048 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1607194113
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1607194113
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1607194113
transform 1 0 4508 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_59
timestamp 1607194113
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_51
timestamp 1607194113
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_52
timestamp 1607194113
transform 1 0 5888 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_40
timestamp 1607194113
transform 1 0 4784 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_74
timestamp 1607194113
transform 1 0 7912 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_62
timestamp 1607194113
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_76
timestamp 1607194113
transform 1 0 8096 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_64
timestamp 1607194113
transform 1 0 6992 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1607194113
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_82
timestamp 1607194113
transform 1 0 8648 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_93
timestamp 1607194113
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_88
timestamp 1607194113
transform 1 0 9200 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1607194113
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1427_
timestamp 1607194113
transform 1 0 8740 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_69_116
timestamp 1607194113
transform 1 0 11776 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_104
timestamp 1607194113
transform 1 0 10672 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_117
timestamp 1607194113
transform 1 0 11868 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_105
timestamp 1607194113
transform 1 0 10764 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1607194113
transform 1 0 10488 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_135
timestamp 1607194113
transform 1 0 13524 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_123
timestamp 1607194113
transform 1 0 12420 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_129
timestamp 1607194113
transform 1 0 12972 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1607194113
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_155
timestamp 1607194113
transform 1 0 15364 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_147
timestamp 1607194113
transform 1 0 14628 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_154
timestamp 1607194113
transform 1 0 15272 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1607194113
transform 1 0 14076 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1607194113
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1192_
timestamp 1607194113
transform 1 0 15640 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_177
timestamp 1607194113
transform 1 0 17388 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_170
timestamp 1607194113
transform 1 0 16744 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_164
timestamp 1607194113
transform 1 0 16192 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_162
timestamp 1607194113
transform 1 0 16008 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1607194113
transform 1 0 17204 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1607194113
transform 1 0 16008 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1387_
timestamp 1607194113
transform 1 0 16100 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1248_
timestamp 1607194113
transform 1 0 16836 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_189
timestamp 1607194113
transform 1 0 18492 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_196
timestamp 1607194113
transform 1 0 19136 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_184
timestamp 1607194113
transform 1 0 18032 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__CLK
timestamp 1607194113
transform 1 0 17848 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1607194113
transform 1 0 18308 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1607194113
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1607194113
transform 1 0 18032 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_213
timestamp 1607194113
transform 1 0 20700 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_201
timestamp 1607194113
transform 1 0 19596 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_215
timestamp 1607194113
transform 1 0 20884 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_208
timestamp 1607194113
transform 1 0 20240 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1607194113
transform 1 0 20976 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1607194113
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1191_
timestamp 1607194113
transform 1 0 21160 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1607194113
transform 1 0 21804 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1607194113
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1607194113
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607194113
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_32
timestamp 1607194113
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1607194113
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1607194113
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_56
timestamp 1607194113
transform 1 0 6256 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_44
timestamp 1607194113
transform 1 0 5152 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0886_
timestamp 1607194113
transform 1 0 5428 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_73
timestamp 1607194113
transform 1 0 7820 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0894_
timestamp 1607194113
transform 1 0 6992 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_70_93
timestamp 1607194113
transform 1 0 9660 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1607194113
transform 1 0 9476 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_85
timestamp 1607194113
transform 1 0 8924 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1607194113
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1607194113
transform 1 0 10212 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_114
timestamp 1607194113
transform 1 0 11592 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_102
timestamp 1607194113
transform 1 0 10488 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_127
timestamp 1607194113
transform 1 0 12788 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_122
timestamp 1607194113
transform 1 0 12328 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1607194113
transform 1 0 12512 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_154
timestamp 1607194113
transform 1 0 15272 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_151
timestamp 1607194113
transform 1 0 14996 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_139
timestamp 1607194113
transform 1 0 13892 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1607194113
transform 1 0 15548 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1607194113
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_178
timestamp 1607194113
transform 1 0 17480 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1428_
timestamp 1607194113
transform 1 0 15732 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_70_190
timestamp 1607194113
transform 1 0 18584 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0885_
timestamp 1607194113
transform 1 0 18768 0 -1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_70_215
timestamp 1607194113
transform 1 0 20884 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_210
timestamp 1607194113
transform 1 0 20424 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B1
timestamp 1607194113
transform 1 0 20240 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A1
timestamp 1607194113
transform 1 0 20056 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1607194113
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_223
timestamp 1607194113
transform 1 0 21620 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1607194113
transform 1 0 21896 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1429_
timestamp 1607194113
transform 1 0 22080 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_71_15
timestamp 1607194113
transform 1 0 2484 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607194113
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607194113
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1509_
timestamp 1607194113
transform 1 0 2576 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_71_37
timestamp 1607194113
transform 1 0 4508 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__CLK
timestamp 1607194113
transform 1 0 4324 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_53
timestamp 1607194113
transform 1 0 5980 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_43
timestamp 1607194113
transform 1 0 5060 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0888_
timestamp 1607194113
transform 1 0 5152 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_71
timestamp 1607194113
transform 1 0 7636 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1607194113
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0892_
timestamp 1607194113
transform 1 0 6808 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_71_95
timestamp 1607194113
transform 1 0 9844 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_83
timestamp 1607194113
transform 1 0 8740 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1607194113
transform 1 0 9936 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1251_
timestamp 1607194113
transform 1 0 10120 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_71_116
timestamp 1607194113
transform 1 0 11776 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A1_N
timestamp 1607194113
transform 1 0 11592 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_123
timestamp 1607194113
transform 1 0 12420 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1607194113
transform 1 0 12604 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1
timestamp 1607194113
transform 1 0 12788 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1607194113
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0893_
timestamp 1607194113
transform 1 0 12972 0 1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_71_155
timestamp 1607194113
transform 1 0 15364 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_143
timestamp 1607194113
transform 1 0 14260 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_167
timestamp 1607194113
transform 1 0 16468 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_190
timestamp 1607194113
transform 1 0 18584 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_184
timestamp 1607194113
transform 1 0 18032 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_179
timestamp 1607194113
transform 1 0 17572 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1607194113
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0883_
timestamp 1607194113
transform 1 0 18676 0 1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_71_217
timestamp 1607194113
transform 1 0 21068 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1607194113
transform 1 0 19964 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_229
timestamp 1607194113
transform 1 0 22172 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1607194113
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607194113
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607194113
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_32
timestamp 1607194113
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1607194113
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1607194113
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_44
timestamp 1607194113
transform 1 0 5152 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0884_
timestamp 1607194113
transform 1 0 5888 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_73
timestamp 1607194113
transform 1 0 7820 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_61
timestamp 1607194113
transform 1 0 6716 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0880_
timestamp 1607194113
transform 1 0 7452 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_93
timestamp 1607194113
transform 1 0 9660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_91
timestamp 1607194113
transform 1 0 9476 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_85
timestamp 1607194113
transform 1 0 8924 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1607194113
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_105
timestamp 1607194113
transform 1 0 10764 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1390_
timestamp 1607194113
transform 1 0 11040 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_129
timestamp 1607194113
transform 1 0 12972 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1607194113
transform 1 0 12788 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_154
timestamp 1607194113
transform 1 0 15272 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1607194113
transform 1 0 14076 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1607194113
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_167
timestamp 1607194113
transform 1 0 16468 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_160
timestamp 1607194113
transform 1 0 15824 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1607194113
transform 1 0 16284 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1607194113
transform 1 0 15916 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_191
timestamp 1607194113
transform 1 0 18676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_179
timestamp 1607194113
transform 1 0 17572 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_215
timestamp 1607194113
transform 1 0 20884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_211
timestamp 1607194113
transform 1 0 20516 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_203
timestamp 1607194113
transform 1 0 19780 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1607194113
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_227
timestamp 1607194113
transform 1 0 21988 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_15
timestamp 1607194113
transform 1 0 2484 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1607194113
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607194113
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1344_
timestamp 1607194113
transform 1 0 2576 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1607194113
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__CLK
timestamp 1607194113
transform 1 0 4508 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__D
timestamp 1607194113
transform 1 0 4324 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_59
timestamp 1607194113
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_51
timestamp 1607194113
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_73
timestamp 1607194113
transform 1 0 7820 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_68
timestamp 1607194113
transform 1 0 7360 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_62
timestamp 1607194113
transform 1 0 6808 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1607194113
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0862_
timestamp 1607194113
transform 1 0 7452 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_97
timestamp 1607194113
transform 1 0 10028 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_85
timestamp 1607194113
transform 1 0 8924 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_109
timestamp 1607194113
transform 1 0 11132 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_135
timestamp 1607194113
transform 1 0 13524 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_123
timestamp 1607194113
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_121
timestamp 1607194113
transform 1 0 12236 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1607194113
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_147
timestamp 1607194113
transform 1 0 14628 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_177
timestamp 1607194113
transform 1 0 17388 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_165
timestamp 1607194113
transform 1 0 16284 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1607194113
transform 1 0 16100 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1607194113
transform 1 0 15732 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_184
timestamp 1607194113
transform 1 0 18032 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1607194113
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0887_
timestamp 1607194113
transform 1 0 18216 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_73_216
timestamp 1607194113
transform 1 0 20976 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_204
timestamp 1607194113
transform 1 0 19872 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1
timestamp 1607194113
transform 1 0 19688 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A1
timestamp 1607194113
transform 1 0 19504 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_228
timestamp 1607194113
transform 1 0 22080 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_15
timestamp 1607194113
transform 1 0 2484 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1607194113
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1607194113
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1607194113
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607194113
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607194113
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1482_
timestamp 1607194113
transform 1 0 2576 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1607194113
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1607194113
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1607194113
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__CLK
timestamp 1607194113
transform 1 0 4508 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__D
timestamp 1607194113
transform 1 0 4324 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1607194113
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_59
timestamp 1607194113
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_51
timestamp 1607194113
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_56
timestamp 1607194113
transform 1 0 6256 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1607194113
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_70
timestamp 1607194113
transform 1 0 7544 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_62
timestamp 1607194113
transform 1 0 6808 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_73
timestamp 1607194113
transform 1 0 7820 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B
timestamp 1607194113
transform 1 0 7636 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1607194113
transform 1 0 7636 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1607194113
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1188_
timestamp 1607194113
transform 1 0 7820 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _0873_
timestamp 1607194113
transform 1 0 6808 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_91
timestamp 1607194113
transform 1 0 9476 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_93
timestamp 1607194113
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1607194113
transform 1 0 9476 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1607194113
transform 1 0 8924 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1_N
timestamp 1607194113
transform 1 0 9292 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1607194113
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_115
timestamp 1607194113
transform 1 0 11684 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_103
timestamp 1607194113
transform 1 0 10580 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_117
timestamp 1607194113
transform 1 0 11868 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_105
timestamp 1607194113
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_123
timestamp 1607194113
transform 1 0 12420 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1607194113
transform 1 0 12236 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_129
timestamp 1607194113
transform 1 0 12972 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B1
timestamp 1607194113
transform 1 0 12604 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1607194113
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1250_
timestamp 1607194113
transform 1 0 12788 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0891_
timestamp 1607194113
transform 1 0 13064 0 -1 42976
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_75_156
timestamp 1607194113
transform 1 0 15456 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_143
timestamp 1607194113
transform 1 0 14260 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_154
timestamp 1607194113
transform 1 0 15272 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_152
timestamp 1607194113
transform 1 0 15088 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_144
timestamp 1607194113
transform 1 0 14352 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1607194113
transform 1 0 15272 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1607194113
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1607194113
transform 1 0 14996 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_168
timestamp 1607194113
transform 1 0 16560 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_178
timestamp 1607194113
transform 1 0 17480 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_166
timestamp 1607194113
transform 1 0 16376 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_180
timestamp 1607194113
transform 1 0 17664 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_190
timestamp 1607194113
transform 1 0 18584 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__B1
timestamp 1607194113
transform 1 0 17756 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1607194113
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1249_
timestamp 1607194113
transform 1 0 18032 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_202
timestamp 1607194113
transform 1 0 19688 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_202
timestamp 1607194113
transform 1 0 19688 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A1_N
timestamp 1607194113
transform 1 0 19504 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__B1
timestamp 1607194113
transform 1 0 20056 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1607194113
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1186_
timestamp 1607194113
transform 1 0 20240 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _0864_
timestamp 1607194113
transform 1 0 20884 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_226
timestamp 1607194113
transform 1 0 21896 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1607194113
transform 1 0 22540 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1607194113
transform 1 0 21436 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1607194113
transform 1 0 22264 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1607194113
transform 1 0 21252 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1_N
timestamp 1607194113
transform 1 0 21712 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1607194113
transform 1 0 22448 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607194113
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607194113
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607194113
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1607194113
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607194113
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1607194113
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_56
timestamp 1607194113
transform 1 0 6256 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1607194113
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_73
timestamp 1607194113
transform 1 0 7820 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1607194113
transform 1 0 7636 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0871_
timestamp 1607194113
transform 1 0 6808 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_76_96
timestamp 1607194113
transform 1 0 9936 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_91
timestamp 1607194113
transform 1 0 9476 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_85
timestamp 1607194113
transform 1 0 8924 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1607194113
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1607194113
transform 1 0 9660 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_108
timestamp 1607194113
transform 1 0 11040 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_124
timestamp 1607194113
transform 1 0 12512 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_120
timestamp 1607194113
transform 1 0 12144 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B1
timestamp 1607194113
transform 1 0 12604 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1187_
timestamp 1607194113
transform 1 0 12788 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_76_151
timestamp 1607194113
transform 1 0 14996 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_143
timestamp 1607194113
transform 1 0 14260 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1607194113
transform 1 0 15548 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1607194113
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1607194113
transform 1 0 15272 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_171
timestamp 1607194113
transform 1 0 16836 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_159
timestamp 1607194113
transform 1 0 15732 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1185_
timestamp 1607194113
transform 1 0 17204 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_193
timestamp 1607194113
transform 1 0 18860 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_181
timestamp 1607194113
transform 1 0 17756 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1607194113
transform 1 0 17572 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_218
timestamp 1607194113
transform 1 0 21160 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_213
timestamp 1607194113
transform 1 0 20700 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_205
timestamp 1607194113
transform 1 0 19964 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1607194113
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1607194113
transform 1 0 20884 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1433_
timestamp 1607194113
transform 1 0 21896 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_77_15
timestamp 1607194113
transform 1 0 2484 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1607194113
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1607194113
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1513_
timestamp 1607194113
transform 1 0 2576 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_77_37
timestamp 1607194113
transform 1 0 4508 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__CLK
timestamp 1607194113
transform 1 0 4324 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_49
timestamp 1607194113
transform 1 0 5612 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_70
timestamp 1607194113
transform 1 0 7544 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_62
timestamp 1607194113
transform 1 0 6808 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1607194113
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1431_
timestamp 1607194113
transform 1 0 7636 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_77_92
timestamp 1607194113
transform 1 0 9568 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1607194113
transform 1 0 9384 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_116
timestamp 1607194113
transform 1 0 11776 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_104
timestamp 1607194113
transform 1 0 10672 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_135
timestamp 1607194113
transform 1 0 13524 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_123
timestamp 1607194113
transform 1 0 12420 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1607194113
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1391_
timestamp 1607194113
transform 1 0 13708 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_77_158
timestamp 1607194113
transform 1 0 15640 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__CLK
timestamp 1607194113
transform 1 0 15456 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_170
timestamp 1607194113
transform 1 0 16744 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_190
timestamp 1607194113
transform 1 0 18584 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_184
timestamp 1607194113
transform 1 0 18032 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_182
timestamp 1607194113
transform 1 0 17848 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1607194113
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1392_
timestamp 1607194113
transform 1 0 18676 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_77_212
timestamp 1607194113
transform 1 0 20608 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__CLK
timestamp 1607194113
transform 1 0 20424 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_224
timestamp 1607194113
transform 1 0 21712 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1607194113
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1607194113
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1607194113
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1607194113
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_27
timestamp 1607194113
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1607194113
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_44
timestamp 1607194113
transform 1 0 5152 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1514_
timestamp 1607194113
transform 1 0 5336 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_78_79
timestamp 1607194113
transform 1 0 8372 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_67
timestamp 1607194113
transform 1 0 7268 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__CLK
timestamp 1607194113
transform 1 0 7084 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_93
timestamp 1607194113
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_91
timestamp 1607194113
transform 1 0 9476 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1607194113
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_117
timestamp 1607194113
transform 1 0 11868 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_105
timestamp 1607194113
transform 1 0 10764 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_129
timestamp 1607194113
transform 1 0 12972 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_154
timestamp 1607194113
transform 1 0 15272 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1607194113
transform 1 0 14076 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1607194113
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_178
timestamp 1607194113
transform 1 0 17480 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_166
timestamp 1607194113
transform 1 0 16376 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_190
timestamp 1607194113
transform 1 0 18584 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_215
timestamp 1607194113
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_202
timestamp 1607194113
transform 1 0 19688 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1607194113
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_227
timestamp 1607194113
transform 1 0 21988 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_15
timestamp 1607194113
transform 1 0 2484 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1607194113
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1607194113
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1511_
timestamp 1607194113
transform 1 0 2576 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_79_37
timestamp 1607194113
transform 1 0 4508 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__CLK
timestamp 1607194113
transform 1 0 4324 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_49
timestamp 1607194113
transform 1 0 5612 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_74
timestamp 1607194113
transform 1 0 7912 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_62
timestamp 1607194113
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1607194113
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_98
timestamp 1607194113
transform 1 0 10120 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_86
timestamp 1607194113
transform 1 0 9016 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_110
timestamp 1607194113
transform 1 0 11224 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_131
timestamp 1607194113
transform 1 0 13156 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_123
timestamp 1607194113
transform 1 0 12420 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1607194113
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1432_
timestamp 1607194113
transform 1 0 13432 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_79_155
timestamp 1607194113
transform 1 0 15364 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1607194113
transform 1 0 15180 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_167
timestamp 1607194113
transform 1 0 16468 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1607194113
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1607194113
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_179
timestamp 1607194113
transform 1 0 17572 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1607194113
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_208
timestamp 1607194113
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_232
timestamp 1607194113
transform 1 0 22448 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_220
timestamp 1607194113
transform 1 0 21344 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_235
timestamp 1607194113
transform 1 0 22724 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B1
timestamp 1607194113
transform 1 0 23000 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1225_
timestamp 1607194113
transform 1 0 23184 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_40_272
timestamp 1607194113
transform 1 0 26128 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_260
timestamp 1607194113
transform 1 0 25024 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B2
timestamp 1607194113
transform 1 0 24840 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A2_N
timestamp 1607194113
transform 1 0 24656 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1607194113
transform 1 0 26956 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1607194113
transform 1 0 26772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607194113
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1607194113
transform 1 0 26496 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_293
timestamp 1607194113
transform 1 0 28060 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[2]
timestamp 1607194113
transform 1 0 28796 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607194113
transform -1 0 29256 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1607194113
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_235
timestamp 1607194113
transform 1 0 22724 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A2
timestamp 1607194113
transform 1 0 23184 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1607194113
transform 1 0 23000 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_248
timestamp 1607194113
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_249
timestamp 1607194113
transform 1 0 24012 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_245
timestamp 1607194113
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1607194113
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__B1
timestamp 1607194113
transform 1 0 24012 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607194113
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1228_
timestamp 1607194113
transform 1 0 24104 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _1231_
timestamp 1607194113
transform 1 0 24196 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_42_269
timestamp 1607194113
transform 1 0 25852 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_254
timestamp 1607194113
transform 1 0 24472 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__CLK
timestamp 1607194113
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A2_N
timestamp 1607194113
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1401_
timestamp 1607194113
transform 1 0 25208 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_42_292
timestamp 1607194113
transform 1 0 27968 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_280
timestamp 1607194113
transform 1 0 26864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1607194113
transform 1 0 26956 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607194113
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1221_
timestamp 1607194113
transform 1 0 26496 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_300
timestamp 1607194113
transform 1 0 28704 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1607194113
transform 1 0 28796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_293
timestamp 1607194113
transform 1 0 28060 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607194113
transform -1 0 29256 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607194113
transform -1 0 29256 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1607194113
transform 1 0 23644 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607194113
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_269
timestamp 1607194113
transform 1 0 25852 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1607194113
transform 1 0 24748 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1607194113
transform 1 0 26956 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_301
timestamp 1607194113
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_293
timestamp 1607194113
transform 1 0 28060 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607194113
transform -1 0 29256 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A2
timestamp 1607194113
transform 1 0 24196 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A1
timestamp 1607194113
transform 1 0 24012 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0979_
timestamp 1607194113
transform 1 0 22724 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_44_272
timestamp 1607194113
transform 1 0 26128 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_260
timestamp 1607194113
transform 1 0 25024 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_255
timestamp 1607194113
transform 1 0 24564 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B1
timestamp 1607194113
transform 1 0 24380 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1607194113
transform 1 0 24748 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1607194113
transform 1 0 27600 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_276
timestamp 1607194113
transform 1 0 26496 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607194113
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1607194113
transform 1 0 27968 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_297
timestamp 1607194113
transform 1 0 28428 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1607194113
transform 1 0 28244 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607194113
transform -1 0 29256 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_249
timestamp 1607194113
transform 1 0 24012 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607194113
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1224_
timestamp 1607194113
transform 1 0 23644 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1607194113
transform 1 0 25116 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1220_
timestamp 1607194113
transform 1 0 24748 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_273
timestamp 1607194113
transform 1 0 26220 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__CLK
timestamp 1607194113
transform 1 0 26312 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1400_
timestamp 1607194113
transform 1 0 26496 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_45_295
timestamp 1607194113
transform 1 0 28244 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607194113
transform -1 0 29256 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_249
timestamp 1607194113
transform 1 0 24012 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1607194113
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B2
timestamp 1607194113
transform 1 0 24104 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0987_
timestamp 1607194113
transform 1 0 24288 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_46_270
timestamp 1607194113
transform 1 0 25944 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B1
timestamp 1607194113
transform 1 0 25760 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 1607194113
transform 1 0 25576 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_292
timestamp 1607194113
transform 1 0 27968 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B1
timestamp 1607194113
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607194113
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1232_
timestamp 1607194113
transform 1 0 26496 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_46_300
timestamp 1607194113
transform 1 0 28704 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607194113
transform -1 0 29256 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_245
timestamp 1607194113
transform 1 0 23644 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_236
timestamp 1607194113
transform 1 0 22816 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607194113
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_269
timestamp 1607194113
transform 1 0 25852 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A2
timestamp 1607194113
transform 1 0 24380 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1015_
timestamp 1607194113
transform 1 0 24564 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1607194113
transform 1 0 26956 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_301
timestamp 1607194113
transform 1 0 28796 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_293
timestamp 1607194113
transform 1 0 28060 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607194113
transform -1 0 29256 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1607194113
transform 1 0 24012 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_241
timestamp 1607194113
transform 1 0 23276 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_251
timestamp 1607194113
transform 1 0 24196 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1607194113
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607194113
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1607194113
transform 1 0 23644 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1607194113
transform 1 0 25116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_263
timestamp 1607194113
transform 1 0 25300 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_285
timestamp 1607194113
transform 1 0 27324 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_273
timestamp 1607194113
transform 1 0 26220 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_288
timestamp 1607194113
transform 1 0 27600 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_276
timestamp 1607194113
transform 1 0 26496 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607194113
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_297
timestamp 1607194113
transform 1 0 28428 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_300
timestamp 1607194113
transform 1 0 28704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607194113
transform -1 0 29256 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607194113
transform -1 0 29256 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_239
timestamp 1607194113
transform 1 0 23092 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__CLK
timestamp 1607194113
transform 1 0 23368 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1517_
timestamp 1607194113
transform 1 0 23552 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_263
timestamp 1607194113
transform 1 0 25300 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_276
timestamp 1607194113
transform 1 0 26496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B1
timestamp 1607194113
transform 1 0 26772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607194113
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1208_
timestamp 1607194113
transform 1 0 26956 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_310
timestamp 1607194113
transform 1 0 29624 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_303
timestamp 1607194113
transform 1 0 28980 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1607194113
transform 1 0 29440 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A2_N
timestamp 1607194113
transform 1 0 28796 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B2
timestamp 1607194113
transform 1 0 28612 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A1_N
timestamp 1607194113
transform 1 0 28428 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1607194113
transform 1 0 29164 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_322
timestamp 1607194113
transform 1 0 30728 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_349
timestamp 1607194113
transform 1 0 33212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_337
timestamp 1607194113
transform 1 0 32108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_334
timestamp 1607194113
transform 1 0 31832 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607194113
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_361
timestamp 1607194113
transform 1 0 34316 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_i
timestamp 1607194113
transform 1 0 35052 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_391
timestamp 1607194113
transform 1 0 37076 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_374
timestamp 1607194113
transform 1 0 35512 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_i_A
timestamp 1607194113
transform 1 0 35328 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1607194113
transform 1 0 36892 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1607194113
transform 1 0 36616 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_410
timestamp 1607194113
transform 1 0 38824 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_398
timestamp 1607194113
transform 1 0 37720 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607194113
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_430
timestamp 1607194113
transform 1 0 40664 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_422
timestamp 1607194113
transform 1 0 39928 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A1_N
timestamp 1607194113
transform 1 0 42504 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B1
timestamp 1607194113
transform 1 0 40848 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1214_
timestamp 1607194113
transform 1 0 41032 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_50_459
timestamp 1607194113
transform 1 0 43332 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_454
timestamp 1607194113
transform 1 0 42872 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A2_N
timestamp 1607194113
transform 1 0 42688 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607194113
transform 1 0 43240 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_245
timestamp 1607194113
transform 1 0 23644 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_241
timestamp 1607194113
transform 1 0 23276 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607194113
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1607194113
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_253
timestamp 1607194113
transform 1 0 24380 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1607194113
transform 1 0 25300 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0683_
timestamp 1607194113
transform 1 0 24472 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_51_277
timestamp 1607194113
transform 1 0 26588 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B1
timestamp 1607194113
transform 1 0 26772 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1209_
timestamp 1607194113
transform 1 0 26956 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_51_303
timestamp 1607194113
transform 1 0 28980 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A2_N
timestamp 1607194113
transform 1 0 28796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B2
timestamp 1607194113
transform 1 0 28612 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A1_N
timestamp 1607194113
transform 1 0 28428 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607194113
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1417_
timestamp 1607194113
transform 1 0 29256 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_327
timestamp 1607194113
transform 1 0 31188 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__CLK
timestamp 1607194113
transform 1 0 31004 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_351
timestamp 1607194113
transform 1 0 33396 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_339
timestamp 1607194113
transform 1 0 32292 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_367
timestamp 1607194113
transform 1 0 34868 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_363
timestamp 1607194113
transform 1 0 34500 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607194113
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1371_
timestamp 1607194113
transform 1 0 35604 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1607194113
transform 1 0 38364 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_398
timestamp 1607194113
transform 1 0 37720 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A
timestamp 1607194113
transform 1 0 37904 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A1_N
timestamp 1607194113
transform 1 0 37352 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B1
timestamp 1607194113
transform 1 0 37536 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1607194113
transform 1 0 38088 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_428
timestamp 1607194113
transform 1 0 40480 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_425
timestamp 1607194113
transform 1 0 40204 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_417
timestamp 1607194113
transform 1 0 39468 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607194113
transform 1 0 40388 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1413_
timestamp 1607194113
transform 1 0 41584 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1404_
timestamp 1607194113
transform 1 0 43332 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_52_252
timestamp 1607194113
transform 1 0 24288 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_247
timestamp 1607194113
transform 1 0 23828 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_239
timestamp 1607194113
transform 1 0 23092 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1607194113
transform 1 0 24012 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_272
timestamp 1607194113
transform 1 0 26128 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_264
timestamp 1607194113
transform 1 0 25392 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1607194113
transform 1 0 25024 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_288
timestamp 1607194113
transform 1 0 27600 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_276
timestamp 1607194113
transform 1 0 26496 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607194113
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_300
timestamp 1607194113
transform 1 0 28704 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1416_
timestamp 1607194113
transform 1 0 29072 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_52_325
timestamp 1607194113
transform 1 0 31004 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__CLK
timestamp 1607194113
transform 1 0 30820 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1607194113
transform 1 0 33212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1607194113
transform 1 0 32108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_333
timestamp 1607194113
transform 1 0 31740 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607194113
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_369
timestamp 1607194113
transform 1 0 35052 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_361
timestamp 1607194113
transform 1 0 34316 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B1
timestamp 1607194113
transform 1 0 35236 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_389
timestamp 1607194113
transform 1 0 36892 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A2_N
timestamp 1607194113
transform 1 0 36984 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1215_
timestamp 1607194113
transform 1 0 35420 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_52_396
timestamp 1607194113
transform 1 0 37536 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B2
timestamp 1607194113
transform 1 0 37168 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1_N
timestamp 1607194113
transform 1 0 37352 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607194113
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1277_
timestamp 1607194113
transform 1 0 37720 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_52_426
timestamp 1607194113
transform 1 0 40296 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_414
timestamp 1607194113
transform 1 0 39192 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A2_N
timestamp 1607194113
transform 1 0 40388 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B2
timestamp 1607194113
transform 1 0 40572 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B1
timestamp 1607194113
transform 1 0 40756 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_451
timestamp 1607194113
transform 1 0 42596 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A1_N
timestamp 1607194113
transform 1 0 42412 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1227_
timestamp 1607194113
transform 1 0 40940 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_464
timestamp 1607194113
transform 1 0 43792 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_457
timestamp 1607194113
transform 1 0 43148 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1607194113
transform 1 0 43608 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607194113
transform 1 0 43240 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1607194113
transform 1 0 43332 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_245
timestamp 1607194113
transform 1 0 23644 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B1
timestamp 1607194113
transform 1 0 23828 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607194113
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0684_
timestamp 1607194113
transform 1 0 24012 0 1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_53_263
timestamp 1607194113
transform 1 0 25300 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_287
timestamp 1607194113
transform 1 0 27508 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_275
timestamp 1607194113
transform 1 0 26404 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_311
timestamp 1607194113
transform 1 0 29716 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_299
timestamp 1607194113
transform 1 0 28612 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1607194113
transform 1 0 29532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607194113
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1607194113
transform 1 0 29256 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_323
timestamp 1607194113
transform 1 0 30820 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_347
timestamp 1607194113
transform 1 0 33028 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_335
timestamp 1607194113
transform 1 0 31924 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_367
timestamp 1607194113
transform 1 0 34868 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_365
timestamp 1607194113
transform 1 0 34684 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_359
timestamp 1607194113
transform 1 0 34132 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A
timestamp 1607194113
transform 1 0 35144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607194113
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_376
timestamp 1607194113
transform 1 0 35696 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1412_
timestamp 1607194113
transform 1 0 36432 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1607194113
transform 1 0 35328 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_403
timestamp 1607194113
transform 1 0 38180 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_428
timestamp 1607194113
transform 1 0 40480 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_415
timestamp 1607194113
transform 1 0 39284 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607194113
transform 1 0 40388 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_449
timestamp 1607194113
transform 1 0 42412 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_440
timestamp 1607194113
transform 1 0 41584 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A
timestamp 1607194113
transform 1 0 41860 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1210_
timestamp 1607194113
transform 1 0 42044 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_462
timestamp 1607194113
transform 1 0 43608 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1607194113
transform 1 0 43424 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1607194113
transform 1 0 43148 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_251
timestamp 1607194113
transform 1 0 24196 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_239
timestamp 1607194113
transform 1 0 23092 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_263
timestamp 1607194113
transform 1 0 25300 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_288
timestamp 1607194113
transform 1 0 27600 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_276
timestamp 1607194113
transform 1 0 26496 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607194113
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_312
timestamp 1607194113
transform 1 0 29808 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_300
timestamp 1607194113
transform 1 0 28704 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_324
timestamp 1607194113
transform 1 0 30912 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1607194113
transform 1 0 33212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_337
timestamp 1607194113
transform 1 0 32108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607194113
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_369
timestamp 1607194113
transform 1 0 35052 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_361
timestamp 1607194113
transform 1 0 34316 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A
timestamp 1607194113
transform 1 0 34500 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1607194113
transform 1 0 34684 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_381
timestamp 1607194113
transform 1 0 36156 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_410
timestamp 1607194113
transform 1 0 38824 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_398
timestamp 1607194113
transform 1 0 37720 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_393
timestamp 1607194113
transform 1 0 37260 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607194113
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_422
timestamp 1607194113
transform 1 0 39928 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A2_N
timestamp 1607194113
transform 1 0 40664 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A1_N
timestamp 1607194113
transform 1 0 42504 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B1
timestamp 1607194113
transform 1 0 40848 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1270_
timestamp 1607194113
transform 1 0 41032 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_454
timestamp 1607194113
transform 1 0 42872 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B2
timestamp 1607194113
transform 1 0 42688 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607194113
transform 1 0 43240 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1377_
timestamp 1607194113
transform 1 0 43332 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_243
timestamp 1607194113
transform 1 0 23460 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_245
timestamp 1607194113
transform 1 0 23644 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_243
timestamp 1607194113
transform 1 0 23460 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_237
timestamp 1607194113
transform 1 0 22908 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607194113
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_267
timestamp 1607194113
transform 1 0 25668 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_255
timestamp 1607194113
transform 1 0 24564 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_253
timestamp 1607194113
transform 1 0 24380 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B1
timestamp 1607194113
transform 1 0 24656 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1280_
timestamp 1607194113
transform 1 0 24840 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_288
timestamp 1607194113
transform 1 0 27600 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1607194113
transform 1 0 26496 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1607194113
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1607194113
transform 1 0 26680 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A2_N
timestamp 1607194113
transform 1 0 26496 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B2
timestamp 1607194113
transform 1 0 26312 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1607194113
transform 1 0 26864 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607194113
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1172_
timestamp 1607194113
transform 1 0 27048 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_300
timestamp 1607194113
transform 1 0 28704 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_298
timestamp 1607194113
transform 1 0 28520 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_304
timestamp 1607194113
transform 1 0 29072 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_304
timestamp 1607194113
transform 1 0 29072 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A2_N
timestamp 1607194113
transform 1 0 29164 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B2
timestamp 1607194113
transform 1 0 29348 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B1
timestamp 1607194113
transform 1 0 29532 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607194113
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_306
timestamp 1607194113
transform 1 0 29256 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1217_
timestamp 1607194113
transform 1 0 29716 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_56_329
timestamp 1607194113
transform 1 0 31372 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_330
timestamp 1607194113
transform 1 0 31464 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_318
timestamp 1607194113
transform 1 0 30360 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1_N
timestamp 1607194113
transform 1 0 31188 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B1
timestamp 1607194113
transform 1 0 31556 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1369_
timestamp 1607194113
transform 1 0 31556 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_56_335
timestamp 1607194113
transform 1 0 31924 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_352
timestamp 1607194113
transform 1 0 33488 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__CLK
timestamp 1607194113
transform 1 0 33304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B2
timestamp 1607194113
transform 1 0 31740 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607194113
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1279_
timestamp 1607194113
transform 1 0 32108 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_367
timestamp 1607194113
transform 1 0 34868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_355
timestamp 1607194113
transform 1 0 33764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_367
timestamp 1607194113
transform 1 0 34868 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_364
timestamp 1607194113
transform 1 0 34592 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A2_N
timestamp 1607194113
transform 1 0 33580 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A
timestamp 1607194113
transform 1 0 35052 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607194113
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1176_
timestamp 1607194113
transform 1 0 35236 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_391
timestamp 1607194113
transform 1 0 37076 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_379
timestamp 1607194113
transform 1 0 35972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_387
timestamp 1607194113
transform 1 0 36708 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_375
timestamp 1607194113
transform 1 0 35604 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A
timestamp 1607194113
transform 1 0 36156 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1206_
timestamp 1607194113
transform 1 0 36340 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_406
timestamp 1607194113
transform 1 0 38456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_398
timestamp 1607194113
transform 1 0 37720 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_411
timestamp 1607194113
transform 1 0 38916 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_399
timestamp 1607194113
transform 1 0 37812 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1607194113
transform 1 0 37904 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A
timestamp 1607194113
transform 1 0 37260 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607194113
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1276_
timestamp 1607194113
transform 1 0 37444 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1266_
timestamp 1607194113
transform 1 0 38088 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_430
timestamp 1607194113
transform 1 0 40664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_418
timestamp 1607194113
transform 1 0 39560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_428
timestamp 1607194113
transform 1 0 40480 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_423
timestamp 1607194113
transform 1 0 40020 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B2
timestamp 1607194113
transform 1 0 40572 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B1
timestamp 1607194113
transform 1 0 40756 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607194113
transform 1 0 40388 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_450
timestamp 1607194113
transform 1 0 42504 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_442
timestamp 1607194113
transform 1 0 41768 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A2_N
timestamp 1607194113
transform 1 0 42596 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1607194113
transform 1 0 41952 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A1_N
timestamp 1607194113
transform 1 0 42412 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1207_
timestamp 1607194113
transform 1 0 40940 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1203_
timestamp 1607194113
transform 1 0 42136 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_463
timestamp 1607194113
transform 1 0 43700 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_459
timestamp 1607194113
transform 1 0 43332 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_461
timestamp 1607194113
transform 1 0 43516 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_453
timestamp 1607194113
transform 1 0 42780 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1607194113
transform 1 0 42964 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607194113
transform 1 0 43240 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1418_
timestamp 1607194113
transform 1 0 43792 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1607194113
transform 1 0 43148 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_245
timestamp 1607194113
transform 1 0 23644 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1607194113
transform 1 0 23460 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607194113
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__CLK
timestamp 1607194113
transform 1 0 24748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1368_
timestamp 1607194113
transform 1 0 24932 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_289
timestamp 1607194113
transform 1 0 27692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_278
timestamp 1607194113
transform 1 0 26680 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1607194113
transform 1 0 27416 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_306
timestamp 1607194113
transform 1 0 29256 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1607194113
transform 1 0 28796 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607194113
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_318
timestamp 1607194113
transform 1 0 30360 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1410_
timestamp 1607194113
transform 1 0 30544 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_352
timestamp 1607194113
transform 1 0 33488 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_341
timestamp 1607194113
transform 1 0 32476 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__CLK
timestamp 1607194113
transform 1 0 32292 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A
timestamp 1607194113
transform 1 0 33304 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1607194113
transform 1 0 33028 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_367
timestamp 1607194113
transform 1 0 34868 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_364
timestamp 1607194113
transform 1 0 34592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607194113
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_387
timestamp 1607194113
transform 1 0 36708 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_379
timestamp 1607194113
transform 1 0 35972 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B2
timestamp 1607194113
transform 1 0 36892 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A2
timestamp 1607194113
transform 1 0 37076 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1607194113
transform 1 0 35420 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1607194113
transform 1 0 35604 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_407
timestamp 1607194113
transform 1 0 38548 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0931_
timestamp 1607194113
transform 1 0 37260 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_57_428
timestamp 1607194113
transform 1 0 40480 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_419
timestamp 1607194113
transform 1 0 39652 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607194113
transform 1 0 40388 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_440
timestamp 1607194113
transform 1 0 41584 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_464
timestamp 1607194113
transform 1 0 43792 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_452
timestamp 1607194113
transform 1 0 42688 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_252
timestamp 1607194113
transform 1 0 24288 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_240
timestamp 1607194113
transform 1 0 23184 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_267
timestamp 1607194113
transform 1 0 25668 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1607194113
transform 1 0 25392 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B2
timestamp 1607194113
transform 1 0 27968 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B1
timestamp 1607194113
transform 1 0 26220 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607194113
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1218_
timestamp 1607194113
transform 1 0 26496 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_308
timestamp 1607194113
transform 1 0 29440 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_296
timestamp 1607194113
transform 1 0 28336 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A2_N
timestamp 1607194113
transform 1 0 28152 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_332
timestamp 1607194113
transform 1 0 31648 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_320
timestamp 1607194113
transform 1 0 30544 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_352
timestamp 1607194113
transform 1 0 33488 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_340
timestamp 1607194113
transform 1 0 32384 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607194113
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1607194113
transform 1 0 32108 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_364
timestamp 1607194113
transform 1 0 34592 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_388
timestamp 1607194113
transform 1 0 36800 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_376
timestamp 1607194113
transform 1 0 35696 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B1
timestamp 1607194113
transform 1 0 36984 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_396
timestamp 1607194113
transform 1 0 37536 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A2_N
timestamp 1607194113
transform 1 0 37168 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B2
timestamp 1607194113
transform 1 0 37352 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607194113
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1202_
timestamp 1607194113
transform 1 0 37720 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_426
timestamp 1607194113
transform 1 0 40296 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_414
timestamp 1607194113
transform 1 0 39192 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_450
timestamp 1607194113
transform 1 0 42504 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_438
timestamp 1607194113
transform 1 0 41400 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_459
timestamp 1607194113
transform 1 0 43332 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607194113
transform 1 0 43240 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1607194113
transform 1 0 23644 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_242
timestamp 1607194113
transform 1 0 23368 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607194113
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_265
timestamp 1607194113
transform 1 0 25484 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_257
timestamp 1607194113
transform 1 0 24748 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1409_
timestamp 1607194113
transform 1 0 25760 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_289
timestamp 1607194113
transform 1 0 27692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__CLK
timestamp 1607194113
transform 1 0 27508 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1607194113
transform 1 0 29256 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1607194113
transform 1 0 28796 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607194113
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_330
timestamp 1607194113
transform 1 0 31464 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1607194113
transform 1 0 30360 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_342
timestamp 1607194113
transform 1 0 32568 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1607194113
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_354
timestamp 1607194113
transform 1 0 33672 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607194113
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_379
timestamp 1607194113
transform 1 0 35972 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B2
timestamp 1607194113
transform 1 0 36340 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1607194113
transform 1 0 36524 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0925_
timestamp 1607194113
transform 1 0 36708 0 1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_59_401
timestamp 1607194113
transform 1 0 37996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_428
timestamp 1607194113
transform 1 0 40480 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_426
timestamp 1607194113
transform 1 0 40296 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_420
timestamp 1607194113
transform 1 0 39744 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_413
timestamp 1607194113
transform 1 0 39100 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1607194113
transform 1 0 39560 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607194113
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1607194113
transform 1 0 39284 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_440
timestamp 1607194113
transform 1 0 41584 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_452
timestamp 1607194113
transform 1 0 42688 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B1
timestamp 1607194113
transform 1 0 42872 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1265_
timestamp 1607194113
transform 1 0 43056 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_245
timestamp 1607194113
transform 1 0 23644 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_269
timestamp 1607194113
transform 1 0 25852 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_257
timestamp 1607194113
transform 1 0 24748 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1607194113
transform 1 0 27968 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B2
timestamp 1607194113
transform 1 0 27784 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607194113
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0706_
timestamp 1607194113
transform 1 0 26496 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_60_306
timestamp 1607194113
transform 1 0 29256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1607194113
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_330
timestamp 1607194113
transform 1 0 31464 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_318
timestamp 1607194113
transform 1 0 30360 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_347
timestamp 1607194113
transform 1 0 33028 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_337
timestamp 1607194113
transform 1 0 32108 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A
timestamp 1607194113
transform 1 0 32844 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607194113
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1196_
timestamp 1607194113
transform 1 0 32476 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_371
timestamp 1607194113
transform 1 0 35236 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_359
timestamp 1607194113
transform 1 0 34132 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_389
timestamp 1607194113
transform 1 0 36892 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1607194113
transform 1 0 36340 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1199_
timestamp 1607194113
transform 1 0 36524 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_398
timestamp 1607194113
transform 1 0 37720 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1607194113
transform 1 0 38272 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607194113
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1421_
timestamp 1607194113
transform 1 0 38456 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_425
timestamp 1607194113
transform 1 0 40204 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_449
timestamp 1607194113
transform 1 0 42412 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_437
timestamp 1607194113
transform 1 0 41308 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_465
timestamp 1607194113
transform 1 0 43884 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_457
timestamp 1607194113
transform 1 0 43148 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1607194113
transform 1 0 43700 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607194113
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1262_
timestamp 1607194113
transform 1 0 43332 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_245
timestamp 1607194113
transform 1 0 23644 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1607194113
transform 1 0 23644 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1607194113
transform 1 0 23460 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_239
timestamp 1607194113
transform 1 0 23092 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1607194113
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1607194113
transform 1 0 25852 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_257
timestamp 1607194113
transform 1 0 24748 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_257
timestamp 1607194113
transform 1 0 24748 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0804_
timestamp 1607194113
transform 1 0 25852 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_285
timestamp 1607194113
transform 1 0 27324 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_287
timestamp 1607194113
transform 1 0 27508 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1607194113
transform 1 0 27324 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1607194113
transform 1 0 27140 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1607194113
transform 1 0 26220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1607194113
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0707_
timestamp 1607194113
transform 1 0 26496 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1607194113
transform 1 0 29532 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_297
timestamp 1607194113
transform 1 0 28428 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_312
timestamp 1607194113
transform 1 0 29808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_299
timestamp 1607194113
transform 1 0 28612 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1607194113
transform 1 0 29624 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1607194113
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1236_
timestamp 1607194113
transform 1 0 29256 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1607194113
transform 1 0 30636 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_324
timestamp 1607194113
transform 1 0 30912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_341
timestamp 1607194113
transform 1 0 32476 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_337
timestamp 1607194113
transform 1 0 32108 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_333
timestamp 1607194113
transform 1 0 31740 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B1
timestamp 1607194113
transform 1 0 33488 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1607194113
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0799_
timestamp 1607194113
transform 1 0 32568 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0701_
timestamp 1607194113
transform 1 0 32016 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_362
timestamp 1607194113
transform 1 0 34408 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1607194113
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_360
timestamp 1607194113
transform 1 0 34224 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A2_N
timestamp 1607194113
transform 1 0 34040 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B2
timestamp 1607194113
transform 1 0 33856 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A2_N
timestamp 1607194113
transform 1 0 34224 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B2
timestamp 1607194113
transform 1 0 34040 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A1_N
timestamp 1607194113
transform 1 0 33672 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1607194113
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_386
timestamp 1607194113
transform 1 0 36616 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_374
timestamp 1607194113
transform 1 0 35512 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_391
timestamp 1607194113
transform 1 0 37076 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1607194113
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_394
timestamp 1607194113
transform 1 0 37352 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_403
timestamp 1607194113
transform 1 0 38180 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B1
timestamp 1607194113
transform 1 0 37444 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1607194113
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1197_
timestamp 1607194113
transform 1 0 37720 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_428
timestamp 1607194113
transform 1 0 40480 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_416
timestamp 1607194113
transform 1 0 39376 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_428
timestamp 1607194113
transform 1 0 40480 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_415
timestamp 1607194113
transform 1 0 39284 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1_N
timestamp 1607194113
transform 1 0 39192 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1607194113
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_440
timestamp 1607194113
transform 1 0 41584 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_440
timestamp 1607194113
transform 1 0 41584 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_459
timestamp 1607194113
transform 1 0 43332 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_452
timestamp 1607194113
transform 1 0 42688 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_452
timestamp 1607194113
transform 1 0 42688 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B1
timestamp 1607194113
transform 1 0 42780 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1607194113
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1263_
timestamp 1607194113
transform 1 0 42964 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1607194113
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_242
timestamp 1607194113
transform 1 0 23368 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_234
timestamp 1607194113
transform 1 0 22632 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1607194113
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_265
timestamp 1607194113
transform 1 0 25484 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_257
timestamp 1607194113
transform 1 0 24748 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A
timestamp 1607194113
transform 1 0 25668 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B
timestamp 1607194113
transform 1 0 25852 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0805_
timestamp 1607194113
transform 1 0 26036 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_292
timestamp 1607194113
transform 1 0 27968 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_280
timestamp 1607194113
transform 1 0 26864 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1607194113
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_304
timestamp 1607194113
transform 1 0 29072 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1607194113
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_330
timestamp 1607194113
transform 1 0 31464 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1607194113
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_351
timestamp 1607194113
transform 1 0 33396 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__B1
timestamp 1607194113
transform 1 0 31740 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1198_
timestamp 1607194113
transform 1 0 31924 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1607194113
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_363
timestamp 1607194113
transform 1 0 34500 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1607194113
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1607194113
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B2
timestamp 1607194113
transform 1 0 37076 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_411
timestamp 1607194113
transform 1 0 38916 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B1
timestamp 1607194113
transform 1 0 37260 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1200_
timestamp 1607194113
transform 1 0 37444 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_428
timestamp 1607194113
transform 1 0 40480 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_423
timestamp 1607194113
transform 1 0 40020 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1607194113
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_440
timestamp 1607194113
transform 1 0 41584 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B1
timestamp 1607194113
transform 1 0 41768 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1260_
timestamp 1607194113
transform 1 0 41952 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_462
timestamp 1607194113
transform 1 0 43608 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A1_N
timestamp 1607194113
transform 1 0 43424 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_247
timestamp 1607194113
transform 1 0 23828 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_235
timestamp 1607194113
transform 1 0 22724 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1607194113
transform 1 0 26036 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_259
timestamp 1607194113
transform 1 0 24932 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1607194113
transform 1 0 26496 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1607194113
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1389_
timestamp 1607194113
transform 1 0 26864 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_301
timestamp 1607194113
transform 1 0 28796 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__CLK
timestamp 1607194113
transform 1 0 28612 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_325
timestamp 1607194113
transform 1 0 31004 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_313
timestamp 1607194113
transform 1 0 29900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_333
timestamp 1607194113
transform 1 0 31740 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__B1
timestamp 1607194113
transform 1 0 31832 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1607194113
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1261_
timestamp 1607194113
transform 1 0 32108 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1607194113
transform 1 0 34684 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_355
timestamp 1607194113
transform 1 0 33764 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A
timestamp 1607194113
transform 1 0 34132 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A1_N
timestamp 1607194113
transform 1 0 33580 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1259_
timestamp 1607194113
transform 1 0 34316 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_389
timestamp 1607194113
transform 1 0 36892 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1607194113
transform 1 0 35788 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_398
timestamp 1607194113
transform 1 0 37720 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__CLK
timestamp 1607194113
transform 1 0 38272 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1607194113
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1423_
timestamp 1607194113
transform 1 0 38456 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_64_425
timestamp 1607194113
transform 1 0 40204 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_448
timestamp 1607194113
transform 1 0 42320 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_436
timestamp 1607194113
transform 1 0 41216 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1607194113
transform 1 0 40940 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_459
timestamp 1607194113
transform 1 0 43332 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_456
timestamp 1607194113
transform 1 0 43056 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1607194113
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_252
timestamp 1607194113
transform 1 0 24288 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_245
timestamp 1607194113
transform 1 0 23644 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_242
timestamp 1607194113
transform 1 0 23368 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1607194113
transform 1 0 23736 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1607194113
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1252_
timestamp 1607194113
transform 1 0 23920 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_260
timestamp 1607194113
transform 1 0 25024 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__B1
timestamp 1607194113
transform 1 0 25300 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1253_
timestamp 1607194113
transform 1 0 25484 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_283
timestamp 1607194113
transform 1 0 27140 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1_N
timestamp 1607194113
transform 1 0 26956 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_306
timestamp 1607194113
transform 1 0 29256 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_303
timestamp 1607194113
transform 1 0 28980 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_295
timestamp 1607194113
transform 1 0 28244 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1607194113
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_330
timestamp 1607194113
transform 1 0 31464 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1607194113
transform 1 0 30360 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_349
timestamp 1607194113
transform 1 0 33212 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_342
timestamp 1607194113
transform 1 0 32568 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk_i
timestamp 1607194113
transform 1 0 32936 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_370
timestamp 1607194113
transform 1 0 35144 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_364
timestamp 1607194113
transform 1 0 34592 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_356
timestamp 1607194113
transform 1 0 33856 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1607194113
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1607194113
transform 1 0 34868 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1607194113
transform 1 0 33580 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_382
timestamp 1607194113
transform 1 0 36248 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_406
timestamp 1607194113
transform 1 0 38456 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_394
timestamp 1607194113
transform 1 0 37352 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0815_
timestamp 1607194113
transform 1 0 38824 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_428
timestamp 1607194113
transform 1 0 40480 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_419
timestamp 1607194113
transform 1 0 39652 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1607194113
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_440
timestamp 1607194113
transform 1 0 41584 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_464
timestamp 1607194113
transform 1 0 43792 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_452
timestamp 1607194113
transform 1 0 42688 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_252
timestamp 1607194113
transform 1 0 24288 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_240
timestamp 1607194113
transform 1 0 23184 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_272
timestamp 1607194113
transform 1 0 26128 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_264
timestamp 1607194113
transform 1 0 25392 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_276
timestamp 1607194113
transform 1 0 26496 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B1
timestamp 1607194113
transform 1 0 26220 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1607194113
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1190_
timestamp 1607194113
transform 1 0 26588 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_307
timestamp 1607194113
transform 1 0 29348 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_295
timestamp 1607194113
transform 1 0 28244 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A1_N
timestamp 1607194113
transform 1 0 28060 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_331
timestamp 1607194113
transform 1 0 31556 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_319
timestamp 1607194113
transform 1 0 30452 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_345
timestamp 1607194113
transform 1 0 32844 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_337
timestamp 1607194113
transform 1 0 32108 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_335
timestamp 1607194113
transform 1 0 31924 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__CLK
timestamp 1607194113
transform 1 0 32936 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1607194113
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1383_
timestamp 1607194113
transform 1 0 33120 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_367
timestamp 1607194113
transform 1 0 34868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_391
timestamp 1607194113
transform 1 0 37076 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_379
timestamp 1607194113
transform 1 0 35972 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_406
timestamp 1607194113
transform 1 0 38456 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_398
timestamp 1607194113
transform 1 0 37720 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1607194113
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0797_
timestamp 1607194113
transform 1 0 38732 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_66_429
timestamp 1607194113
transform 1 0 40572 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B2
timestamp 1607194113
transform 1 0 40388 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__C
timestamp 1607194113
transform 1 0 40756 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A2_N
timestamp 1607194113
transform 1 0 40204 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_442
timestamp 1607194113
transform 1 0 41768 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0720_
timestamp 1607194113
transform 1 0 40940 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_459
timestamp 1607194113
transform 1 0 43332 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_454
timestamp 1607194113
transform 1 0 42872 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1607194113
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_248
timestamp 1607194113
transform 1 0 23920 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1607194113
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1607194113
transform 1 0 23644 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_272
timestamp 1607194113
transform 1 0 26128 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_260
timestamp 1607194113
transform 1 0 25024 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_284
timestamp 1607194113
transform 1 0 27232 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1189_
timestamp 1607194113
transform 1 0 27968 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_306
timestamp 1607194113
transform 1 0 29256 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_304
timestamp 1607194113
transform 1 0 29072 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_298
timestamp 1607194113
transform 1 0 28520 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1607194113
transform 1 0 28336 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1607194113
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_330
timestamp 1607194113
transform 1 0 31464 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_318
timestamp 1607194113
transform 1 0 30360 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_342
timestamp 1607194113
transform 1 0 32568 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1607194113
transform 1 0 34868 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_354
timestamp 1607194113
transform 1 0 33672 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1607194113
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_388
timestamp 1607194113
transform 1 0 36800 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_379
timestamp 1607194113
transform 1 0 35972 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_i_A
timestamp 1607194113
transform 1 0 36616 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_i
timestamp 1607194113
transform 1 0 36340 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_400
timestamp 1607194113
transform 1 0 37904 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_428
timestamp 1607194113
transform 1 0 40480 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_424
timestamp 1607194113
transform 1 0 40112 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_412
timestamp 1607194113
transform 1 0 39008 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1607194113
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_440
timestamp 1607194113
transform 1 0 41584 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_464
timestamp 1607194113
transform 1 0 43792 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_452
timestamp 1607194113
transform 1 0 42688 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_248
timestamp 1607194113
transform 1 0 23920 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_243
timestamp 1607194113
transform 1 0 23460 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_237
timestamp 1607194113
transform 1 0 22908 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_248
timestamp 1607194113
transform 1 0 23920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_236
timestamp 1607194113
transform 1 0 22816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1_N
timestamp 1607194113
transform 1 0 22632 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1607194113
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1607194113
transform 1 0 23644 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_272
timestamp 1607194113
transform 1 0 26128 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_260
timestamp 1607194113
transform 1 0 25024 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_272
timestamp 1607194113
transform 1 0 26128 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_260
timestamp 1607194113
transform 1 0 25024 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_284
timestamp 1607194113
transform 1 0 27232 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_288
timestamp 1607194113
transform 1 0 27600 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_276
timestamp 1607194113
transform 1 0 26496 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1607194113
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1430_
timestamp 1607194113
transform 1 0 27968 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_312
timestamp 1607194113
transform 1 0 29808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_304
timestamp 1607194113
transform 1 0 29072 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_296
timestamp 1607194113
transform 1 0 28336 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__CLK
timestamp 1607194113
transform 1 0 29716 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1607194113
transform 1 0 29624 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1607194113
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1182_
timestamp 1607194113
transform 1 0 29256 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_324
timestamp 1607194113
transform 1 0 30912 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_325
timestamp 1607194113
transform 1 0 31004 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_313
timestamp 1607194113
transform 1 0 29900 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_348
timestamp 1607194113
transform 1 0 33120 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_336
timestamp 1607194113
transform 1 0 32016 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_337
timestamp 1607194113
transform 1 0 32108 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1607194113
transform 1 0 31740 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1607194113
transform 1 0 32844 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1607194113
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1424_
timestamp 1607194113
transform 1 0 33028 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1607194113
transform 1 0 34868 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_360
timestamp 1607194113
transform 1 0 34224 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_366
timestamp 1607194113
transform 1 0 34776 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1607194113
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_391
timestamp 1607194113
transform 1 0 37076 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1607194113
transform 1 0 35972 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_390
timestamp 1607194113
transform 1 0 36984 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_378
timestamp 1607194113
transform 1 0 35880 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_403
timestamp 1607194113
transform 1 0 38180 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_398
timestamp 1607194113
transform 1 0 37720 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_396
timestamp 1607194113
transform 1 0 37536 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1607194113
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0698_
timestamp 1607194113
transform 1 0 38824 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_415
timestamp 1607194113
transform 1 0 39284 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_430
timestamp 1607194113
transform 1 0 40664 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B2
timestamp 1607194113
transform 1 0 40480 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A2_N
timestamp 1607194113
transform 1 0 40296 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1607194113
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0814_
timestamp 1607194113
transform 1 0 40480 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1607194113
transform 1 0 42412 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_437
timestamp 1607194113
transform 1 0 41308 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_442
timestamp 1607194113
transform 1 0 41768 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1607194113
transform 1 0 43516 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_459
timestamp 1607194113
transform 1 0 43332 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_454
timestamp 1607194113
transform 1 0 42872 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B1
timestamp 1607194113
transform 1 0 43884 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1607194113
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_247
timestamp 1607194113
transform 1 0 23828 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_271
timestamp 1607194113
transform 1 0 26036 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_259
timestamp 1607194113
transform 1 0 24932 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_285
timestamp 1607194113
transform 1 0 27324 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1607194113
transform 1 0 27140 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1607194113
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0703_
timestamp 1607194113
transform 1 0 26496 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_70_297
timestamp 1607194113
transform 1 0 28428 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B1
timestamp 1607194113
transform 1 0 29164 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1184_
timestamp 1607194113
transform 1 0 29348 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_70_325
timestamp 1607194113
transform 1 0 31004 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1_N
timestamp 1607194113
transform 1 0 30820 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_345
timestamp 1607194113
transform 1 0 32844 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_337
timestamp 1607194113
transform 1 0 32108 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_333
timestamp 1607194113
transform 1 0 31740 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__CLK
timestamp 1607194113
transform 1 0 32936 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1607194113
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1393_
timestamp 1607194113
transform 1 0 33120 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_367
timestamp 1607194113
transform 1 0 34868 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_391
timestamp 1607194113
transform 1 0 37076 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_379
timestamp 1607194113
transform 1 0 35972 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_398
timestamp 1607194113
transform 1 0 37720 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B1
timestamp 1607194113
transform 1 0 38456 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1607194113
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0711_
timestamp 1607194113
transform 1 0 38640 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_428
timestamp 1607194113
transform 1 0 40480 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B2
timestamp 1607194113
transform 1 0 40296 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A2_N
timestamp 1607194113
transform 1 0 40112 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_441
timestamp 1607194113
transform 1 0 41676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0719_
timestamp 1607194113
transform 1 0 40848 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_459
timestamp 1607194113
transform 1 0 43332 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_457
timestamp 1607194113
transform 1 0 43148 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_453
timestamp 1607194113
transform 1 0 42780 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1607194113
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_245
timestamp 1607194113
transform 1 0 23644 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_241
timestamp 1607194113
transform 1 0 23276 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__B1
timestamp 1607194113
transform 1 0 23736 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1607194113
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1183_
timestamp 1607194113
transform 1 0 23920 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_264
timestamp 1607194113
transform 1 0 25392 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1435_
timestamp 1607194113
transform 1 0 26128 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__CLK
timestamp 1607194113
transform 1 0 27876 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_306
timestamp 1607194113
transform 1 0 29256 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1607194113
transform 1 0 28060 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B1
timestamp 1607194113
transform 1 0 29440 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1607194113
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1247_
timestamp 1607194113
transform 1 0 29624 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_328
timestamp 1607194113
transform 1 0 31280 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1_N
timestamp 1607194113
transform 1 0 31096 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_352
timestamp 1607194113
transform 1 0 33488 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_340
timestamp 1607194113
transform 1 0 32384 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1607194113
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_364
timestamp 1607194113
transform 1 0 34592 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1607194113
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_391
timestamp 1607194113
transform 1 0 37076 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1607194113
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_399
timestamp 1607194113
transform 1 0 37812 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1607194113
transform 1 0 37996 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0807_
timestamp 1607194113
transform 1 0 38180 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_71_423
timestamp 1607194113
transform 1 0 40020 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B2
timestamp 1607194113
transform 1 0 39836 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1_N
timestamp 1607194113
transform 1 0 40204 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2_N
timestamp 1607194113
transform 1 0 39652 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1607194113
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0811_
timestamp 1607194113
transform 1 0 40480 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_446
timestamp 1607194113
transform 1 0 42136 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1607194113
transform 1 0 41952 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_458
timestamp 1607194113
transform 1 0 43240 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_251
timestamp 1607194113
transform 1 0 24196 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_239
timestamp 1607194113
transform 1 0 23092 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_263
timestamp 1607194113
transform 1 0 25300 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_285
timestamp 1607194113
transform 1 0 27324 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1607194113
transform 1 0 27692 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1607194113
transform 1 0 27140 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1607194113
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0802_
timestamp 1607194113
transform 1 0 26496 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1607194113
transform 1 0 27876 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_306
timestamp 1607194113
transform 1 0 29256 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_294
timestamp 1607194113
transform 1 0 28152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A
timestamp 1607194113
transform 1 0 29808 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1245_
timestamp 1607194113
transform 1 0 29440 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_326
timestamp 1607194113
transform 1 0 31096 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_314
timestamp 1607194113
transform 1 0 29992 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_345
timestamp 1607194113
transform 1 0 32844 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_337
timestamp 1607194113
transform 1 0 32108 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_334
timestamp 1607194113
transform 1 0 31832 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1607194113
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1434_
timestamp 1607194113
transform 1 0 33120 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_369
timestamp 1607194113
transform 1 0 35052 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1607194113
transform 1 0 34868 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_381
timestamp 1607194113
transform 1 0 36156 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_410
timestamp 1607194113
transform 1 0 38824 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_398
timestamp 1607194113
transform 1 0 37720 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_393
timestamp 1607194113
transform 1 0 37260 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1607194113
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1_N
timestamp 1607194113
transform 1 0 39100 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B2
timestamp 1607194113
transform 1 0 40756 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0716_
timestamp 1607194113
transform 1 0 39284 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1607194113
transform 1 0 42044 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1607194113
transform 1 0 40940 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_459
timestamp 1607194113
transform 1 0 43332 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_457
timestamp 1607194113
transform 1 0 43148 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1607194113
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_245
timestamp 1607194113
transform 1 0 23644 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_240
timestamp 1607194113
transform 1 0 23184 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B1
timestamp 1607194113
transform 1 0 24012 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1607194113
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1246_
timestamp 1607194113
transform 1 0 24196 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_267
timestamp 1607194113
transform 1 0 25668 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_285
timestamp 1607194113
transform 1 0 27324 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1607194113
transform 1 0 26772 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1607194113
transform 1 0 27140 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1607194113
transform 1 0 26864 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_306
timestamp 1607194113
transform 1 0 29256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_297
timestamp 1607194113
transform 1 0 28428 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1607194113
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_330
timestamp 1607194113
transform 1 0 31464 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_318
timestamp 1607194113
transform 1 0 30360 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A
timestamp 1607194113
transform 1 0 30912 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1173_
timestamp 1607194113
transform 1 0 31096 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_342
timestamp 1607194113
transform 1 0 32568 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1607194113
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_354
timestamp 1607194113
transform 1 0 33672 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1607194113
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_391
timestamp 1607194113
transform 1 0 37076 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1607194113
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_403
timestamp 1607194113
transform 1 0 38180 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_428
timestamp 1607194113
transform 1 0 40480 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_415
timestamp 1607194113
transform 1 0 39284 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1607194113
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_440
timestamp 1607194113
transform 1 0 41584 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_464
timestamp 1607194113
transform 1 0 43792 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_452
timestamp 1607194113
transform 1 0 42688 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_248
timestamp 1607194113
transform 1 0 23920 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_236
timestamp 1607194113
transform 1 0 22816 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_245
timestamp 1607194113
transform 1 0 23644 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1607194113
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1607194113
transform 1 0 23644 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_262
timestamp 1607194113
transform 1 0 25208 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_256
timestamp 1607194113
transform 1 0 24656 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_269
timestamp 1607194113
transform 1 0 25852 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_257
timestamp 1607194113
transform 1 0 24748 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1607194113
transform 1 0 25760 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1607194113
transform 1 0 24748 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1394_
timestamp 1607194113
transform 1 0 25944 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1607194113
transform 1 0 24932 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_289
timestamp 1607194113
transform 1 0 27692 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_288
timestamp 1607194113
transform 1 0 27600 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_276
timestamp 1607194113
transform 1 0 26496 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1607194113
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_306
timestamp 1607194113
transform 1 0 29256 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_301
timestamp 1607194113
transform 1 0 28796 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_312
timestamp 1607194113
transform 1 0 29808 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_300
timestamp 1607194113
transform 1 0 28704 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1607194113
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_330
timestamp 1607194113
transform 1 0 31464 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_318
timestamp 1607194113
transform 1 0 30360 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_328
timestamp 1607194113
transform 1 0 31280 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_320
timestamp 1607194113
transform 1 0 30544 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A
timestamp 1607194113
transform 1 0 30728 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1237_
timestamp 1607194113
transform 1 0 30912 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_337
timestamp 1607194113
transform 1 0 32108 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B1
timestamp 1607194113
transform 1 0 32200 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1607194113
transform 1 0 32476 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1607194113
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1239_
timestamp 1607194113
transform 1 0 32660 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1175_
timestamp 1607194113
transform 1 0 32384 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_75_367
timestamp 1607194113
transform 1 0 34868 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_358
timestamp 1607194113
transform 1 0 34040 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_361
timestamp 1607194113
transform 1 0 34316 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1_N
timestamp 1607194113
transform 1 0 34132 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1_N
timestamp 1607194113
transform 1 0 33856 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1607194113
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_385
timestamp 1607194113
transform 1 0 36524 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_373
timestamp 1607194113
transform 1 0 35420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1398_
timestamp 1607194113
transform 1 0 35420 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_75_394
timestamp 1607194113
transform 1 0 37352 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_410
timestamp 1607194113
transform 1 0 38824 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_398
timestamp 1607194113
transform 1 0 37720 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__CLK
timestamp 1607194113
transform 1 0 37720 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__CLK
timestamp 1607194113
transform 1 0 37168 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1607194113
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1439_
timestamp 1607194113
transform 1 0 37904 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1607194113
transform 1 0 38916 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_428
timestamp 1607194113
transform 1 0 40480 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_419
timestamp 1607194113
transform 1 0 39652 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_426
timestamp 1607194113
transform 1 0 40296 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_414
timestamp 1607194113
transform 1 0 39192 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1607194113
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_440
timestamp 1607194113
transform 1 0 41584 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_450
timestamp 1607194113
transform 1 0 42504 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_438
timestamp 1607194113
transform 1 0 41400 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_464
timestamp 1607194113
transform 1 0 43792 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_452
timestamp 1607194113
transform 1 0 42688 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_459
timestamp 1607194113
transform 1 0 43332 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1607194113
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_245
timestamp 1607194113
transform 1 0 23644 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_269
timestamp 1607194113
transform 1 0 25852 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_257
timestamp 1607194113
transform 1 0 24748 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_276
timestamp 1607194113
transform 1 0 26496 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1607194113
transform 1 0 26404 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0872_
timestamp 1607194113
transform 1 0 27232 0 -1 44064
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_76_302
timestamp 1607194113
transform 1 0 28888 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B1
timestamp 1607194113
transform 1 0 28704 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A1
timestamp 1607194113
transform 1 0 28520 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_326
timestamp 1607194113
transform 1 0 31096 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_314
timestamp 1607194113
transform 1 0 29992 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_337
timestamp 1607194113
transform 1 0 32108 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B1
timestamp 1607194113
transform 1 0 31832 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1607194113
transform 1 0 32016 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1174_
timestamp 1607194113
transform 1 0 32200 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_368
timestamp 1607194113
transform 1 0 34960 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_356
timestamp 1607194113
transform 1 0 33856 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A1_N
timestamp 1607194113
transform 1 0 33672 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_391
timestamp 1607194113
transform 1 0 37076 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_380
timestamp 1607194113
transform 1 0 36064 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk_i
timestamp 1607194113
transform 1 0 36800 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_409
timestamp 1607194113
transform 1 0 38732 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_398
timestamp 1607194113
transform 1 0 37720 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1607194113
transform 1 0 37628 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1607194113
transform 1 0 38456 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__CLK
timestamp 1607194113
transform 1 0 39468 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1440_
timestamp 1607194113
transform 1 0 39652 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_76_449
timestamp 1607194113
transform 1 0 42412 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_438
timestamp 1607194113
transform 1 0 41400 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1607194113
transform 1 0 42136 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_459
timestamp 1607194113
transform 1 0 43332 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_457
timestamp 1607194113
transform 1 0 43148 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1607194113
transform 1 0 43240 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_245
timestamp 1607194113
transform 1 0 23644 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_236
timestamp 1607194113
transform 1 0 22816 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1607194113
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_269
timestamp 1607194113
transform 1 0 25852 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_257
timestamp 1607194113
transform 1 0 24748 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1607194113
transform 1 0 26956 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0870_
timestamp 1607194113
transform 1 0 27140 0 1 44064
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_77_306
timestamp 1607194113
transform 1 0 29256 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_301
timestamp 1607194113
transform 1 0 28796 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1607194113
transform 1 0 28612 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1607194113
transform 1 0 28428 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1607194113
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_330
timestamp 1607194113
transform 1 0 31464 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_318
timestamp 1607194113
transform 1 0 30360 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_338
timestamp 1607194113
transform 1 0 32200 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B1
timestamp 1607194113
transform 1 0 32292 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1238_
timestamp 1607194113
transform 1 0 32476 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_367
timestamp 1607194113
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_365
timestamp 1607194113
transform 1 0 34684 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_359
timestamp 1607194113
transform 1 0 34132 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A1_N
timestamp 1607194113
transform 1 0 33948 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1607194113
transform 1 0 34776 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_391
timestamp 1607194113
transform 1 0 37076 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_379
timestamp 1607194113
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_403
timestamp 1607194113
transform 1 0 38180 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_428
timestamp 1607194113
transform 1 0 40480 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_415
timestamp 1607194113
transform 1 0 39284 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1607194113
transform 1 0 40388 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_441
timestamp 1607194113
transform 1 0 41676 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_436
timestamp 1607194113
transform 1 0 41216 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1607194113
transform 1 0 41400 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_465
timestamp 1607194113
transform 1 0 43884 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_453
timestamp 1607194113
transform 1 0 42780 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_247
timestamp 1607194113
transform 1 0 23828 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_239
timestamp 1607194113
transform 1 0 23092 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A
timestamp 1607194113
transform 1 0 24012 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1241_
timestamp 1607194113
transform 1 0 24196 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_267
timestamp 1607194113
transform 1 0 25668 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_255
timestamp 1607194113
transform 1 0 24564 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_288
timestamp 1607194113
transform 1 0 27600 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_276
timestamp 1607194113
transform 1 0 26496 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1607194113
transform 1 0 26404 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1607194113
transform 1 0 29532 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_300
timestamp 1607194113
transform 1 0 28704 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1607194113
transform 1 0 29348 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1177_
timestamp 1607194113
transform 1 0 28980 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1607194113
transform 1 0 30636 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_349
timestamp 1607194113
transform 1 0 33212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_337
timestamp 1607194113
transform 1 0 32108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_333
timestamp 1607194113
transform 1 0 31740 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1607194113
transform 1 0 32016 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_361
timestamp 1607194113
transform 1 0 34316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_385
timestamp 1607194113
transform 1 0 36524 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_373
timestamp 1607194113
transform 1 0 35420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_406
timestamp 1607194113
transform 1 0 38456 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_398
timestamp 1607194113
transform 1 0 37720 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__CLK
timestamp 1607194113
transform 1 0 38732 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1607194113
transform 1 0 37628 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1399_
timestamp 1607194113
transform 1 0 38916 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_78_430
timestamp 1607194113
transform 1 0 40664 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_442
timestamp 1607194113
transform 1 0 41768 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_459
timestamp 1607194113
transform 1 0 43332 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_454
timestamp 1607194113
transform 1 0 42872 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1607194113
transform 1 0 43240 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_245
timestamp 1607194113
transform 1 0 23644 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1607194113
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_269
timestamp 1607194113
transform 1 0 25852 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_257
timestamp 1607194113
transform 1 0 24748 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1607194113
transform 1 0 26956 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_306
timestamp 1607194113
transform 1 0 29256 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1607194113
transform 1 0 28060 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1607194113
transform 1 0 29164 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_318
timestamp 1607194113
transform 1 0 30360 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B2
timestamp 1607194113
transform 1 0 30636 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B1
timestamp 1607194113
transform 1 0 30820 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1242_
timestamp 1607194113
transform 1 0 31004 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_343
timestamp 1607194113
transform 1 0 32660 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1_N
timestamp 1607194113
transform 1 0 32476 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1607194113
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_363
timestamp 1607194113
transform 1 0 34500 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_355
timestamp 1607194113
transform 1 0 33764 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1607194113
transform 1 0 34776 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_391
timestamp 1607194113
transform 1 0 37076 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1607194113
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_403
timestamp 1607194113
transform 1 0 38180 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_428
timestamp 1607194113
transform 1 0 40480 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_415
timestamp 1607194113
transform 1 0 39284 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1607194113
transform 1 0 40388 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_440
timestamp 1607194113
transform 1 0 41584 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_464
timestamp 1607194113
transform 1 0 43792 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_452
timestamp 1607194113
transform 1 0 42688 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_478
timestamp 1607194113
transform 1 0 45080 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_470
timestamp 1607194113
transform 1 0 44344 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1607194113
transform 1 0 45264 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk_i
timestamp 1607194113
transform 1 0 44068 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 45448 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_50_502
timestamp 1607194113
transform 1 0 47288 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_520
timestamp 1607194113
transform 1 0 48944 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_513
timestamp 1607194113
transform 1 0 48300 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_i_A
timestamp 1607194113
transform 1 0 47840 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_i
timestamp 1607194113
transform 1 0 48024 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607194113
transform 1 0 48852 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_544
timestamp 1607194113
transform 1 0 51152 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_532
timestamp 1607194113
transform 1 0 50048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A2_N
timestamp 1607194113
transform 1 0 51336 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B2
timestamp 1607194113
transform 1 0 51520 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_570
timestamp 1607194113
transform 1 0 53544 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A1_N
timestamp 1607194113
transform 1 0 53360 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B1
timestamp 1607194113
transform 1 0 51704 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1211_
timestamp 1607194113
transform 1 0 51888 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1607194113
transform 1 0 54556 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_578
timestamp 1607194113
transform 1 0 54280 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_i_A
timestamp 1607194113
transform 1 0 55108 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_i
timestamp 1607194113
transform 1 0 55292 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607194113
transform 1 0 54464 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_600
timestamp 1607194113
transform 1 0 56304 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_592
timestamp 1607194113
transform 1 0 55568 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A2_N
timestamp 1607194113
transform 1 0 56396 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B2
timestamp 1607194113
transform 1 0 56580 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B1
timestamp 1607194113
transform 1 0 56764 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1226_
timestamp 1607194113
transform 1 0 56948 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_50_625
timestamp 1607194113
transform 1 0 58604 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[8]
timestamp 1607194113
transform 1 0 59156 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[3]
timestamp 1607194113
transform 1 0 58788 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[1]
timestamp 1607194113
transform 1 0 58972 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A1_N
timestamp 1607194113
transform 1 0 58420 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_inp_i
timestamp 1607194113
transform 1 0 59524 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[7]
timestamp 1607194113
transform 1 0 59340 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[6]
timestamp 1607194113
transform 1 0 59892 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[4]
timestamp 1607194113
transform 1 0 59708 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607194113
transform 1 0 60076 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1405_
timestamp 1607194113
transform 1 0 60168 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_663
timestamp 1607194113
transform 1 0 62100 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__CLK
timestamp 1607194113
transform 1 0 61916 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_687
timestamp 1607194113
transform 1 0 64308 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_675
timestamp 1607194113
transform 1 0 63204 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_699
timestamp 1607194113
transform 1 0 65412 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_486
timestamp 1607194113
transform 1 0 45816 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_478
timestamp 1607194113
transform 1 0 45080 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_497
timestamp 1607194113
transform 1 0 46828 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_489
timestamp 1607194113
transform 1 0 46092 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607194113
transform 1 0 46000 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1411_
timestamp 1607194113
transform 1 0 46920 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_519
timestamp 1607194113
transform 1 0 48852 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__CLK
timestamp 1607194113
transform 1 0 48668 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_543
timestamp 1607194113
transform 1 0 51060 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_531
timestamp 1607194113
transform 1 0 49956 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607194113
transform 1 0 51612 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_558
timestamp 1607194113
transform 1 0 52440 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_550
timestamp 1607194113
transform 1 0 51704 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__CLK
timestamp 1607194113
transform 1 0 52532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1415_
timestamp 1607194113
transform 1 0 52716 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_580
timestamp 1607194113
transform 1 0 54464 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_611
timestamp 1607194113
transform 1 0 57316 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_604
timestamp 1607194113
transform 1 0 56672 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_592
timestamp 1607194113
transform 1 0 55568 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607194113
transform 1 0 57224 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__CLK
timestamp 1607194113
transform 1 0 59156 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1374_
timestamp 1607194113
transform 1 0 57408 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_51_639
timestamp 1607194113
transform 1 0 59892 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_633
timestamp 1607194113
transform 1 0 59340 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1607194113
transform 1 0 59984 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[2]
timestamp 1607194113
transform 1 0 59708 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[0]
timestamp 1607194113
transform 1 0 59524 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1_N
timestamp 1607194113
transform 1 0 60168 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0760_
timestamp 1607194113
transform 1 0 60352 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_672
timestamp 1607194113
transform 1 0 62928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_670
timestamp 1607194113
transform 1 0 62744 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_664
timestamp 1607194113
transform 1 0 62192 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2_N
timestamp 1607194113
transform 1 0 62008 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B2
timestamp 1607194113
transform 1 0 61824 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607194113
transform 1 0 62836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_684
timestamp 1607194113
transform 1 0 64032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_696
timestamp 1607194113
transform 1 0 65136 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_476
timestamp 1607194113
transform 1 0 44896 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_506
timestamp 1607194113
transform 1 0 47656 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B1
timestamp 1607194113
transform 1 0 46000 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1216_
timestamp 1607194113
transform 1 0 46184 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_52_514
timestamp 1607194113
transform 1 0 48392 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__CLK
timestamp 1607194113
transform 1 0 48668 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607194113
transform 1 0 48852 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1370_
timestamp 1607194113
transform 1 0 48944 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_52_539
timestamp 1607194113
transform 1 0 50692 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_563
timestamp 1607194113
transform 1 0 52900 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_551
timestamp 1607194113
transform 1 0 51796 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_584
timestamp 1607194113
transform 1 0 54832 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_579
timestamp 1607194113
transform 1 0 54372 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_575
timestamp 1607194113
transform 1 0 54004 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607194113
transform 1 0 54464 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1607194113
transform 1 0 54556 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_596
timestamp 1607194113
transform 1 0 55936 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A2_N
timestamp 1607194113
transform 1 0 56120 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B2
timestamp 1607194113
transform 1 0 56304 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B1
timestamp 1607194113
transform 1 0 56488 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1273_
timestamp 1607194113
transform 1 0 56672 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_620
timestamp 1607194113
transform 1 0 58144 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1607194113
transform 1 0 59156 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1607194113
transform 1 0 58880 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_642
timestamp 1607194113
transform 1 0 60168 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_633
timestamp 1607194113
transform 1 0 59340 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1_N
timestamp 1607194113
transform 1 0 60720 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1607194113
transform 1 0 60904 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607194113
transform 1 0 60076 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0740_
timestamp 1607194113
transform 1 0 61088 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_672
timestamp 1607194113
transform 1 0 62928 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B2
timestamp 1607194113
transform 1 0 62744 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2_N
timestamp 1607194113
transform 1 0 62560 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_684
timestamp 1607194113
transform 1 0 64032 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_696
timestamp 1607194113
transform 1 0 65136 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_486
timestamp 1607194113
transform 1 0 45816 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_474
timestamp 1607194113
transform 1 0 44712 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_493
timestamp 1607194113
transform 1 0 46460 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_489
timestamp 1607194113
transform 1 0 46092 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A2_N
timestamp 1607194113
transform 1 0 46552 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B2
timestamp 1607194113
transform 1 0 46736 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B1
timestamp 1607194113
transform 1 0 46920 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607194113
transform 1 0 46000 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1278_
timestamp 1607194113
transform 1 0 47104 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_528
timestamp 1607194113
transform 1 0 49680 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_516
timestamp 1607194113
transform 1 0 48576 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_548
timestamp 1607194113
transform 1 0 51520 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_540
timestamp 1607194113
transform 1 0 50784 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607194113
transform 1 0 51612 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_568
timestamp 1607194113
transform 1 0 53360 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_562
timestamp 1607194113
transform 1 0 52808 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_550
timestamp 1607194113
transform 1 0 51704 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0783_
timestamp 1607194113
transform 1 0 53452 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_589
timestamp 1607194113
transform 1 0 55292 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A2_N
timestamp 1607194113
transform 1 0 55108 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B2
timestamp 1607194113
transform 1 0 54924 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_611
timestamp 1607194113
transform 1 0 57316 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_609
timestamp 1607194113
transform 1 0 57132 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_601
timestamp 1607194113
transform 1 0 56396 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607194113
transform 1 0 57224 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_632
timestamp 1607194113
transform 1 0 59248 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_623
timestamp 1607194113
transform 1 0 58420 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1607194113
transform 1 0 58972 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_640
timestamp 1607194113
transform 1 0 59984 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A1_N
timestamp 1607194113
transform 1 0 60260 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1607194113
transform 1 0 60444 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0736_
timestamp 1607194113
transform 1 0 60628 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_53_667
timestamp 1607194113
transform 1 0 62468 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B2
timestamp 1607194113
transform 1 0 62284 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2_N
timestamp 1607194113
transform 1 0 62100 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607194113
transform 1 0 62836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0741_
timestamp 1607194113
transform 1 0 62928 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_53_693
timestamp 1607194113
transform 1 0 64860 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_681
timestamp 1607194113
transform 1 0 63756 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_478
timestamp 1607194113
transform 1 0 45080 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_502
timestamp 1607194113
transform 1 0 47288 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_490
timestamp 1607194113
transform 1 0 46184 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_520
timestamp 1607194113
transform 1 0 48944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_518
timestamp 1607194113
transform 1 0 48760 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_514
timestamp 1607194113
transform 1 0 48392 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607194113
transform 1 0 48852 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_544
timestamp 1607194113
transform 1 0 51152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_532
timestamp 1607194113
transform 1 0 50048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_570
timestamp 1607194113
transform 1 0 53544 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_564
timestamp 1607194113
transform 1 0 52992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_556
timestamp 1607194113
transform 1 0 52256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1607194113
transform 1 0 53084 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1607194113
transform 1 0 53268 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_586
timestamp 1607194113
transform 1 0 55016 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_578
timestamp 1607194113
transform 1 0 54280 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1607194113
transform 1 0 54832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607194113
transform 1 0 54464 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1607194113
transform 1 0 54556 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_610
timestamp 1607194113
transform 1 0 57224 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_598
timestamp 1607194113
transform 1 0 56120 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_622
timestamp 1607194113
transform 1 0 58328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_642
timestamp 1607194113
transform 1 0 60168 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_640
timestamp 1607194113
transform 1 0 59984 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_634
timestamp 1607194113
transform 1 0 59432 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607194113
transform 1 0 60076 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_666
timestamp 1607194113
transform 1 0 62376 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_654
timestamp 1607194113
transform 1 0 61272 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_690
timestamp 1607194113
transform 1 0 64584 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_678
timestamp 1607194113
transform 1 0 63480 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_483
timestamp 1607194113
transform 1 0 45540 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_485
timestamp 1607194113
transform 1 0 45724 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1607194113
transform 1 0 44620 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_469
timestamp 1607194113
transform 1 0 44252 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1607194113
transform 1 0 44344 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_506
timestamp 1607194113
transform 1 0 47656 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_494
timestamp 1607194113
transform 1 0 46552 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_501
timestamp 1607194113
transform 1 0 47196 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_489
timestamp 1607194113
transform 1 0 46092 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607194113
transform 1 0 46000 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1607194113
transform 1 0 46276 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_518
timestamp 1607194113
transform 1 0 48760 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_524
timestamp 1607194113
transform 1 0 49312 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_512
timestamp 1607194113
transform 1 0 48208 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B2
timestamp 1607194113
transform 1 0 48944 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1607194113
transform 1 0 49128 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk_i
timestamp 1607194113
transform 1 0 47932 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607194113
transform 1 0 48852 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0935_
timestamp 1607194113
transform 1 0 49312 0 -1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_56_538
timestamp 1607194113
transform 1 0 50600 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_548
timestamp 1607194113
transform 1 0 51520 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_536
timestamp 1607194113
transform 1 0 50416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607194113
transform 1 0 51612 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_562
timestamp 1607194113
transform 1 0 52808 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_550
timestamp 1607194113
transform 1 0 51704 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_562
timestamp 1607194113
transform 1 0 52808 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1607194113
transform 1 0 51704 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0854_
timestamp 1607194113
transform 1 0 53084 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_581
timestamp 1607194113
transform 1 0 54556 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_574
timestamp 1607194113
transform 1 0 53912 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_587
timestamp 1607194113
transform 1 0 55108 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2_N
timestamp 1607194113
transform 1 0 54924 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B1
timestamp 1607194113
transform 1 0 54740 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B2
timestamp 1607194113
transform 1 0 54556 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607194113
transform 1 0 54464 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_605
timestamp 1607194113
transform 1 0 56764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_593
timestamp 1607194113
transform 1 0 55660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_611
timestamp 1607194113
transform 1 0 57316 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_607
timestamp 1607194113
transform 1 0 56948 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_599
timestamp 1607194113
transform 1 0 56212 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607194113
transform 1 0 57224 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_629
timestamp 1607194113
transform 1 0 58972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_617
timestamp 1607194113
transform 1 0 57868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_623
timestamp 1607194113
transform 1 0 58420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_642
timestamp 1607194113
transform 1 0 60168 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_643
timestamp 1607194113
transform 1 0 60260 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_635
timestamp 1607194113
transform 1 0 59524 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1607194113
transform 1 0 60352 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607194113
transform 1 0 60076 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0759_
timestamp 1607194113
transform 1 0 60536 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_654
timestamp 1607194113
transform 1 0 61272 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_672
timestamp 1607194113
transform 1 0 62928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_668
timestamp 1607194113
transform 1 0 62560 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B2
timestamp 1607194113
transform 1 0 62376 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2_N
timestamp 1607194113
transform 1 0 62192 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1_N
timestamp 1607194113
transform 1 0 62008 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A1_N
timestamp 1607194113
transform 1 0 61640 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607194113
transform 1 0 62836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0732_
timestamp 1607194113
transform 1 0 61824 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_694
timestamp 1607194113
transform 1 0 64952 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_682
timestamp 1607194113
transform 1 0 63848 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_684
timestamp 1607194113
transform 1 0 64032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B2
timestamp 1607194113
transform 1 0 63664 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B1
timestamp 1607194113
transform 1 0 63480 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A2_N
timestamp 1607194113
transform 1 0 63296 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_696
timestamp 1607194113
transform 1 0 65136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_476
timestamp 1607194113
transform 1 0 44896 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_501
timestamp 1607194113
transform 1 0 47196 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_489
timestamp 1607194113
transform 1 0 46092 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607194113
transform 1 0 46000 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_513
timestamp 1607194113
transform 1 0 48300 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A2_N
timestamp 1607194113
transform 1 0 48852 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B2
timestamp 1607194113
transform 1 0 49036 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B1
timestamp 1607194113
transform 1 0 49220 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1205_
timestamp 1607194113
transform 1 0 49404 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_541
timestamp 1607194113
transform 1 0 50876 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B2
timestamp 1607194113
transform 1 0 51244 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1607194113
transform 1 0 51428 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607194113
transform 1 0 51612 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_550
timestamp 1607194113
transform 1 0 51704 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A2_N
timestamp 1607194113
transform 1 0 53452 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1
timestamp 1607194113
transform 1 0 53268 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1607194113
transform 1 0 53084 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0933_
timestamp 1607194113
transform 1 0 51796 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B2
timestamp 1607194113
transform 1 0 53636 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A1_N
timestamp 1607194113
transform 1 0 55476 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B1
timestamp 1607194113
transform 1 0 53820 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1204_
timestamp 1607194113
transform 1 0 54004 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_57_609
timestamp 1607194113
transform 1 0 57132 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_593
timestamp 1607194113
transform 1 0 55660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A1_N
timestamp 1607194113
transform 1 0 56948 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1607194113
transform 1 0 56764 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607194113
transform 1 0 57224 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0763_
timestamp 1607194113
transform 1 0 57316 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_631
timestamp 1607194113
transform 1 0 59156 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B2
timestamp 1607194113
transform 1 0 58972 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A2_N
timestamp 1607194113
transform 1 0 58788 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_643
timestamp 1607194113
transform 1 0 60260 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0764_
timestamp 1607194113
transform 1 0 60628 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_672
timestamp 1607194113
transform 1 0 62928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_668
timestamp 1607194113
transform 1 0 62560 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_656
timestamp 1607194113
transform 1 0 61456 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607194113
transform 1 0 62836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_684
timestamp 1607194113
transform 1 0 64032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_696
timestamp 1607194113
transform 1 0 65136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_467
timestamp 1607194113
transform 1 0 44068 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1380_
timestamp 1607194113
transform 1 0 44344 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1607194113
transform 1 0 47196 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1607194113
transform 1 0 46092 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_513
timestamp 1607194113
transform 1 0 48300 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A2_N
timestamp 1607194113
transform 1 0 48944 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B2
timestamp 1607194113
transform 1 0 49128 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B1
timestamp 1607194113
transform 1 0 48668 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607194113
transform 1 0 48852 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1268_
timestamp 1607194113
transform 1 0 49312 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_540
timestamp 1607194113
transform 1 0 50784 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_564
timestamp 1607194113
transform 1 0 52992 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_552
timestamp 1607194113
transform 1 0 51888 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_579
timestamp 1607194113
transform 1 0 54372 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_572
timestamp 1607194113
transform 1 0 53728 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A2_N
timestamp 1607194113
transform 1 0 54004 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B2
timestamp 1607194113
transform 1 0 54188 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607194113
transform 1 0 54464 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1267_
timestamp 1607194113
transform 1 0 54556 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_599
timestamp 1607194113
transform 1 0 56212 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1_N
timestamp 1607194113
transform 1 0 56580 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B1
timestamp 1607194113
transform 1 0 56764 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1_N
timestamp 1607194113
transform 1 0 56028 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0840_
timestamp 1607194113
transform 1 0 56948 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_627
timestamp 1607194113
transform 1 0 58788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B2
timestamp 1607194113
transform 1 0 58604 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A2_N
timestamp 1607194113
transform 1 0 58420 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_642
timestamp 1607194113
transform 1 0 60168 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_639
timestamp 1607194113
transform 1 0 59892 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607194113
transform 1 0 60076 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_670
timestamp 1607194113
transform 1 0 62744 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_666
timestamp 1607194113
transform 1 0 62376 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_654
timestamp 1607194113
transform 1 0 61272 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__CLK
timestamp 1607194113
transform 1 0 62836 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1379_
timestamp 1607194113
transform 1 0 63020 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_58_692
timestamp 1607194113
transform 1 0 64768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_476
timestamp 1607194113
transform 1 0 44896 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A2_N
timestamp 1607194113
transform 1 0 44712 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B2
timestamp 1607194113
transform 1 0 44528 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_501
timestamp 1607194113
transform 1 0 47196 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_489
timestamp 1607194113
transform 1 0 46092 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607194113
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_525
timestamp 1607194113
transform 1 0 49404 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_513
timestamp 1607194113
transform 1 0 48300 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_545
timestamp 1607194113
transform 1 0 51244 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_537
timestamp 1607194113
transform 1 0 50508 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1607194113
transform 1 0 51428 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607194113
transform 1 0 51612 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_568
timestamp 1607194113
transform 1 0 53360 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B2
timestamp 1607194113
transform 1 0 51704 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B1
timestamp 1607194113
transform 1 0 53176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0927_
timestamp 1607194113
transform 1 0 51888 0 1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_59_581
timestamp 1607194113
transform 1 0 54556 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_576
timestamp 1607194113
transform 1 0 54096 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B1
timestamp 1607194113
transform 1 0 54372 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_611
timestamp 1607194113
transform 1 0 57316 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_609
timestamp 1607194113
transform 1 0 57132 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_605
timestamp 1607194113
transform 1 0 56764 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_593
timestamp 1607194113
transform 1 0 55660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607194113
transform 1 0 57224 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_631
timestamp 1607194113
transform 1 0 59156 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_623
timestamp 1607194113
transform 1 0 58420 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__CLK
timestamp 1607194113
transform 1 0 61180 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1515_
timestamp 1607194113
transform 1 0 59432 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_59_670
timestamp 1607194113
transform 1 0 62744 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_663
timestamp 1607194113
transform 1 0 62100 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_655
timestamp 1607194113
transform 1 0 61364 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A1_N
timestamp 1607194113
transform 1 0 62560 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1607194113
transform 1 0 62376 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607194113
transform 1 0 62836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0758_
timestamp 1607194113
transform 1 0 62928 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_692
timestamp 1607194113
transform 1 0 64768 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2_N
timestamp 1607194113
transform 1 0 64584 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B2
timestamp 1607194113
transform 1 0 64400 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_476
timestamp 1607194113
transform 1 0 44896 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1607194113
transform 1 0 44712 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1607194113
transform 1 0 44436 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_500
timestamp 1607194113
transform 1 0 47104 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_488
timestamp 1607194113
transform 1 0 46000 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_520
timestamp 1607194113
transform 1 0 48944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_518
timestamp 1607194113
transform 1 0 48760 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_512
timestamp 1607194113
transform 1 0 48208 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607194113
transform 1 0 48852 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_544
timestamp 1607194113
transform 1 0 51152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_532
timestamp 1607194113
transform 1 0 50048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_568
timestamp 1607194113
transform 1 0 53360 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_556
timestamp 1607194113
transform 1 0 52256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_589
timestamp 1607194113
transform 1 0 55292 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_581
timestamp 1607194113
transform 1 0 54556 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A2_N
timestamp 1607194113
transform 1 0 55476 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607194113
transform 1 0 54464 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B2
timestamp 1607194113
transform 1 0 55660 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B1
timestamp 1607194113
transform 1 0 55844 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1264_
timestamp 1607194113
transform 1 0 56028 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_627
timestamp 1607194113
transform 1 0 58788 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_615
timestamp 1607194113
transform 1 0 57684 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A1_N
timestamp 1607194113
transform 1 0 57500 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_642
timestamp 1607194113
transform 1 0 60168 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_639
timestamp 1607194113
transform 1 0 59892 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1607194113
transform 1 0 60076 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_666
timestamp 1607194113
transform 1 0 62376 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_654
timestamp 1607194113
transform 1 0 61272 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_690
timestamp 1607194113
transform 1 0 64584 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_678
timestamp 1607194113
transform 1 0 63480 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_471
timestamp 1607194113
transform 1 0 44436 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_485
timestamp 1607194113
transform 1 0 45724 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1607194113
transform 1 0 44620 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B2
timestamp 1607194113
transform 1 0 44436 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1425_
timestamp 1607194113
transform 1 0 45172 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_61_495
timestamp 1607194113
transform 1 0 46644 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_489
timestamp 1607194113
transform 1 0 46092 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1607194113
transform 1 0 46736 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1607194113
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_506
timestamp 1607194113
transform 1 0 47656 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_500
timestamp 1607194113
transform 1 0 47104 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1607194113
transform 1 0 46920 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1607194113
transform 1 0 47748 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1607194113
transform 1 0 46920 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_501
timestamp 1607194113
transform 1 0 47196 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_520
timestamp 1607194113
transform 1 0 48944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_518
timestamp 1607194113
transform 1 0 48760 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_512
timestamp 1607194113
transform 1 0 48208 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_525
timestamp 1607194113
transform 1 0 49404 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_513
timestamp 1607194113
transform 1 0 48300 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1607194113
transform 1 0 48024 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1607194113
transform 1 0 48852 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_532
timestamp 1607194113
transform 1 0 50048 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_537
timestamp 1607194113
transform 1 0 50508 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__CLK
timestamp 1607194113
transform 1 0 50600 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1607194113
transform 1 0 51612 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1378_
timestamp 1607194113
transform 1 0 50784 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_559
timestamp 1607194113
transform 1 0 52532 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_567
timestamp 1607194113
transform 1 0 53268 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_555
timestamp 1607194113
transform 1 0 52164 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_550
timestamp 1607194113
transform 1 0 51704 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1607194113
transform 1 0 51888 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_581
timestamp 1607194113
transform 1 0 54556 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_579
timestamp 1607194113
transform 1 0 54372 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_571
timestamp 1607194113
transform 1 0 53636 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_591
timestamp 1607194113
transform 1 0 55476 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_579
timestamp 1607194113
transform 1 0 54372 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1607194113
transform 1 0 54464 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_599
timestamp 1607194113
transform 1 0 56212 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_593
timestamp 1607194113
transform 1 0 55660 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A2_N
timestamp 1607194113
transform 1 0 56304 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_609
timestamp 1607194113
transform 1 0 57132 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_603
timestamp 1607194113
transform 1 0 56580 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B2
timestamp 1607194113
transform 1 0 56488 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B1
timestamp 1607194113
transform 1 0 56672 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1607194113
transform 1 0 57224 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_611
timestamp 1607194113
transform 1 0 57316 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1201_
timestamp 1607194113
transform 1 0 56856 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_622
timestamp 1607194113
transform 1 0 58328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1422_
timestamp 1607194113
transform 1 0 58420 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_642
timestamp 1607194113
transform 1 0 60168 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_640
timestamp 1607194113
transform 1 0 59984 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_634
timestamp 1607194113
transform 1 0 59432 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_644
timestamp 1607194113
transform 1 0 60352 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__CLK
timestamp 1607194113
transform 1 0 60168 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1607194113
transform 1 0 60076 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_666
timestamp 1607194113
transform 1 0 62376 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_654
timestamp 1607194113
transform 1 0 61272 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_672
timestamp 1607194113
transform 1 0 62928 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_668
timestamp 1607194113
transform 1 0 62560 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_656
timestamp 1607194113
transform 1 0 61456 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1607194113
transform 1 0 62836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1607194113
transform 1 0 63112 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1607194113
transform 1 0 63112 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_689
timestamp 1607194113
transform 1 0 64492 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_677
timestamp 1607194113
transform 1 0 63388 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_689
timestamp 1607194113
transform 1 0 64492 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_677
timestamp 1607194113
transform 1 0 63388 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_486
timestamp 1607194113
transform 1 0 45816 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_474
timestamp 1607194113
transform 1 0 44712 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_489
timestamp 1607194113
transform 1 0 46092 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1607194113
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1384_
timestamp 1607194113
transform 1 0 46644 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_63_528
timestamp 1607194113
transform 1 0 49680 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_516
timestamp 1607194113
transform 1 0 48576 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__CLK
timestamp 1607194113
transform 1 0 48392 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_541
timestamp 1607194113
transform 1 0 50876 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_536
timestamp 1607194113
transform 1 0 50416 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1607194113
transform 1 0 51428 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1607194113
transform 1 0 51612 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1607194113
transform 1 0 50600 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_569
timestamp 1607194113
transform 1 0 53452 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1419_
timestamp 1607194113
transform 1 0 51704 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_581
timestamp 1607194113
transform 1 0 54556 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_611
timestamp 1607194113
transform 1 0 57316 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_609
timestamp 1607194113
transform 1 0 57132 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_605
timestamp 1607194113
transform 1 0 56764 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_593
timestamp 1607194113
transform 1 0 55660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1607194113
transform 1 0 57224 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_619
timestamp 1607194113
transform 1 0 58052 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1381_
timestamp 1607194113
transform 1 0 58144 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1607194113
transform 1 0 61180 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1607194113
transform 1 0 60076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__CLK
timestamp 1607194113
transform 1 0 59892 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_672
timestamp 1607194113
transform 1 0 62928 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1607194113
transform 1 0 62284 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1607194113
transform 1 0 62836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_680
timestamp 1607194113
transform 1 0 63664 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0691_
timestamp 1607194113
transform 1 0 63940 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A2
timestamp 1607194113
transform 1 0 65412 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B2
timestamp 1607194113
transform 1 0 65228 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_i_A
timestamp 1607194113
transform 1 0 44436 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_i
timestamp 1607194113
transform 1 0 44620 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1382_
timestamp 1607194113
transform 1 0 44896 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_497
timestamp 1607194113
transform 1 0 46828 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1607194113
transform 1 0 46644 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_520
timestamp 1607194113
transform 1 0 48944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_517
timestamp 1607194113
transform 1 0 48668 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_509
timestamp 1607194113
transform 1 0 47932 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1607194113
transform 1 0 48852 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_544
timestamp 1607194113
transform 1 0 51152 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_532
timestamp 1607194113
transform 1 0 50048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_550
timestamp 1607194113
transform 1 0 51704 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B2
timestamp 1607194113
transform 1 0 53452 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2_N
timestamp 1607194113
transform 1 0 53268 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0746_
timestamp 1607194113
transform 1 0 51796 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_581
timestamp 1607194113
transform 1 0 54556 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_579
timestamp 1607194113
transform 1 0 54372 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_571
timestamp 1607194113
transform 1 0 53636 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1607194113
transform 1 0 54464 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_605
timestamp 1607194113
transform 1 0 56764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_593
timestamp 1607194113
transform 1 0 55660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_629
timestamp 1607194113
transform 1 0 58972 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_617
timestamp 1607194113
transform 1 0 57868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_645
timestamp 1607194113
transform 1 0 60444 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1607194113
transform 1 0 60076 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1607194113
transform 1 0 60168 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_669
timestamp 1607194113
transform 1 0 62652 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_657
timestamp 1607194113
transform 1 0 61548 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_677
timestamp 1607194113
transform 1 0 63388 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B1
timestamp 1607194113
transform 1 0 63480 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B2
timestamp 1607194113
transform 1 0 64952 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0792_
timestamp 1607194113
transform 1 0 63664 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_64_698
timestamp 1607194113
transform 1 0 65320 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A2
timestamp 1607194113
transform 1 0 65136 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_476
timestamp 1607194113
transform 1 0 44896 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_504
timestamp 1607194113
transform 1 0 47472 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_492
timestamp 1607194113
transform 1 0 46368 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1607194113
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1607194113
transform 1 0 46092 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_528
timestamp 1607194113
transform 1 0 49680 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_516
timestamp 1607194113
transform 1 0 48576 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_548
timestamp 1607194113
transform 1 0 51520 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_540
timestamp 1607194113
transform 1 0 50784 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1607194113
transform 1 0 51612 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_570
timestamp 1607194113
transform 1 0 53544 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B2
timestamp 1607194113
transform 1 0 53360 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A2_N
timestamp 1607194113
transform 1 0 53176 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0828_
timestamp 1607194113
transform 1 0 51704 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_582
timestamp 1607194113
transform 1 0 54648 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_611
timestamp 1607194113
transform 1 0 57316 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_606
timestamp 1607194113
transform 1 0 56856 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_594
timestamp 1607194113
transform 1 0 55752 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1607194113
transform 1 0 57224 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1607194113
transform 1 0 58420 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0858_
timestamp 1607194113
transform 1 0 58604 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_653
timestamp 1607194113
transform 1 0 61180 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_646
timestamp 1607194113
transform 1 0 60536 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_634
timestamp 1607194113
transform 1 0 59432 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk_i
timestamp 1607194113
transform 1 0 60904 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_672
timestamp 1607194113
transform 1 0 62928 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1607194113
transform 1 0 62284 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1607194113
transform 1 0 62836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_681
timestamp 1607194113
transform 1 0 63756 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1607194113
transform 1 0 63296 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1
timestamp 1607194113
transform 1 0 64124 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1607194113
transform 1 0 64308 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0790_
timestamp 1607194113
transform 1 0 64492 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1607194113
transform 1 0 63480 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_483
timestamp 1607194113
transform 1 0 45540 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_471
timestamp 1607194113
transform 1 0 44436 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_507
timestamp 1607194113
transform 1 0 47748 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_495
timestamp 1607194113
transform 1 0 46644 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_520
timestamp 1607194113
transform 1 0 48944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1607194113
transform 1 0 48852 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_544
timestamp 1607194113
transform 1 0 51152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_532
timestamp 1607194113
transform 1 0 50048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_567
timestamp 1607194113
transform 1 0 53268 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_556
timestamp 1607194113
transform 1 0 52256 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0756_
timestamp 1607194113
transform 1 0 52440 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_581
timestamp 1607194113
transform 1 0 54556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_579
timestamp 1607194113
transform 1 0 54372 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1607194113
transform 1 0 54464 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_605
timestamp 1607194113
transform 1 0 56764 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_593
timestamp 1607194113
transform 1 0 55660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_629
timestamp 1607194113
transform 1 0 58972 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_617
timestamp 1607194113
transform 1 0 57868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_651
timestamp 1607194113
transform 1 0 60996 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_637
timestamp 1607194113
transform 1 0 59708 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B
timestamp 1607194113
transform 1 0 59892 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1607194113
transform 1 0 60076 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0787_
timestamp 1607194113
transform 1 0 60168 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_663
timestamp 1607194113
transform 1 0 62100 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_691
timestamp 1607194113
transform 1 0 64676 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_683
timestamp 1607194113
transform 1 0 63940 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_675
timestamp 1607194113
transform 1 0 63204 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1607194113
transform 1 0 64216 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1607194113
transform 1 0 64400 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_i_A
timestamp 1607194113
transform 1 0 65228 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_i
timestamp 1607194113
transform 1 0 65412 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_476
timestamp 1607194113
transform 1 0 44896 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A1_N
timestamp 1607194113
transform 1 0 47748 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B1
timestamp 1607194113
transform 1 0 46092 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1607194113
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0755_
timestamp 1607194113
transform 1 0 46276 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_525
timestamp 1607194113
transform 1 0 49404 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_513
timestamp 1607194113
transform 1 0 48300 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B2
timestamp 1607194113
transform 1 0 48116 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A2_N
timestamp 1607194113
transform 1 0 47932 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_545
timestamp 1607194113
transform 1 0 51244 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_537
timestamp 1607194113
transform 1 0 50508 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1_N
timestamp 1607194113
transform 1 0 51428 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1607194113
transform 1 0 51612 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_550
timestamp 1607194113
transform 1 0 51704 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B2
timestamp 1607194113
transform 1 0 53452 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1607194113
transform 1 0 51796 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0749_
timestamp 1607194113
transform 1 0 51980 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_586
timestamp 1607194113
transform 1 0 55016 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_573
timestamp 1607194113
transform 1 0 53820 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2_N
timestamp 1607194113
transform 1 0 53636 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0835_
timestamp 1607194113
transform 1 0 54188 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_67_611
timestamp 1607194113
transform 1 0 57316 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_598
timestamp 1607194113
transform 1 0 56120 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1607194113
transform 1 0 57224 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_619
timestamp 1607194113
transform 1 0 58052 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A1_N
timestamp 1607194113
transform 1 0 58144 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1607194113
transform 1 0 58328 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0817_
timestamp 1607194113
transform 1 0 58512 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_67_642
timestamp 1607194113
transform 1 0 60168 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A1
timestamp 1607194113
transform 1 0 60536 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2_N
timestamp 1607194113
transform 1 0 59984 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0827_
timestamp 1607194113
transform 1 0 60720 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_67_672
timestamp 1607194113
transform 1 0 62928 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_670
timestamp 1607194113
transform 1 0 62744 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_664
timestamp 1607194113
transform 1 0 62192 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__C1
timestamp 1607194113
transform 1 0 62008 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1607194113
transform 1 0 62836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_684
timestamp 1607194113
transform 1 0 64032 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A1
timestamp 1607194113
transform 1 0 64308 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0688_
timestamp 1607194113
transform 1 0 64492 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_69_485
timestamp 1607194113
transform 1 0 45724 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1607194113
transform 1 0 44620 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B2
timestamp 1607194113
transform 1 0 45724 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A1_N
timestamp 1607194113
transform 1 0 44068 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0714_
timestamp 1607194113
transform 1 0 44252 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_69_489
timestamp 1607194113
transform 1 0 46092 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1607194113
transform 1 0 46092 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A2_N
timestamp 1607194113
transform 1 0 45908 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1607194113
transform 1 0 46828 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B1
timestamp 1607194113
transform 1 0 46276 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1_N
timestamp 1607194113
transform 1 0 47012 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1607194113
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0855_
timestamp 1607194113
transform 1 0 47196 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0834_
timestamp 1607194113
transform 1 0 46460 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_521
timestamp 1607194113
transform 1 0 49036 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_520
timestamp 1607194113
transform 1 0 48944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_515
timestamp 1607194113
transform 1 0 48484 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B2
timestamp 1607194113
transform 1 0 48300 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2_N
timestamp 1607194113
transform 1 0 48852 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A2_N
timestamp 1607194113
transform 1 0 48116 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A1_N
timestamp 1607194113
transform 1 0 47932 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B2
timestamp 1607194113
transform 1 0 48668 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1607194113
transform 1 0 48852 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_545
timestamp 1607194113
transform 1 0 51244 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_533
timestamp 1607194113
transform 1 0 50140 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_544
timestamp 1607194113
transform 1 0 51152 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_532
timestamp 1607194113
transform 1 0 50048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1607194113
transform 1 0 51612 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_562
timestamp 1607194113
transform 1 0 52808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_550
timestamp 1607194113
transform 1 0 51704 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A1_N
timestamp 1607194113
transform 1 0 51704 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B1
timestamp 1607194113
transform 1 0 51888 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B2
timestamp 1607194113
transform 1 0 53544 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0830_
timestamp 1607194113
transform 1 0 52072 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_585
timestamp 1607194113
transform 1 0 54924 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_590
timestamp 1607194113
transform 1 0 55384 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_574
timestamp 1607194113
transform 1 0 53912 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__B
timestamp 1607194113
transform 1 0 54740 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A2_N
timestamp 1607194113
transform 1 0 53728 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1607194113
transform 1 0 54464 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0857_
timestamp 1607194113
transform 1 0 53912 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0786_
timestamp 1607194113
transform 1 0 54556 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_69_611
timestamp 1607194113
transform 1 0 57316 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_609
timestamp 1607194113
transform 1 0 57132 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_597
timestamp 1607194113
transform 1 0 56028 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_602
timestamp 1607194113
transform 1 0 56488 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1607194113
transform 1 0 57224 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_621
timestamp 1607194113
transform 1 0 58236 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1607194113
transform 1 0 57684 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_626
timestamp 1607194113
transform 1 0 58696 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_614
timestamp 1607194113
transform 1 0 57592 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A1_N
timestamp 1607194113
transform 1 0 58604 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 1607194113
transform 1 0 57776 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B1
timestamp 1607194113
transform 1 0 58788 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1607194113
transform 1 0 57960 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0724_
timestamp 1607194113
transform 1 0 58972 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_647
timestamp 1607194113
transform 1 0 60628 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_638
timestamp 1607194113
transform 1 0 59800 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A1
timestamp 1607194113
transform 1 0 59892 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A2_N
timestamp 1607194113
transform 1 0 60444 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1607194113
transform 1 0 60076 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0742_
timestamp 1607194113
transform 1 0 60168 0 -1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_69_672
timestamp 1607194113
transform 1 0 62928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_659
timestamp 1607194113
transform 1 0 61732 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_668
timestamp 1607194113
transform 1 0 62560 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_656
timestamp 1607194113
transform 1 0 61456 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1607194113
transform 1 0 62836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_684
timestamp 1607194113
transform 1 0 64032 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_692
timestamp 1607194113
transform 1 0 64768 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_680
timestamp 1607194113
transform 1 0 63664 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_696
timestamp 1607194113
transform 1 0 65136 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_467
timestamp 1607194113
transform 1 0 44068 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1_N
timestamp 1607194113
transform 1 0 44344 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0809_
timestamp 1607194113
transform 1 0 44528 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_506
timestamp 1607194113
transform 1 0 47656 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_494
timestamp 1607194113
transform 1 0 46552 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2_N
timestamp 1607194113
transform 1 0 46368 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B1
timestamp 1607194113
transform 1 0 46184 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1607194113
transform 1 0 46000 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_520
timestamp 1607194113
transform 1 0 48944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_518
timestamp 1607194113
transform 1 0 48760 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1607194113
transform 1 0 48852 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_544
timestamp 1607194113
transform 1 0 51152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_532
timestamp 1607194113
transform 1 0 50048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_569
timestamp 1607194113
transform 1 0 53452 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_556
timestamp 1607194113
transform 1 0 52256 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0856_
timestamp 1607194113
transform 1 0 52624 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_581
timestamp 1607194113
transform 1 0 54556 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_577
timestamp 1607194113
transform 1 0 54188 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1607194113
transform 1 0 54464 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_605
timestamp 1607194113
transform 1 0 56764 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_593
timestamp 1607194113
transform 1 0 55660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_628
timestamp 1607194113
transform 1 0 58880 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_617
timestamp 1607194113
transform 1 0 57868 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1607194113
transform 1 0 58420 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1607194113
transform 1 0 58604 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_645
timestamp 1607194113
transform 1 0 60444 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_640
timestamp 1607194113
transform 1 0 59984 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1607194113
transform 1 0 60076 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1607194113
transform 1 0 60168 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_669
timestamp 1607194113
transform 1 0 62652 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_657
timestamp 1607194113
transform 1 0 61548 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1607194113
transform 1 0 64860 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_681
timestamp 1607194113
transform 1 0 63756 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1607194113
transform 1 0 65412 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_482
timestamp 1607194113
transform 1 0 45448 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_470
timestamp 1607194113
transform 1 0 44344 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_489
timestamp 1607194113
transform 1 0 46092 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B1
timestamp 1607194113
transform 1 0 46828 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1_N
timestamp 1607194113
transform 1 0 47012 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1607194113
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0784_
timestamp 1607194113
transform 1 0 47196 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_521
timestamp 1607194113
transform 1 0 49036 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2_N
timestamp 1607194113
transform 1 0 48852 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B2
timestamp 1607194113
transform 1 0 48668 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_545
timestamp 1607194113
transform 1 0 51244 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_533
timestamp 1607194113
transform 1 0 50140 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1607194113
transform 1 0 51612 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_562
timestamp 1607194113
transform 1 0 52808 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_550
timestamp 1607194113
transform 1 0 51704 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0785_
timestamp 1607194113
transform 1 0 53084 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_586
timestamp 1607194113
transform 1 0 55016 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_574
timestamp 1607194113
transform 1 0 53912 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_611
timestamp 1607194113
transform 1 0 57316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_598
timestamp 1607194113
transform 1 0 56120 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1607194113
transform 1 0 57224 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_631
timestamp 1607194113
transform 1 0 59156 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_623
timestamp 1607194113
transform 1 0 58420 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_i_A
timestamp 1607194113
transform 1 0 58696 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_i
timestamp 1607194113
transform 1 0 58880 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1476_
timestamp 1607194113
transform 1 0 59248 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_653
timestamp 1607194113
transform 1 0 61180 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__CLK
timestamp 1607194113
transform 1 0 60996 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_672
timestamp 1607194113
transform 1 0 62928 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1607194113
transform 1 0 62284 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1607194113
transform 1 0 62836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_684
timestamp 1607194113
transform 1 0 64032 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_696
timestamp 1607194113
transform 1 0 65136 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1607194113
transform 1 0 65320 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_479
timestamp 1607194113
transform 1 0 45172 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_471
timestamp 1607194113
transform 1 0 44436 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1_N
timestamp 1607194113
transform 1 0 45448 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1607194113
transform 1 0 45632 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0780_
timestamp 1607194113
transform 1 0 45816 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_504
timestamp 1607194113
transform 1 0 47472 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2_N
timestamp 1607194113
transform 1 0 47288 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_520
timestamp 1607194113
transform 1 0 48944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_516
timestamp 1607194113
transform 1 0 48576 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1607194113
transform 1 0 48852 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_548
timestamp 1607194113
transform 1 0 51520 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_544
timestamp 1607194113
transform 1 0 51152 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_532
timestamp 1607194113
transform 1 0 50048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1
timestamp 1607194113
transform 1 0 51612 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2_N
timestamp 1607194113
transform 1 0 53452 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1_N
timestamp 1607194113
transform 1 0 51796 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0777_
timestamp 1607194113
transform 1 0 51980 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_581
timestamp 1607194113
transform 1 0 54556 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_579
timestamp 1607194113
transform 1 0 54372 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_571
timestamp 1607194113
transform 1 0 53636 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1607194113
transform 1 0 54464 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_605
timestamp 1607194113
transform 1 0 56764 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_593
timestamp 1607194113
transform 1 0 55660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_629
timestamp 1607194113
transform 1 0 58972 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_617
timestamp 1607194113
transform 1 0 57868 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_647
timestamp 1607194113
transform 1 0 60628 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1607194113
transform 1 0 60444 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1607194113
transform 1 0 60076 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1607194113
transform 1 0 60168 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_671
timestamp 1607194113
transform 1 0 62836 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_659
timestamp 1607194113
transform 1 0 61732 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_695
timestamp 1607194113
transform 1 0 65044 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_683
timestamp 1607194113
transform 1 0 63940 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_482
timestamp 1607194113
transform 1 0 45448 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_476
timestamp 1607194113
transform 1 0 44896 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1_N
timestamp 1607194113
transform 1 0 45724 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B1
timestamp 1607194113
transform 1 0 45540 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_507
timestamp 1607194113
transform 1 0 47748 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_487
timestamp 1607194113
transform 1 0 45908 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A2_N
timestamp 1607194113
transform 1 0 47564 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1607194113
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0852_
timestamp 1607194113
transform 1 0 46092 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_519
timestamp 1607194113
transform 1 0 48852 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_548
timestamp 1607194113
transform 1 0 51520 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_543
timestamp 1607194113
transform 1 0 51060 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_531
timestamp 1607194113
transform 1 0 49956 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B1
timestamp 1607194113
transform 1 0 51336 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A1_N
timestamp 1607194113
transform 1 0 51152 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1607194113
transform 1 0 51612 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_568
timestamp 1607194113
transform 1 0 53360 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A2_N
timestamp 1607194113
transform 1 0 53176 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0851_
timestamp 1607194113
transform 1 0 51704 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_580
timestamp 1607194113
transform 1 0 54464 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_611
timestamp 1607194113
transform 1 0 57316 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_604
timestamp 1607194113
transform 1 0 56672 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_592
timestamp 1607194113
transform 1 0 55568 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1607194113
transform 1 0 57224 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_619
timestamp 1607194113
transform 1 0 58052 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1607194113
transform 1 0 58144 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_73_641
timestamp 1607194113
transform 1 0 60076 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__CLK
timestamp 1607194113
transform 1 0 59892 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1077_
timestamp 1607194113
transform 1 0 60628 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_73_672
timestamp 1607194113
transform 1 0 62928 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_670
timestamp 1607194113
transform 1 0 62744 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_666
timestamp 1607194113
transform 1 0 62376 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_654
timestamp 1607194113
transform 1 0 61272 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1607194113
transform 1 0 62836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_684
timestamp 1607194113
transform 1 0 64032 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__CLK
timestamp 1607194113
transform 1 0 64216 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1472_
timestamp 1607194113
transform 1 0 64400 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_476
timestamp 1607194113
transform 1 0 44896 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_471
timestamp 1607194113
transform 1 0 44436 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A1_N
timestamp 1607194113
transform 1 0 44620 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1
timestamp 1607194113
transform 1 0 44804 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0832_
timestamp 1607194113
transform 1 0 44988 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_501
timestamp 1607194113
transform 1 0 47196 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_489
timestamp 1607194113
transform 1 0 46092 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_497
timestamp 1607194113
transform 1 0 46828 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B2
timestamp 1607194113
transform 1 0 46644 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A2_N
timestamp 1607194113
transform 1 0 46460 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1607194113
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_525
timestamp 1607194113
transform 1 0 49404 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_513
timestamp 1607194113
transform 1 0 48300 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_520
timestamp 1607194113
transform 1 0 48944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_517
timestamp 1607194113
transform 1 0 48668 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_509
timestamp 1607194113
transform 1 0 47932 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1607194113
transform 1 0 48852 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_537
timestamp 1607194113
transform 1 0 50508 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_532
timestamp 1607194113
transform 1 0 50048 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_548
timestamp 1607194113
transform 1 0 51520 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_543
timestamp 1607194113
transform 1 0 51060 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_540
timestamp 1607194113
transform 1 0 50784 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B1
timestamp 1607194113
transform 1 0 51336 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A1_N
timestamp 1607194113
transform 1 0 51152 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B1
timestamp 1607194113
transform 1 0 51060 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1_N
timestamp 1607194113
transform 1 0 51244 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1607194113
transform 1 0 51612 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0769_
timestamp 1607194113
transform 1 0 51428 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_570
timestamp 1607194113
transform 1 0 53544 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_567
timestamp 1607194113
transform 1 0 53268 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A2_N
timestamp 1607194113
transform 1 0 53084 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A2_N
timestamp 1607194113
transform 1 0 53360 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B2
timestamp 1607194113
transform 1 0 52900 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B2
timestamp 1607194113
transform 1 0 53176 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0845_
timestamp 1607194113
transform 1 0 51704 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_582
timestamp 1607194113
transform 1 0 54648 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_581
timestamp 1607194113
transform 1 0 54556 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_579
timestamp 1607194113
transform 1 0 54372 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1607194113
transform 1 0 54464 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_611
timestamp 1607194113
transform 1 0 57316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_606
timestamp 1607194113
transform 1 0 56856 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_594
timestamp 1607194113
transform 1 0 55752 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_605
timestamp 1607194113
transform 1 0 56764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_593
timestamp 1607194113
transform 1 0 55660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1607194113
transform 1 0 57224 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_630
timestamp 1607194113
transform 1 0 59064 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_623
timestamp 1607194113
transform 1 0 58420 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_623
timestamp 1607194113
transform 1 0 58420 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_617
timestamp 1607194113
transform 1 0 57868 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1078_
timestamp 1607194113
transform 1 0 58512 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1607194113
transform 1 0 58788 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_649
timestamp 1607194113
transform 1 0 60812 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_651
timestamp 1607194113
transform 1 0 60996 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_635
timestamp 1607194113
transform 1 0 59524 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1607194113
transform 1 0 60628 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1607194113
transform 1 0 59340 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1607194113
transform 1 0 60076 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1075_
timestamp 1607194113
transform 1 0 59800 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 60168 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_672
timestamp 1607194113
transform 1 0 62928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_670
timestamp 1607194113
transform 1 0 62744 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_662
timestamp 1607194113
transform 1 0 62008 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_663
timestamp 1607194113
transform 1 0 62100 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1607194113
transform 1 0 62836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1069_
timestamp 1607194113
transform 1 0 61364 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_75_684
timestamp 1607194113
transform 1 0 64032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_687
timestamp 1607194113
transform 1 0 64308 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_675
timestamp 1607194113
transform 1 0 63204 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_696
timestamp 1607194113
transform 1 0 65136 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_699
timestamp 1607194113
transform 1 0 65412 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_76_471
timestamp 1607194113
transform 1 0 44436 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1_N
timestamp 1607194113
transform 1 0 44712 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1607194113
transform 1 0 44896 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0753_
timestamp 1607194113
transform 1 0 45080 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_498
timestamp 1607194113
transform 1 0 46920 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B2
timestamp 1607194113
transform 1 0 46736 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2_N
timestamp 1607194113
transform 1 0 46552 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_520
timestamp 1607194113
transform 1 0 48944 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_518
timestamp 1607194113
transform 1 0 48760 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_510
timestamp 1607194113
transform 1 0 48024 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1607194113
transform 1 0 48852 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_540
timestamp 1607194113
transform 1 0 50784 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_532
timestamp 1607194113
transform 1 0 50048 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _0772_
timestamp 1607194113
transform 1 0 51060 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_561
timestamp 1607194113
transform 1 0 52716 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2_N
timestamp 1607194113
transform 1 0 52532 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_590
timestamp 1607194113
transform 1 0 55384 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_579
timestamp 1607194113
transform 1 0 54372 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_573
timestamp 1607194113
transform 1 0 53820 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1607194113
transform 1 0 54464 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0850_
timestamp 1607194113
transform 1 0 54556 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_76_602
timestamp 1607194113
transform 1 0 56488 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_626
timestamp 1607194113
transform 1 0 58696 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_614
timestamp 1607194113
transform 1 0 57592 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1607194113
transform 1 0 59156 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1607194113
transform 1 0 58880 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_649
timestamp 1607194113
transform 1 0 60812 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_633
timestamp 1607194113
transform 1 0 59340 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1607194113
transform 1 0 60076 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1068_
timestamp 1607194113
transform 1 0 60168 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_76_664
timestamp 1607194113
transform 1 0 62192 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1070_
timestamp 1607194113
transform 1 0 61548 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_76_688
timestamp 1607194113
transform 1 0 64400 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_676
timestamp 1607194113
transform 1 0 63296 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_477
timestamp 1607194113
transform 1 0 44988 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1607194113
transform 1 0 45724 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1_N
timestamp 1607194113
transform 1 0 45540 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_507
timestamp 1607194113
transform 1 0 47748 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_487
timestamp 1607194113
transform 1 0 45908 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B2
timestamp 1607194113
transform 1 0 47564 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1607194113
transform 1 0 46000 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0849_
timestamp 1607194113
transform 1 0 46092 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_519
timestamp 1607194113
transform 1 0 48852 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_543
timestamp 1607194113
transform 1 0 51060 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_531
timestamp 1607194113
transform 1 0 49956 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1607194113
transform 1 0 51612 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_568
timestamp 1607194113
transform 1 0 53360 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2_N
timestamp 1607194113
transform 1 0 53176 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0847_
timestamp 1607194113
transform 1 0 51704 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_580
timestamp 1607194113
transform 1 0 54464 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_611
timestamp 1607194113
transform 1 0 57316 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_604
timestamp 1607194113
transform 1 0 56672 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_592
timestamp 1607194113
transform 1 0 55568 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1607194113
transform 1 0 57224 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1079_
timestamp 1607194113
transform 1 0 58420 0 1 44064
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_77_639
timestamp 1607194113
transform 1 0 59892 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1607194113
transform 1 0 59708 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1050_
timestamp 1607194113
transform 1 0 60444 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_77_672
timestamp 1607194113
transform 1 0 62928 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_670
timestamp 1607194113
transform 1 0 62744 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_666
timestamp 1607194113
transform 1 0 62376 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_654
timestamp 1607194113
transform 1 0 61272 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1607194113
transform 1 0 62836 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_692
timestamp 1607194113
transform 1 0 64768 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_684
timestamp 1607194113
transform 1 0 64032 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0751_
timestamp 1607194113
transform 1 0 65044 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1607194113
transform 1 0 65412 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1607194113
transform 1 0 44436 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1_N
timestamp 1607194113
transform 1 0 44620 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0774_
timestamp 1607194113
transform 1 0 44804 0 -1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_78_505
timestamp 1607194113
transform 1 0 47564 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_493
timestamp 1607194113
transform 1 0 46460 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B2
timestamp 1607194113
transform 1 0 46276 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_520
timestamp 1607194113
transform 1 0 48944 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_517
timestamp 1607194113
transform 1 0 48668 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1607194113
transform 1 0 48852 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_544
timestamp 1607194113
transform 1 0 51152 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_532
timestamp 1607194113
transform 1 0 50048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_565
timestamp 1607194113
transform 1 0 53084 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0775_
timestamp 1607194113
transform 1 0 52256 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_78_581
timestamp 1607194113
transform 1 0 54556 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_577
timestamp 1607194113
transform 1 0 54188 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1607194113
transform 1 0 54464 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_611
timestamp 1607194113
transform 1 0 57316 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_605
timestamp 1607194113
transform 1 0 56764 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_593
timestamp 1607194113
transform 1 0 55660 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__CLK
timestamp 1607194113
transform 1 0 59156 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1474_
timestamp 1607194113
transform 1 0 57408 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_78_649
timestamp 1607194113
transform 1 0 60812 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_633
timestamp 1607194113
transform 1 0 59340 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1607194113
transform 1 0 60076 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1032_
timestamp 1607194113
transform 1 0 60168 0 -1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_78_660
timestamp 1607194113
transform 1 0 61824 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk_i
timestamp 1607194113
transform 1 0 61548 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1072_
timestamp 1607194113
transform 1 0 62376 0 -1 45152
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_78_693
timestamp 1607194113
transform 1 0 64860 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_681
timestamp 1607194113
transform 1 0 63756 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1607194113
transform 1 0 63572 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_486
timestamp 1607194113
transform 1 0 45816 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_474
timestamp 1607194113
transform 1 0 44712 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_470
timestamp 1607194113
transform 1 0 44344 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1607194113
transform 1 0 44436 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_504
timestamp 1607194113
transform 1 0 47472 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_492
timestamp 1607194113
transform 1 0 46368 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1607194113
transform 1 0 46000 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1607194113
transform 1 0 46092 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_528
timestamp 1607194113
transform 1 0 49680 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_516
timestamp 1607194113
transform 1 0 48576 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_544
timestamp 1607194113
transform 1 0 51152 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_540
timestamp 1607194113
transform 1 0 50784 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A1_N
timestamp 1607194113
transform 1 0 51244 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B1
timestamp 1607194113
transform 1 0 51428 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1607194113
transform 1 0 51612 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_566
timestamp 1607194113
transform 1 0 53176 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0843_
timestamp 1607194113
transform 1 0 51704 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_79_590
timestamp 1607194113
transform 1 0 55384 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_578
timestamp 1607194113
transform 1 0 54280 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_611
timestamp 1607194113
transform 1 0 57316 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_602
timestamp 1607194113
transform 1 0 56488 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_596
timestamp 1607194113
transform 1 0 55936 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1607194113
transform 1 0 56304 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1607194113
transform 1 0 57224 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1607194113
transform 1 0 56028 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_622
timestamp 1607194113
transform 1 0 58328 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1607194113
transform 1 0 58052 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_646
timestamp 1607194113
transform 1 0 60536 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_634
timestamp 1607194113
transform 1 0 59432 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_672
timestamp 1607194113
transform 1 0 62928 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_670
timestamp 1607194113
transform 1 0 62744 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_658
timestamp 1607194113
transform 1 0 61640 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1607194113
transform 1 0 62836 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_684
timestamp 1607194113
transform 1 0 64032 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_696
timestamp 1607194113
transform 1 0 65136 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_715
timestamp 1607194113
transform 1 0 66884 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_703
timestamp 1607194113
transform 1 0 65780 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607194113
transform 1 0 65688 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1373_
timestamp 1607194113
transform 1 0 67620 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_756
timestamp 1607194113
transform 1 0 70656 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_744
timestamp 1607194113
transform 1 0 69552 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1607194113
transform 1 0 69368 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_762
timestamp 1607194113
transform 1 0 71208 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A2_N
timestamp 1607194113
transform 1 0 71024 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B2
timestamp 1607194113
transform 1 0 71392 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607194113
transform 1 0 71300 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1212_
timestamp 1607194113
transform 1 0 71576 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_50_784
timestamp 1607194113
transform 1 0 73232 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A1_N
timestamp 1607194113
transform 1 0 73048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1414_
timestamp 1607194113
transform 1 0 73784 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_811
timestamp 1607194113
transform 1 0 75716 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__CLK
timestamp 1607194113
transform 1 0 75532 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_837
timestamp 1607194113
transform 1 0 78108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_825
timestamp 1607194113
transform 1 0 77004 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_823
timestamp 1607194113
transform 1 0 76820 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607194113
transform 1 0 76912 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_852
timestamp 1607194113
transform 1 0 79488 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1607194113
transform 1 0 79212 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_866
timestamp 1607194113
transform 1 0 80776 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_860
timestamp 1607194113
transform 1 0 80224 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1607194113
transform 1 0 80500 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_886
timestamp 1607194113
transform 1 0 82616 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_884
timestamp 1607194113
transform 1 0 82432 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_878
timestamp 1607194113
transform 1 0 81880 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607194113
transform 1 0 82524 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_910
timestamp 1607194113
transform 1 0 84824 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_898
timestamp 1607194113
transform 1 0 83720 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_922
timestamp 1607194113
transform 1 0 85928 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[4]
timestamp 1607194113
transform 1 0 86664 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[2]
timestamp 1607194113
transform 1 0 86296 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[0]
timestamp 1607194113
transform 1 0 86480 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_inp_i
timestamp 1607194113
transform 1 0 86848 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A2_N
timestamp 1607194113
transform 1 0 65688 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B2
timestamp 1607194113
transform 1 0 65872 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B1
timestamp 1607194113
transform 1 0 66056 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1274_
timestamp 1607194113
transform 1 0 66240 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_738
timestamp 1607194113
transform 1 0 69000 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_724
timestamp 1607194113
transform 1 0 67712 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1607194113
transform 1 0 68816 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607194113
transform 1 0 68448 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1607194113
transform 1 0 68540 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_750
timestamp 1607194113
transform 1 0 70104 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_778
timestamp 1607194113
transform 1 0 72680 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_766
timestamp 1607194113
transform 1 0 71576 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_762
timestamp 1607194113
transform 1 0 71208 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B1
timestamp 1607194113
transform 1 0 71392 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_794
timestamp 1607194113
transform 1 0 74152 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_790
timestamp 1607194113
transform 1 0 73784 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607194113
transform 1 0 74060 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1607194113
transform 1 0 74336 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_811
timestamp 1607194113
transform 1 0 75716 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_799
timestamp 1607194113
transform 1 0 74612 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_835
timestamp 1607194113
transform 1 0 77924 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_823
timestamp 1607194113
transform 1 0 76820 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_851
timestamp 1607194113
transform 1 0 79396 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_847
timestamp 1607194113
transform 1 0 79028 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__CLK
timestamp 1607194113
transform 1 0 79488 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607194113
transform 1 0 79672 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1607194113
transform 1 0 79764 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_874
timestamp 1607194113
transform 1 0 81512 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_886
timestamp 1607194113
transform 1 0 82616 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_916
timestamp 1607194113
transform 1 0 85376 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_909
timestamp 1607194113
transform 1 0 84732 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_898
timestamp 1607194113
transform 1 0 83720 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1607194113
transform 1 0 84548 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607194113
transform 1 0 85284 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1607194113
transform 1 0 84272 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_931
timestamp 1607194113
transform 1 0 86756 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[1]
timestamp 1607194113
transform 1 0 86848 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1141_
timestamp 1607194113
transform 1 0 86112 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_52_703
timestamp 1607194113
transform 1 0 65780 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1_N
timestamp 1607194113
transform 1 0 66056 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607194113
transform 1 0 65688 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0825_
timestamp 1607194113
transform 1 0 66240 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B2
timestamp 1607194113
transform 1 0 67896 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1607194113
transform 1 0 68080 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1_N
timestamp 1607194113
transform 1 0 68264 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A2_N
timestamp 1607194113
transform 1 0 67712 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0838_
timestamp 1607194113
transform 1 0 68448 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_752
timestamp 1607194113
transform 1 0 70288 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A2_N
timestamp 1607194113
transform 1 0 70104 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B2
timestamp 1607194113
transform 1 0 69920 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_776
timestamp 1607194113
transform 1 0 72496 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_764
timestamp 1607194113
transform 1 0 71392 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_760
timestamp 1607194113
transform 1 0 71024 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607194113
transform 1 0 71300 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_782
timestamp 1607194113
transform 1 0 73048 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A1_N
timestamp 1607194113
transform 1 0 73140 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B1
timestamp 1607194113
transform 1 0 73324 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0727_
timestamp 1607194113
transform 1 0 73508 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_807
timestamp 1607194113
transform 1 0 75348 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A2_N
timestamp 1607194113
transform 1 0 75164 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B2
timestamp 1607194113
transform 1 0 74980 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_837
timestamp 1607194113
transform 1 0 78108 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_825
timestamp 1607194113
transform 1 0 77004 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_823
timestamp 1607194113
transform 1 0 76820 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_819
timestamp 1607194113
transform 1 0 76452 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607194113
transform 1 0 76912 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 1607194113
transform 1 0 78660 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1147_
timestamp 1607194113
transform 1 0 78844 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_52_871
timestamp 1607194113
transform 1 0 81236 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_861
timestamp 1607194113
transform 1 0 80316 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A1
timestamp 1607194113
transform 1 0 80132 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1607194113
transform 1 0 80684 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0738_
timestamp 1607194113
transform 1 0 80868 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_886
timestamp 1607194113
transform 1 0 82616 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_883
timestamp 1607194113
transform 1 0 82340 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607194113
transform 1 0 82524 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__CLK
timestamp 1607194113
transform 1 0 83720 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1607194113
transform 1 0 83904 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_52_919
timestamp 1607194113
transform 1 0 85652 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1607194113
transform 1 0 86204 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1043_
timestamp 1607194113
transform 1 0 86388 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_53_717
timestamp 1607194113
transform 1 0 67068 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_705
timestamp 1607194113
transform 1 0 65964 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_729
timestamp 1607194113
transform 1 0 68172 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607194113
transform 1 0 68448 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0826_
timestamp 1607194113
transform 1 0 68540 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_53_754
timestamp 1607194113
transform 1 0 70472 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_742
timestamp 1607194113
transform 1 0 69368 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_778
timestamp 1607194113
transform 1 0 72680 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_766
timestamp 1607194113
transform 1 0 71576 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_786
timestamp 1607194113
transform 1 0 73416 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1_N
timestamp 1607194113
transform 1 0 73692 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1
timestamp 1607194113
transform 1 0 73876 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607194113
transform 1 0 74060 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0818_
timestamp 1607194113
transform 1 0 74152 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_814
timestamp 1607194113
transform 1 0 75992 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2_N
timestamp 1607194113
transform 1 0 75808 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1607194113
transform 1 0 75624 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_826
timestamp 1607194113
transform 1 0 77096 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_850
timestamp 1607194113
transform 1 0 79304 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_838
timestamp 1607194113
transform 1 0 78200 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607194113
transform 1 0 79672 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1137_
timestamp 1607194113
transform 1 0 79764 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_876
timestamp 1607194113
transform 1 0 81696 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_864
timestamp 1607194113
transform 1 0 80592 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1607194113
transform 1 0 80408 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_888
timestamp 1607194113
transform 1 0 82800 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_880
timestamp 1607194113
transform 1 0 82064 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1607194113
transform 1 0 83536 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1138_
timestamp 1607194113
transform 1 0 82156 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_53_907
timestamp 1607194113
transform 1 0 84548 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1607194113
transform 1 0 85100 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607194113
transform 1 0 85284 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1143_
timestamp 1607194113
transform 1 0 83720 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1142_
timestamp 1607194113
transform 1 0 85376 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_53_925
timestamp 1607194113
transform 1 0 86204 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_703
timestamp 1607194113
transform 1 0 65780 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1_N
timestamp 1607194113
transform 1 0 66884 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B1
timestamp 1607194113
transform 1 0 67068 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607194113
transform 1 0 65688 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B2
timestamp 1607194113
transform 1 0 68908 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A2_N
timestamp 1607194113
transform 1 0 68724 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0823_
timestamp 1607194113
transform 1 0 67252 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_54_751
timestamp 1607194113
transform 1 0 70196 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_739
timestamp 1607194113
transform 1 0 69092 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_776
timestamp 1607194113
transform 1 0 72496 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_764
timestamp 1607194113
transform 1 0 71392 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607194113
transform 1 0 71300 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_788
timestamp 1607194113
transform 1 0 73600 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1607194113
transform 1 0 74336 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_818
timestamp 1607194113
transform 1 0 76360 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_54_809
timestamp 1607194113
transform 1 0 75532 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_801
timestamp 1607194113
transform 1 0 74796 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1607194113
transform 1 0 74612 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1607194113
transform 1 0 76176 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0726_
timestamp 1607194113
transform 1 0 75808 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_837
timestamp 1607194113
transform 1 0 78108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_825
timestamp 1607194113
transform 1 0 77004 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607194113
transform 1 0 76912 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_849
timestamp 1607194113
transform 1 0 79212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_874
timestamp 1607194113
transform 1 0 81512 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_861
timestamp 1607194113
transform 1 0 80316 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1607194113
transform 1 0 81328 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1047_
timestamp 1607194113
transform 1 0 80500 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_886
timestamp 1607194113
transform 1 0 82616 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_882
timestamp 1607194113
transform 1 0 82248 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607194113
transform 1 0 82524 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_910
timestamp 1607194113
transform 1 0 84824 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_898
timestamp 1607194113
transform 1 0 83720 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1607194113
transform 1 0 85376 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_919
timestamp 1607194113
transform 1 0 85652 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1145_
timestamp 1607194113
transform 1 0 86756 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_56_715
timestamp 1607194113
transform 1 0 66884 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_703
timestamp 1607194113
transform 1 0 65780 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_708
timestamp 1607194113
transform 1 0 66240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1_N
timestamp 1607194113
transform 1 0 66976 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607194113
transform 1 0 65688 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0821_
timestamp 1607194113
transform 1 0 67160 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_738
timestamp 1607194113
transform 1 0 69000 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_728
timestamp 1607194113
transform 1 0 68080 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_720
timestamp 1607194113
transform 1 0 67344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B1
timestamp 1607194113
transform 1 0 68264 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1607194113
transform 1 0 68816 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2_N
timestamp 1607194113
transform 1 0 68632 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607194113
transform 1 0 68448 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0837_
timestamp 1607194113
transform 1 0 68540 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_750
timestamp 1607194113
transform 1 0 70104 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_751
timestamp 1607194113
transform 1 0 70196 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A2_N
timestamp 1607194113
transform 1 0 70012 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_776
timestamp 1607194113
transform 1 0 72496 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_764
timestamp 1607194113
transform 1 0 71392 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_762
timestamp 1607194113
transform 1 0 71208 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_775
timestamp 1607194113
transform 1 0 72404 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_763
timestamp 1607194113
transform 1 0 71300 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607194113
transform 1 0 71300 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_798
timestamp 1607194113
transform 1 0 74520 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_784
timestamp 1607194113
transform 1 0 73232 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_787
timestamp 1607194113
transform 1 0 73508 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607194113
transform 1 0 74060 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1607194113
transform 1 0 74152 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1152_
timestamp 1607194113
transform 1 0 73416 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_813
timestamp 1607194113
transform 1 0 75900 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_806
timestamp 1607194113
transform 1 0 75256 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_815
timestamp 1607194113
transform 1 0 76084 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__CLK
timestamp 1607194113
transform 1 0 75900 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1607194113
transform 1 0 75716 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1607194113
transform 1 0 75440 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_836
timestamp 1607194113
transform 1 0 78016 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_825
timestamp 1607194113
transform 1 0 77004 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_821
timestamp 1607194113
transform 1 0 76636 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_827
timestamp 1607194113
transform 1 0 77188 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk_i
timestamp 1607194113
transform 1 0 77740 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607194113
transform 1 0 76912 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_848
timestamp 1607194113
transform 1 0 79120 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_855
timestamp 1607194113
transform 1 0 79764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_851
timestamp 1607194113
transform 1 0 79396 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_839
timestamp 1607194113
transform 1 0 78292 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607194113
transform 1 0 79672 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_877
timestamp 1607194113
transform 1 0 81788 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_865
timestamp 1607194113
transform 1 0 80684 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_860
timestamp 1607194113
transform 1 0 80224 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_873
timestamp 1607194113
transform 1 0 81420 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_867
timestamp 1607194113
transform 1 0 80868 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1140_
timestamp 1607194113
transform 1 0 81512 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0734_
timestamp 1607194113
transform 1 0 81420 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1607194113
transform 1 0 80408 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_888
timestamp 1607194113
transform 1 0 82800 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B1
timestamp 1607194113
transform 1 0 82156 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1607194113
transform 1 0 82340 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1607194113
transform 1 0 82616 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607194113
transform 1 0 82524 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1139_
timestamp 1607194113
transform 1 0 82616 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_56_911
timestamp 1607194113
transform 1 0 84916 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_899
timestamp 1607194113
transform 1 0 83812 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_916
timestamp 1607194113
transform 1 0 85376 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_912
timestamp 1607194113
transform 1 0 85008 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_900
timestamp 1607194113
transform 1 0 83904 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 1607194113
transform 1 0 85284 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A1
timestamp 1607194113
transform 1 0 85468 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607194113
transform 1 0 85284 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_928
timestamp 1607194113
transform 1 0 86480 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _1135_
timestamp 1607194113
transform 1 0 85652 0 -1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_57_708
timestamp 1607194113
transform 1 0 66240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_720
timestamp 1607194113
transform 1 0 67344 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607194113
transform 1 0 68448 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0841_
timestamp 1607194113
transform 1 0 68540 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_754
timestamp 1607194113
transform 1 0 70472 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_742
timestamp 1607194113
transform 1 0 69368 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_778
timestamp 1607194113
transform 1 0 72680 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_766
timestamp 1607194113
transform 1 0 71576 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_794
timestamp 1607194113
transform 1 0 74152 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_790
timestamp 1607194113
transform 1 0 73784 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607194113
transform 1 0 74060 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_806
timestamp 1607194113
transform 1 0 75256 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1607194113
transform 1 0 75992 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_835
timestamp 1607194113
transform 1 0 77924 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1607194113
transform 1 0 77740 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_855
timestamp 1607194113
transform 1 0 79764 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_853
timestamp 1607194113
transform 1 0 79580 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_847
timestamp 1607194113
transform 1 0 79028 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607194113
transform 1 0 79672 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_863
timestamp 1607194113
transform 1 0 80500 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__CLK
timestamp 1607194113
transform 1 0 80684 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1457_
timestamp 1607194113
transform 1 0 80868 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_886
timestamp 1607194113
transform 1 0 82616 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_914
timestamp 1607194113
transform 1 0 85192 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_910
timestamp 1607194113
transform 1 0 84824 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_898
timestamp 1607194113
transform 1 0 83720 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607194113
transform 1 0 85284 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1607194113
transform 1 0 85376 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_927
timestamp 1607194113
transform 1 0 86388 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_919
timestamp 1607194113
transform 1 0 85652 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1607194113
transform 1 0 86572 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1130_
timestamp 1607194113
transform 1 0 86756 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_58_715
timestamp 1607194113
transform 1 0 66884 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_703
timestamp 1607194113
transform 1 0 65780 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_700
timestamp 1607194113
transform 1 0 65504 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607194113
transform 1 0 65688 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1420_
timestamp 1607194113
transform 1 0 67160 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__CLK
timestamp 1607194113
transform 1 0 68908 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_751
timestamp 1607194113
transform 1 0 70196 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_739
timestamp 1607194113
transform 1 0 69092 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_776
timestamp 1607194113
transform 1 0 72496 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_764
timestamp 1607194113
transform 1 0 71392 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607194113
transform 1 0 71300 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B1
timestamp 1607194113
transform 1 0 74428 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1151_
timestamp 1607194113
transform 1 0 73232 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_58_818
timestamp 1607194113
transform 1 0 76360 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_799
timestamp 1607194113
transform 1 0 74612 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1607194113
transform 1 0 76176 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1607194113
transform 1 0 75164 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1046_
timestamp 1607194113
transform 1 0 75348 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_834
timestamp 1607194113
transform 1 0 77832 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607194113
transform 1 0 76912 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1154_
timestamp 1607194113
transform 1 0 77004 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_846
timestamp 1607194113
transform 1 0 78936 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_870
timestamp 1607194113
transform 1 0 81144 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_858
timestamp 1607194113
transform 1 0 80040 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_886
timestamp 1607194113
transform 1 0 82616 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_882
timestamp 1607194113
transform 1 0 82248 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__CLK
timestamp 1607194113
transform 1 0 83168 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607194113
transform 1 0 82524 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1607194113
transform 1 0 83352 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_58_913
timestamp 1607194113
transform 1 0 85100 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_925
timestamp 1607194113
transform 1 0 86204 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_716
timestamp 1607194113
transform 1 0 66976 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_704
timestamp 1607194113
transform 1 0 65872 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_700
timestamp 1607194113
transform 1 0 65504 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1607194113
transform 1 0 65596 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_729
timestamp 1607194113
transform 1 0 68172 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_724
timestamp 1607194113
transform 1 0 67712 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A1_N
timestamp 1607194113
transform 1 0 67988 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B1
timestamp 1607194113
transform 1 0 67804 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A2_N
timestamp 1607194113
transform 1 0 68264 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607194113
transform 1 0 68448 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0836_
timestamp 1607194113
transform 1 0 68540 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_751
timestamp 1607194113
transform 1 0 70196 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B2
timestamp 1607194113
transform 1 0 70012 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_775
timestamp 1607194113
transform 1 0 72404 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_763
timestamp 1607194113
transform 1 0 71300 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_794
timestamp 1607194113
transform 1 0 74152 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_787
timestamp 1607194113
transform 1 0 73508 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607194113
transform 1 0 74060 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_817
timestamp 1607194113
transform 1 0 76268 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1607194113
transform 1 0 76084 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1153_
timestamp 1607194113
transform 1 0 75256 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_59_830
timestamp 1607194113
transform 1 0 77464 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A
timestamp 1607194113
transform 1 0 76636 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1149_
timestamp 1607194113
transform 1 0 76820 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_59_855
timestamp 1607194113
transform 1 0 79764 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_842
timestamp 1607194113
transform 1 0 78568 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607194113
transform 1 0 79672 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_867
timestamp 1607194113
transform 1 0 80868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_891
timestamp 1607194113
transform 1 0 83076 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_879
timestamp 1607194113
transform 1 0 81972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_903
timestamp 1607194113
transform 1 0 84180 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607194113
transform 1 0 85284 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1607194113
transform 1 0 85376 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_931
timestamp 1607194113
transform 1 0 86756 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_919
timestamp 1607194113
transform 1 0 85652 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_715
timestamp 1607194113
transform 1 0 66884 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_703
timestamp 1607194113
transform 1 0 65780 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1607194113
transform 1 0 65688 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_729
timestamp 1607194113
transform 1 0 68172 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_723
timestamp 1607194113
transform 1 0 67620 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1607194113
transform 1 0 67896 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_753
timestamp 1607194113
transform 1 0 70380 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_741
timestamp 1607194113
transform 1 0 69276 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_776
timestamp 1607194113
transform 1 0 72496 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_770
timestamp 1607194113
transform 1 0 71944 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_764
timestamp 1607194113
transform 1 0 71392 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_761
timestamp 1607194113
transform 1 0 71116 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1607194113
transform 1 0 72312 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1607194113
transform 1 0 71300 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1607194113
transform 1 0 72036 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_788
timestamp 1607194113
transform 1 0 73600 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_812
timestamp 1607194113
transform 1 0 75808 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_800
timestamp 1607194113
transform 1 0 74704 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1607194113
transform 1 0 75624 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1150_
timestamp 1607194113
transform 1 0 74980 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_60_828
timestamp 1607194113
transform 1 0 77280 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1607194113
transform 1 0 76912 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1607194113
transform 1 0 77004 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_854
timestamp 1607194113
transform 1 0 79672 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_848
timestamp 1607194113
transform 1 0 79120 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_840
timestamp 1607194113
transform 1 0 78384 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1117_
timestamp 1607194113
transform 1 0 79304 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_866
timestamp 1607194113
transform 1 0 80776 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_886
timestamp 1607194113
transform 1 0 82616 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_884
timestamp 1607194113
transform 1 0 82432 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_878
timestamp 1607194113
transform 1 0 81880 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1607194113
transform 1 0 82524 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_910
timestamp 1607194113
transform 1 0 84824 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_898
timestamp 1607194113
transform 1 0 83720 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_922
timestamp 1607194113
transform 1 0 85928 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_715
timestamp 1607194113
transform 1 0 66884 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_703
timestamp 1607194113
transform 1 0 65780 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_701
timestamp 1607194113
transform 1 0 65596 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B1
timestamp 1607194113
transform 1 0 65596 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B2
timestamp 1607194113
transform 1 0 67068 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1607194113
transform 1 0 65688 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0794_
timestamp 1607194113
transform 1 0 65780 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _0694_
timestamp 1607194113
transform 1 0 66976 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_736
timestamp 1607194113
transform 1 0 68816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_733
timestamp 1607194113
transform 1 0 68540 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_729
timestamp 1607194113
transform 1 0 68172 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_721
timestamp 1607194113
transform 1 0 67436 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A2
timestamp 1607194113
transform 1 0 68632 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A2
timestamp 1607194113
transform 1 0 67252 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B2
timestamp 1607194113
transform 1 0 68448 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B1
timestamp 1607194113
transform 1 0 68264 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1607194113
transform 1 0 68448 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_748
timestamp 1607194113
transform 1 0 69920 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_757
timestamp 1607194113
transform 1 0 70748 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_745
timestamp 1607194113
transform 1 0 69644 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_764
timestamp 1607194113
transform 1 0 71392 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_760
timestamp 1607194113
transform 1 0 71024 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_775
timestamp 1607194113
transform 1 0 72404 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_763
timestamp 1607194113
transform 1 0 71300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A
timestamp 1607194113
transform 1 0 72220 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B
timestamp 1607194113
transform 1 0 72036 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1607194113
transform 1 0 71300 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1450_
timestamp 1607194113
transform 1 0 71484 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1157_
timestamp 1607194113
transform 1 0 71392 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_62_794
timestamp 1607194113
transform 1 0 74152 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_786
timestamp 1607194113
transform 1 0 73416 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_787
timestamp 1607194113
transform 1 0 73508 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1607194113
transform 1 0 73232 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_i_A
timestamp 1607194113
transform 1 0 74428 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1607194113
transform 1 0 74060 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1155_
timestamp 1607194113
transform 1 0 74152 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_62_813
timestamp 1607194113
transform 1 0 75900 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_802
timestamp 1607194113
transform 1 0 74888 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_805
timestamp 1607194113
transform 1 0 75164 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1607194113
transform 1 0 74796 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1607194113
transform 1 0 74980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_i
timestamp 1607194113
transform 1 0 74612 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1451_
timestamp 1607194113
transform 1 0 75532 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1156_
timestamp 1607194113
transform 1 0 75072 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_837
timestamp 1607194113
transform 1 0 78108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_825
timestamp 1607194113
transform 1 0 77004 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_821
timestamp 1607194113
transform 1 0 76636 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_830
timestamp 1607194113
transform 1 0 77464 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1607194113
transform 1 0 77280 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1607194113
transform 1 0 76912 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_849
timestamp 1607194113
transform 1 0 79212 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_850
timestamp 1607194113
transform 1 0 79304 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_842
timestamp 1607194113
transform 1 0 78568 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__CLK
timestamp 1607194113
transform 1 0 79488 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1607194113
transform 1 0 79580 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1607194113
transform 1 0 79672 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1463_
timestamp 1607194113
transform 1 0 79764 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1120_
timestamp 1607194113
transform 1 0 79764 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_62_876
timestamp 1607194113
transform 1 0 81696 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_864
timestamp 1607194113
transform 1 0 80592 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_874
timestamp 1607194113
transform 1 0 81512 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_886
timestamp 1607194113
transform 1 0 82616 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_884
timestamp 1607194113
transform 1 0 82432 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_886
timestamp 1607194113
transform 1 0 82616 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1607194113
transform 1 0 82524 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_910
timestamp 1607194113
transform 1 0 84824 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_898
timestamp 1607194113
transform 1 0 83720 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_914
timestamp 1607194113
transform 1 0 85192 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_910
timestamp 1607194113
transform 1 0 84824 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_898
timestamp 1607194113
transform 1 0 83720 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1607194113
transform 1 0 85284 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1108_
timestamp 1607194113
transform 1 0 85376 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_62_925
timestamp 1607194113
transform 1 0 86204 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_918
timestamp 1607194113
transform 1 0 85560 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_927
timestamp 1607194113
transform 1 0 86388 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1607194113
transform 1 0 86020 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1607194113
transform 1 0 86572 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1607194113
transform 1 0 86204 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1123_
timestamp 1607194113
transform 1 0 86756 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1607194113
transform 1 0 85744 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_714
timestamp 1607194113
transform 1 0 66792 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_701
timestamp 1607194113
transform 1 0 65596 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _0795_
timestamp 1607194113
transform 1 0 65964 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_733
timestamp 1607194113
transform 1 0 68540 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_726
timestamp 1607194113
transform 1 0 67896 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1607194113
transform 1 0 68448 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_757
timestamp 1607194113
transform 1 0 70748 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_745
timestamp 1607194113
transform 1 0 69644 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1516_
timestamp 1607194113
transform 1 0 70840 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__CLK
timestamp 1607194113
transform 1 0 72588 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_794
timestamp 1607194113
transform 1 0 74152 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_791
timestamp 1607194113
transform 1 0 73876 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_779
timestamp 1607194113
transform 1 0 72772 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1607194113
transform 1 0 74060 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_817
timestamp 1607194113
transform 1 0 76268 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_812
timestamp 1607194113
transform 1 0 75808 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_806
timestamp 1607194113
transform 1 0 75256 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0700_
timestamp 1607194113
transform 1 0 75900 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_829
timestamp 1607194113
transform 1 0 77372 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_848
timestamp 1607194113
transform 1 0 79120 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_841
timestamp 1607194113
transform 1 0 78476 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1607194113
transform 1 0 78936 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1607194113
transform 1 0 79672 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1114_
timestamp 1607194113
transform 1 0 79764 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1607194113
transform 1 0 78660 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_872
timestamp 1607194113
transform 1 0 81328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_864
timestamp 1607194113
transform 1 0 80592 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1607194113
transform 1 0 80408 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1048_
timestamp 1607194113
transform 1 0 81420 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_63_894
timestamp 1607194113
transform 1 0 83352 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_882
timestamp 1607194113
transform 1 0 82248 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_916
timestamp 1607194113
transform 1 0 85376 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_913
timestamp 1607194113
transform 1 0 85100 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1607194113
transform 1 0 84916 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__C
timestamp 1607194113
transform 1 0 84732 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__D
timestamp 1607194113
transform 1 0 84548 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1607194113
transform 1 0 85284 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1040_
timestamp 1607194113
transform 1 0 83720 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B1
timestamp 1607194113
transform 1 0 85744 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A1
timestamp 1607194113
transform 1 0 85928 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1128_
timestamp 1607194113
transform 1 0 86112 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_64_712
timestamp 1607194113
transform 1 0 66608 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1607194113
transform 1 0 65688 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0695_
timestamp 1607194113
transform 1 0 65780 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_736
timestamp 1607194113
transform 1 0 68816 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_724
timestamp 1607194113
transform 1 0 67712 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_753
timestamp 1607194113
transform 1 0 70380 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_748
timestamp 1607194113
transform 1 0 69920 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1607194113
transform 1 0 70104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_777
timestamp 1607194113
transform 1 0 72588 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_772
timestamp 1607194113
transform 1 0 72128 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_764
timestamp 1607194113
transform 1 0 71392 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_761
timestamp 1607194113
transform 1 0 71116 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1607194113
transform 1 0 71300 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1607194113
transform 1 0 72220 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_789
timestamp 1607194113
transform 1 0 73692 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1607194113
transform 1 0 73324 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_813
timestamp 1607194113
transform 1 0 75900 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_801
timestamp 1607194113
transform 1 0 74796 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_837
timestamp 1607194113
transform 1 0 78108 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_825
timestamp 1607194113
transform 1 0 77004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_821
timestamp 1607194113
transform 1 0 76636 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1607194113
transform 1 0 76912 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_845
timestamp 1607194113
transform 1 0 78844 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 1607194113
transform 1 0 78936 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1607194113
transform 1 0 79120 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1041_
timestamp 1607194113
transform 1 0 79304 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_64_876
timestamp 1607194113
transform 1 0 81696 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_861
timestamp 1607194113
transform 1 0 80316 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1607194113
transform 1 0 81512 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__D
timestamp 1607194113
transform 1 0 80132 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1119_
timestamp 1607194113
transform 1 0 80868 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_64_886
timestamp 1607194113
transform 1 0 82616 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_884
timestamp 1607194113
transform 1 0 82432 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1607194113
transform 1 0 82524 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_916
timestamp 1607194113
transform 1 0 85376 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_910
timestamp 1607194113
transform 1 0 84824 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_898
timestamp 1607194113
transform 1 0 83720 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1607194113
transform 1 0 85468 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_930
timestamp 1607194113
transform 1 0 86664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B
timestamp 1607194113
transform 1 0 86480 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1109_
timestamp 1607194113
transform 1 0 85652 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_715
timestamp 1607194113
transform 1 0 66884 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_703
timestamp 1607194113
transform 1 0 65780 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_733
timestamp 1607194113
transform 1 0 68540 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_731
timestamp 1607194113
transform 1 0 68356 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_727
timestamp 1607194113
transform 1 0 67988 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1607194113
transform 1 0 68448 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_757
timestamp 1607194113
transform 1 0 70748 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_745
timestamp 1607194113
transform 1 0 69644 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_778
timestamp 1607194113
transform 1 0 72680 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_769
timestamp 1607194113
transform 1 0 71852 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1607194113
transform 1 0 72128 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1607194113
transform 1 0 72312 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_798
timestamp 1607194113
transform 1 0 74520 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_790
timestamp 1607194113
transform 1 0 73784 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1607194113
transform 1 0 74060 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1607194113
transform 1 0 74152 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_810
timestamp 1607194113
transform 1 0 75624 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_834
timestamp 1607194113
transform 1 0 77832 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_828
timestamp 1607194113
transform 1 0 77280 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_822
timestamp 1607194113
transform 1 0 76728 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1607194113
transform 1 0 77648 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1607194113
transform 1 0 77372 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_846
timestamp 1607194113
transform 1 0 78936 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1607194113
transform 1 0 79672 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1113_
timestamp 1607194113
transform 1 0 79764 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_65_874
timestamp 1607194113
transform 1 0 81512 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_864
timestamp 1607194113
transform 1 0 80592 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1607194113
transform 1 0 80408 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0744_
timestamp 1607194113
transform 1 0 81144 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_886
timestamp 1607194113
transform 1 0 82616 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_916
timestamp 1607194113
transform 1 0 85376 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_914
timestamp 1607194113
transform 1 0 85192 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_910
timestamp 1607194113
transform 1 0 84824 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_898
timestamp 1607194113
transform 1 0 83720 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1607194113
transform 1 0 85284 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_932
timestamp 1607194113
transform 1 0 86848 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_928
timestamp 1607194113
transform 1 0 86480 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1607194113
transform 1 0 86572 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_715
timestamp 1607194113
transform 1 0 66884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_703
timestamp 1607194113
transform 1 0 65780 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1607194113
transform 1 0 65688 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_727
timestamp 1607194113
transform 1 0 67988 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_751
timestamp 1607194113
transform 1 0 70196 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_739
timestamp 1607194113
transform 1 0 69092 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_777
timestamp 1607194113
transform 1 0 72588 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_772
timestamp 1607194113
transform 1 0 72128 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_764
timestamp 1607194113
transform 1 0 71392 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1607194113
transform 1 0 71300 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1607194113
transform 1 0 72220 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_789
timestamp 1607194113
transform 1 0 73692 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1607194113
transform 1 0 73324 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_813
timestamp 1607194113
transform 1 0 75900 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_801
timestamp 1607194113
transform 1 0 74796 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_825
timestamp 1607194113
transform 1 0 77004 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk_i
timestamp 1607194113
transform 1 0 76636 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1607194113
transform 1 0 76912 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1115_
timestamp 1607194113
transform 1 0 77372 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_66_857
timestamp 1607194113
transform 1 0 79948 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_840
timestamp 1607194113
transform 1 0 78384 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1607194113
transform 1 0 78568 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1607194113
transform 1 0 78200 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__C
timestamp 1607194113
transform 1 0 79764 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1607194113
transform 1 0 78752 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1110_
timestamp 1607194113
transform 1 0 78936 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_866
timestamp 1607194113
transform 1 0 80776 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1607194113
transform 1 0 80500 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_886
timestamp 1607194113
transform 1 0 82616 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_884
timestamp 1607194113
transform 1 0 82432 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_878
timestamp 1607194113
transform 1 0 81880 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B1
timestamp 1607194113
transform 1 0 82892 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1607194113
transform 1 0 82524 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1121_
timestamp 1607194113
transform 1 0 83076 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_66_907
timestamp 1607194113
transform 1 0 84548 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1607194113
transform 1 0 84364 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_931
timestamp 1607194113
transform 1 0 86756 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_919
timestamp 1607194113
transform 1 0 85652 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_713
timestamp 1607194113
transform 1 0 66700 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_705
timestamp 1607194113
transform 1 0 65964 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1607194113
transform 1 0 67160 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B1
timestamp 1607194113
transform 1 0 65780 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1607194113
transform 1 0 66884 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_738
timestamp 1607194113
transform 1 0 69000 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_733
timestamp 1607194113
transform 1 0 68540 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_720
timestamp 1607194113
transform 1 0 67344 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1607194113
transform 1 0 68448 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1607194113
transform 1 0 68724 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_750
timestamp 1607194113
transform 1 0 70104 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A1
timestamp 1607194113
transform 1 0 70840 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_778
timestamp 1607194113
transform 1 0 72680 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 1607194113
transform 1 0 72496 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A2
timestamp 1607194113
transform 1 0 72312 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1106_
timestamp 1607194113
transform 1 0 71024 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_67_794
timestamp 1607194113
transform 1 0 74152 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_785
timestamp 1607194113
transform 1 0 73324 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1607194113
transform 1 0 72864 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1607194113
transform 1 0 74060 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1607194113
transform 1 0 73048 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_818
timestamp 1607194113
transform 1 0 76360 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_806
timestamp 1607194113
transform 1 0 75256 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__CLK
timestamp 1607194113
transform 1 0 76912 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1464_
timestamp 1607194113
transform 1 0 77096 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_67_853
timestamp 1607194113
transform 1 0 79580 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_845
timestamp 1607194113
transform 1 0 78844 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1607194113
transform 1 0 79672 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1607194113
transform 1 0 79764 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_872
timestamp 1607194113
transform 1 0 81328 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_860
timestamp 1607194113
transform 1 0 80224 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1607194113
transform 1 0 80040 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_884
timestamp 1607194113
transform 1 0 82432 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1607194113
transform 1 0 83536 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0722_
timestamp 1607194113
transform 1 0 83168 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_907
timestamp 1607194113
transform 1 0 84548 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_898
timestamp 1607194113
transform 1 0 83720 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1607194113
transform 1 0 85284 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1607194113
transform 1 0 84272 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1607194113
transform 1 0 85376 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_925
timestamp 1607194113
transform 1 0 86204 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_919
timestamp 1607194113
transform 1 0 85652 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__CLK
timestamp 1607194113
transform 1 0 86296 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1460_
timestamp 1607194113
transform 1 0 86480 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_708
timestamp 1607194113
transform 1 0 66240 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_707
timestamp 1607194113
transform 1 0 66148 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_703
timestamp 1607194113
transform 1 0 65780 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_700
timestamp 1607194113
transform 1 0 65504 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__CLK
timestamp 1607194113
transform 1 0 66884 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1607194113
transform 1 0 65688 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1466_
timestamp 1607194113
transform 1 0 67068 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1607194113
transform 1 0 65872 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_733
timestamp 1607194113
transform 1 0 68540 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_720
timestamp 1607194113
transform 1 0 67344 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_736
timestamp 1607194113
transform 1 0 68816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1607194113
transform 1 0 68448 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_757
timestamp 1607194113
transform 1 0 70748 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_745
timestamp 1607194113
transform 1 0 69644 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_748
timestamp 1607194113
transform 1 0 69920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_765
timestamp 1607194113
transform 1 0 71484 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_761
timestamp 1607194113
transform 1 0 71116 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_760
timestamp 1607194113
transform 1 0 71024 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1607194113
transform 1 0 71392 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1607194113
transform 1 0 71300 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1607194113
transform 1 0 71208 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1095_
timestamp 1607194113
transform 1 0 71576 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_68_775
timestamp 1607194113
transform 1 0 72404 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B
timestamp 1607194113
transform 1 0 72220 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1104_
timestamp 1607194113
transform 1 0 72220 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_69_797
timestamp 1607194113
transform 1 0 74428 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_792
timestamp 1607194113
transform 1 0 73968 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_784
timestamp 1607194113
transform 1 0 73232 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_788
timestamp 1607194113
transform 1 0 73600 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1607194113
transform 1 0 73048 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1607194113
transform 1 0 72772 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1607194113
transform 1 0 74060 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1103_
timestamp 1607194113
transform 1 0 72956 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1607194113
transform 1 0 74152 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_809
timestamp 1607194113
transform 1 0 75532 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_812
timestamp 1607194113
transform 1 0 75808 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_800
timestamp 1607194113
transform 1 0 74704 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_833
timestamp 1607194113
transform 1 0 77740 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_821
timestamp 1607194113
transform 1 0 76636 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_825
timestamp 1607194113
transform 1 0 77004 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A
timestamp 1607194113
transform 1 0 77740 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1607194113
transform 1 0 76912 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1116_
timestamp 1607194113
transform 1 0 77924 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1087_
timestamp 1607194113
transform 1 0 77372 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_855
timestamp 1607194113
transform 1 0 79764 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_853
timestamp 1607194113
transform 1 0 79580 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_845
timestamp 1607194113
transform 1 0 78844 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_856
timestamp 1607194113
transform 1 0 79856 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_844
timestamp 1607194113
transform 1 0 78752 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1607194113
transform 1 0 79672 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_867
timestamp 1607194113
transform 1 0 80868 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_868
timestamp 1607194113
transform 1 0 80960 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_879
timestamp 1607194113
transform 1 0 81972 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_886
timestamp 1607194113
transform 1 0 82616 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_884
timestamp 1607194113
transform 1 0 82432 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_880
timestamp 1607194113
transform 1 0 82064 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1607194113
transform 1 0 82248 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A1
timestamp 1607194113
transform 1 0 83628 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1607194113
transform 1 0 82524 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1111_
timestamp 1607194113
transform 1 0 82432 0 1 39712
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_69_916
timestamp 1607194113
transform 1 0 85376 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_911
timestamp 1607194113
transform 1 0 84916 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_899
timestamp 1607194113
transform 1 0 83812 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_898
timestamp 1607194113
transform 1 0 83720 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__CLK
timestamp 1607194113
transform 1 0 83996 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1607194113
transform 1 0 85284 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1462_
timestamp 1607194113
transform 1 0 84180 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_928
timestamp 1607194113
transform 1 0 86480 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_922
timestamp 1607194113
transform 1 0 85928 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__CLK
timestamp 1607194113
transform 1 0 65504 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1607194113
transform 1 0 65688 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1471_
timestamp 1607194113
transform 1 0 65780 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_734
timestamp 1607194113
transform 1 0 68632 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_722
timestamp 1607194113
transform 1 0 67528 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_758
timestamp 1607194113
transform 1 0 70840 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_746
timestamp 1607194113
transform 1 0 69736 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_764
timestamp 1607194113
transform 1 0 71392 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_762
timestamp 1607194113
transform 1 0 71208 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__CLK
timestamp 1607194113
transform 1 0 71944 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1607194113
transform 1 0 71300 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1467_
timestamp 1607194113
transform 1 0 72128 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_791
timestamp 1607194113
transform 1 0 73876 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_815
timestamp 1607194113
transform 1 0 76084 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_803
timestamp 1607194113
transform 1 0 74980 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_836
timestamp 1607194113
transform 1 0 78016 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_825
timestamp 1607194113
transform 1 0 77004 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_823
timestamp 1607194113
transform 1 0 76820 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1607194113
transform 1 0 76912 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1097_
timestamp 1607194113
transform 1 0 77372 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_70_848
timestamp 1607194113
transform 1 0 79120 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_872
timestamp 1607194113
transform 1 0 81328 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_860
timestamp 1607194113
transform 1 0 80224 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_886
timestamp 1607194113
transform 1 0 82616 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_884
timestamp 1607194113
transform 1 0 82432 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1607194113
transform 1 0 82524 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1112_
timestamp 1607194113
transform 1 0 82708 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_910
timestamp 1607194113
transform 1 0 84824 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_901
timestamp 1607194113
transform 1 0 83996 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1607194113
transform 1 0 83812 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1607194113
transform 1 0 84548 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_922
timestamp 1607194113
transform 1 0 85928 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_703
timestamp 1607194113
transform 1 0 65780 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1607194113
transform 1 0 65596 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1607194113
transform 1 0 67160 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1092_
timestamp 1607194113
transform 1 0 66332 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_733
timestamp 1607194113
transform 1 0 68540 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_720
timestamp 1607194113
transform 1 0 67344 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1607194113
transform 1 0 68448 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_757
timestamp 1607194113
transform 1 0 70748 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_745
timestamp 1607194113
transform 1 0 69644 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_765
timestamp 1607194113
transform 1 0 71484 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1607194113
transform 1 0 71760 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1035_
timestamp 1607194113
transform 1 0 71944 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_794
timestamp 1607194113
transform 1 0 74152 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_781
timestamp 1607194113
transform 1 0 72956 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__D
timestamp 1607194113
transform 1 0 72772 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1607194113
transform 1 0 74060 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_814
timestamp 1607194113
transform 1 0 75992 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_806
timestamp 1607194113
transform 1 0 75256 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1607194113
transform 1 0 76176 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_836
timestamp 1607194113
transform 1 0 78016 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_821
timestamp 1607194113
transform 1 0 76636 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1607194113
transform 1 0 76452 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1100_
timestamp 1607194113
transform 1 0 77188 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_855
timestamp 1607194113
transform 1 0 79764 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_848
timestamp 1607194113
transform 1 0 79120 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1607194113
transform 1 0 79672 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_867
timestamp 1607194113
transform 1 0 80868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_896
timestamp 1607194113
transform 1 0 83536 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_887
timestamp 1607194113
transform 1 0 82708 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_879
timestamp 1607194113
transform 1 0 81972 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1607194113
transform 1 0 83352 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0709_
timestamp 1607194113
transform 1 0 82984 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_916
timestamp 1607194113
transform 1 0 85376 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_914
timestamp 1607194113
transform 1 0 85192 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_908
timestamp 1607194113
transform 1 0 84640 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1607194113
transform 1 0 85284 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_928
timestamp 1607194113
transform 1 0 86480 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_711
timestamp 1607194113
transform 1 0 66516 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_703
timestamp 1607194113
transform 1 0 65780 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_701
timestamp 1607194113
transform 1 0 65596 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1607194113
transform 1 0 65688 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1091_
timestamp 1607194113
transform 1 0 66608 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_72_731
timestamp 1607194113
transform 1 0 68356 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_719
timestamp 1607194113
transform 1 0 67252 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_755
timestamp 1607194113
transform 1 0 70564 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_743
timestamp 1607194113
transform 1 0 69460 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_772
timestamp 1607194113
transform 1 0 72128 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_764
timestamp 1607194113
transform 1 0 71392 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1607194113
transform 1 0 71300 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1096_
timestamp 1607194113
transform 1 0 72312 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_72_793
timestamp 1607194113
transform 1 0 74060 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_781
timestamp 1607194113
transform 1 0 72956 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_818
timestamp 1607194113
transform 1 0 76360 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_811
timestamp 1607194113
transform 1 0 75716 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_805
timestamp 1607194113
transform 1 0 75164 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1607194113
transform 1 0 76176 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0779_
timestamp 1607194113
transform 1 0 75808 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_825
timestamp 1607194113
transform 1 0 77004 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__CLK
timestamp 1607194113
transform 1 0 77372 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1607194113
transform 1 0 76912 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1468_
timestamp 1607194113
transform 1 0 77556 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_850
timestamp 1607194113
transform 1 0 79304 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_874
timestamp 1607194113
transform 1 0 81512 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_862
timestamp 1607194113
transform 1 0 80408 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_886
timestamp 1607194113
transform 1 0 82616 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_72_882
timestamp 1607194113
transform 1 0 82248 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__CLK
timestamp 1607194113
transform 1 0 83168 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1607194113
transform 1 0 82524 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1465_
timestamp 1607194113
transform 1 0 83352 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_913
timestamp 1607194113
transform 1 0 85100 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_925
timestamp 1607194113
transform 1 0 86204 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_707
timestamp 1607194113
transform 1 0 66148 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1088_
timestamp 1607194113
transform 1 0 66884 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_73_733
timestamp 1607194113
transform 1 0 68540 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_724
timestamp 1607194113
transform 1 0 67712 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1607194113
transform 1 0 68448 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1083_
timestamp 1607194113
transform 1 0 68632 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_73_753
timestamp 1607194113
transform 1 0 70380 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_741
timestamp 1607194113
transform 1 0 69276 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1607194113
transform 1 0 70656 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_778
timestamp 1607194113
transform 1 0 72680 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_767
timestamp 1607194113
transform 1 0 71668 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_759
timestamp 1607194113
transform 1 0 70932 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1607194113
transform 1 0 72496 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1081_
timestamp 1607194113
transform 1 0 71852 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_73_794
timestamp 1607194113
transform 1 0 74152 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_790
timestamp 1607194113
transform 1 0 73784 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1607194113
transform 1 0 74060 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_818
timestamp 1607194113
transform 1 0 76360 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_806
timestamp 1607194113
transform 1 0 75256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_830
timestamp 1607194113
transform 1 0 77464 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1101_
timestamp 1607194113
transform 1 0 77556 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_73_855
timestamp 1607194113
transform 1 0 79764 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_842
timestamp 1607194113
transform 1 0 78568 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A
timestamp 1607194113
transform 1 0 78384 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1607194113
transform 1 0 79672 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_867
timestamp 1607194113
transform 1 0 80868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_891
timestamp 1607194113
transform 1 0 83076 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_879
timestamp 1607194113
transform 1 0 81972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_916
timestamp 1607194113
transform 1 0 85376 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_903
timestamp 1607194113
transform 1 0 84180 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1607194113
transform 1 0 85284 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_928
timestamp 1607194113
transform 1 0 86480 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_712
timestamp 1607194113
transform 1 0 66608 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_708
timestamp 1607194113
transform 1 0 66240 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_718
timestamp 1607194113
transform 1 0 67160 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_703
timestamp 1607194113
transform 1 0 65780 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1607194113
transform 1 0 66976 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1607194113
transform 1 0 65688 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1089_
timestamp 1607194113
transform 1 0 66148 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1084_
timestamp 1607194113
transform 1 0 66700 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_75_733
timestamp 1607194113
transform 1 0 68540 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_720
timestamp 1607194113
transform 1 0 67344 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_734
timestamp 1607194113
transform 1 0 68632 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_730
timestamp 1607194113
transform 1 0 68264 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__D
timestamp 1607194113
transform 1 0 68724 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1607194113
transform 1 0 68448 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1038_
timestamp 1607194113
transform 1 0 68908 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_75_757
timestamp 1607194113
transform 1 0 70748 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_745
timestamp 1607194113
transform 1 0 69644 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_758
timestamp 1607194113
transform 1 0 70840 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_746
timestamp 1607194113
transform 1 0 69736 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_772
timestamp 1607194113
transform 1 0 72128 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_762
timestamp 1607194113
transform 1 0 71208 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1607194113
transform 1 0 72680 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__C
timestamp 1607194113
transform 1 0 71944 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1607194113
transform 1 0 71300 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1093_
timestamp 1607194113
transform 1 0 71392 0 -1 42976
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1049_
timestamp 1607194113
transform 1 0 71116 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1607194113
transform 1 0 72680 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_794
timestamp 1607194113
transform 1 0 74152 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_791
timestamp 1607194113
transform 1 0 73876 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_783
timestamp 1607194113
transform 1 0 73140 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_792
timestamp 1607194113
transform 1 0 73968 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_780
timestamp 1607194113
transform 1 0 72864 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1607194113
transform 1 0 72956 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1607194113
transform 1 0 74060 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_818
timestamp 1607194113
transform 1 0 76360 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_806
timestamp 1607194113
transform 1 0 75256 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_816
timestamp 1607194113
transform 1 0 76176 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_804
timestamp 1607194113
transform 1 0 75072 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_826
timestamp 1607194113
transform 1 0 77096 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_825
timestamp 1607194113
transform 1 0 77004 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1607194113
transform 1 0 77372 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A1
timestamp 1607194113
transform 1 0 77556 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1607194113
transform 1 0 77372 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1607194113
transform 1 0 76912 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1099_
timestamp 1607194113
transform 1 0 77556 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _1098_
timestamp 1607194113
transform 1 0 77740 0 -1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_75_855
timestamp 1607194113
transform 1 0 79764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_851
timestamp 1607194113
transform 1 0 79396 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_843
timestamp 1607194113
transform 1 0 78660 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_857
timestamp 1607194113
transform 1 0 79948 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_846
timestamp 1607194113
transform 1 0 78936 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1607194113
transform 1 0 79672 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1607194113
transform 1 0 79672 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_867
timestamp 1607194113
transform 1 0 80868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_869
timestamp 1607194113
transform 1 0 81052 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_891
timestamp 1607194113
transform 1 0 83076 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_879
timestamp 1607194113
transform 1 0 81972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_886
timestamp 1607194113
transform 1 0 82616 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_881
timestamp 1607194113
transform 1 0 82156 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1607194113
transform 1 0 82524 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_916
timestamp 1607194113
transform 1 0 85376 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_903
timestamp 1607194113
transform 1 0 84180 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_910
timestamp 1607194113
transform 1 0 84824 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_898
timestamp 1607194113
transform 1 0 83720 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1607194113
transform 1 0 85284 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_928
timestamp 1607194113
transform 1 0 86480 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_922
timestamp 1607194113
transform 1 0 85928 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_703
timestamp 1607194113
transform 1 0 65780 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_700
timestamp 1607194113
transform 1 0 65504 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1607194113
transform 1 0 65964 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1607194113
transform 1 0 65688 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1086_
timestamp 1607194113
transform 1 0 66148 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_731
timestamp 1607194113
transform 1 0 68356 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_719
timestamp 1607194113
transform 1 0 67252 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_755
timestamp 1607194113
transform 1 0 70564 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_743
timestamp 1607194113
transform 1 0 69460 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_771
timestamp 1607194113
transform 1 0 72036 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1607194113
transform 1 0 71300 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1607194113
transform 1 0 71392 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_76_794
timestamp 1607194113
transform 1 0 74152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_782
timestamp 1607194113
transform 1 0 73048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1607194113
transform 1 0 72772 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_818
timestamp 1607194113
transform 1 0 76360 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_806
timestamp 1607194113
transform 1 0 75256 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_825
timestamp 1607194113
transform 1 0 77004 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__CLK
timestamp 1607194113
transform 1 0 77372 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1607194113
transform 1 0 76912 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1469_
timestamp 1607194113
transform 1 0 77556 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_76_850
timestamp 1607194113
transform 1 0 79304 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_874
timestamp 1607194113
transform 1 0 81512 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_862
timestamp 1607194113
transform 1 0 80408 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_886
timestamp 1607194113
transform 1 0 82616 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_882
timestamp 1607194113
transform 1 0 82248 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1607194113
transform 1 0 82524 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_910
timestamp 1607194113
transform 1 0 84824 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_898
timestamp 1607194113
transform 1 0 83720 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_922
timestamp 1607194113
transform 1 0 85928 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_701
timestamp 1607194113
transform 1 0 65596 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A1
timestamp 1607194113
transform 1 0 65964 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1085_
timestamp 1607194113
transform 1 0 66148 0 1 44064
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_77_736
timestamp 1607194113
transform 1 0 68816 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_730
timestamp 1607194113
transform 1 0 68264 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_722
timestamp 1607194113
transform 1 0 67528 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B1
timestamp 1607194113
transform 1 0 67344 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1607194113
transform 1 0 68448 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1607194113
transform 1 0 68540 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_748
timestamp 1607194113
transform 1 0 69920 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_760
timestamp 1607194113
transform 1 0 71024 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1470_
timestamp 1607194113
transform 1 0 71392 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_77_794
timestamp 1607194113
transform 1 0 74152 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_785
timestamp 1607194113
transform 1 0 73324 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__CLK
timestamp 1607194113
transform 1 0 73140 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1607194113
transform 1 0 74060 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_818
timestamp 1607194113
transform 1 0 76360 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_806
timestamp 1607194113
transform 1 0 75256 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_830
timestamp 1607194113
transform 1 0 77464 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_855
timestamp 1607194113
transform 1 0 79764 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_842
timestamp 1607194113
transform 1 0 78568 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1607194113
transform 1 0 79672 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_867
timestamp 1607194113
transform 1 0 80868 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_891
timestamp 1607194113
transform 1 0 83076 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_879
timestamp 1607194113
transform 1 0 81972 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_916
timestamp 1607194113
transform 1 0 85376 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_903
timestamp 1607194113
transform 1 0 84180 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1607194113
transform 1 0 85284 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_928
timestamp 1607194113
transform 1 0 86480 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_703
timestamp 1607194113
transform 1 0 65780 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_701
timestamp 1607194113
transform 1 0 65596 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__CLK
timestamp 1607194113
transform 1 0 66516 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1607194113
transform 1 0 65688 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1473_
timestamp 1607194113
transform 1 0 66700 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_78_732
timestamp 1607194113
transform 1 0 68448 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_756
timestamp 1607194113
transform 1 0 70656 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_744
timestamp 1607194113
transform 1 0 69552 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_776
timestamp 1607194113
transform 1 0 72496 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_764
timestamp 1607194113
transform 1 0 71392 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_762
timestamp 1607194113
transform 1 0 71208 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1607194113
transform 1 0 71300 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_788
timestamp 1607194113
transform 1 0 73600 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_812
timestamp 1607194113
transform 1 0 75808 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_800
timestamp 1607194113
transform 1 0 74704 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_837
timestamp 1607194113
transform 1 0 78108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_825
timestamp 1607194113
transform 1 0 77004 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1607194113
transform 1 0 76912 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_849
timestamp 1607194113
transform 1 0 79212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_873
timestamp 1607194113
transform 1 0 81420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_861
timestamp 1607194113
transform 1 0 80316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_886
timestamp 1607194113
transform 1 0 82616 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1607194113
transform 1 0 82524 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_910
timestamp 1607194113
transform 1 0 84824 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_898
timestamp 1607194113
transform 1 0 83720 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_922
timestamp 1607194113
transform 1 0 85928 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_708
timestamp 1607194113
transform 1 0 66240 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_733
timestamp 1607194113
transform 1 0 68540 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_720
timestamp 1607194113
transform 1 0 67344 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1607194113
transform 1 0 68448 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_757
timestamp 1607194113
transform 1 0 70748 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_745
timestamp 1607194113
transform 1 0 69644 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_769
timestamp 1607194113
transform 1 0 71852 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_794
timestamp 1607194113
transform 1 0 74152 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_781
timestamp 1607194113
transform 1 0 72956 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1607194113
transform 1 0 74060 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_818
timestamp 1607194113
transform 1 0 76360 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_806
timestamp 1607194113
transform 1 0 75256 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_830
timestamp 1607194113
transform 1 0 77464 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_855
timestamp 1607194113
transform 1 0 79764 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_842
timestamp 1607194113
transform 1 0 78568 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1607194113
transform 1 0 79672 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_867
timestamp 1607194113
transform 1 0 80868 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_891
timestamp 1607194113
transform 1 0 83076 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_879
timestamp 1607194113
transform 1 0 81972 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_916
timestamp 1607194113
transform 1 0 85376 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_903
timestamp 1607194113
transform 1 0 84180 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1607194113
transform 1 0 85284 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_928
timestamp 1607194113
transform 1 0 86480 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_947
timestamp 1607194113
transform 1 0 88228 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_942
timestamp 1607194113
transform 1 0 87768 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[8]
timestamp 1607194113
transform 1 0 87584 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[7]
timestamp 1607194113
transform 1 0 87400 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[6]
timestamp 1607194113
transform 1 0 87216 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[5]
timestamp 1607194113
transform 1 0 87032 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607194113
transform 1 0 88136 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_971
timestamp 1607194113
transform 1 0 90436 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_959
timestamp 1607194113
transform 1 0 89332 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_983
timestamp 1607194113
transform 1 0 91540 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1008
timestamp 1607194113
transform 1 0 93840 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_995
timestamp 1607194113
transform 1 0 92644 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607194113
transform 1 0 93748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1020
timestamp 1607194113
transform 1 0 94944 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1044
timestamp 1607194113
transform 1 0 97152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1032
timestamp 1607194113
transform 1 0 96048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1069
timestamp 1607194113
transform 1 0 99452 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1056
timestamp 1607194113
transform 1 0 98256 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607194113
transform 1 0 99360 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1081
timestamp 1607194113
transform 1 0 100556 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1105
timestamp 1607194113
transform 1 0 102764 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1093
timestamp 1607194113
transform 1 0 101660 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1130
timestamp 1607194113
transform 1 0 105064 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1117
timestamp 1607194113
transform 1 0 103868 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607194113
transform 1 0 104972 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1142
timestamp 1607194113
transform 1 0 106168 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1158
timestamp 1607194113
transform 1 0 107640 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_1154
timestamp 1607194113
transform 1 0 107272 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607194113
transform -1 0 108008 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_943
timestamp 1607194113
transform 1 0 87860 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_936
timestamp 1607194113
transform 1 0 87216 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[3]
timestamp 1607194113
transform 1 0 87032 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1607194113
transform 1 0 87584 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_967
timestamp 1607194113
transform 1 0 90068 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_955
timestamp 1607194113
transform 1 0 88964 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_989
timestamp 1607194113
transform 1 0 92092 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_977
timestamp 1607194113
transform 1 0 90988 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_975
timestamp 1607194113
transform 1 0 90804 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607194113
transform 1 0 90896 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1001
timestamp 1607194113
transform 1 0 93196 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1025
timestamp 1607194113
transform 1 0 95404 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1013
timestamp 1607194113
transform 1 0 94300 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1050
timestamp 1607194113
transform 1 0 97704 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1038
timestamp 1607194113
transform 1 0 96600 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607194113
transform 1 0 96508 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1062
timestamp 1607194113
transform 1 0 98808 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1086
timestamp 1607194113
transform 1 0 101016 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1074
timestamp 1607194113
transform 1 0 99912 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1099
timestamp 1607194113
transform 1 0 102212 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607194113
transform 1 0 102120 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1123
timestamp 1607194113
transform 1 0 104420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1111
timestamp 1607194113
transform 1 0 103316 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1147
timestamp 1607194113
transform 1 0 106628 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1135
timestamp 1607194113
transform 1 0 105524 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607194113
transform -1 0 108008 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_947
timestamp 1607194113
transform 1 0 88228 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_942
timestamp 1607194113
transform 1 0 87768 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_934
timestamp 1607194113
transform 1 0 87032 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__CLK
timestamp 1607194113
transform 1 0 87952 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607194113
transform 1 0 88136 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1607194113
transform 1 0 88320 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_52_967
timestamp 1607194113
transform 1 0 90068 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_991
timestamp 1607194113
transform 1 0 92276 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_979
timestamp 1607194113
transform 1 0 91172 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1008
timestamp 1607194113
transform 1 0 93840 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_1003
timestamp 1607194113
transform 1 0 93380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607194113
transform 1 0 93748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1020
timestamp 1607194113
transform 1 0 94944 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1044
timestamp 1607194113
transform 1 0 97152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1032
timestamp 1607194113
transform 1 0 96048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1069
timestamp 1607194113
transform 1 0 99452 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1056
timestamp 1607194113
transform 1 0 98256 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607194113
transform 1 0 99360 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1081
timestamp 1607194113
transform 1 0 100556 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1105
timestamp 1607194113
transform 1 0 102764 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1093
timestamp 1607194113
transform 1 0 101660 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1130
timestamp 1607194113
transform 1 0 105064 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1117
timestamp 1607194113
transform 1 0 103868 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607194113
transform 1 0 104972 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1142
timestamp 1607194113
transform 1 0 106168 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1158
timestamp 1607194113
transform 1 0 107640 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_1154
timestamp 1607194113
transform 1 0 107272 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607194113
transform -1 0 108008 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_947
timestamp 1607194113
transform 1 0 88228 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_933
timestamp 1607194113
transform 1 0 86940 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1607194113
transform 1 0 87216 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1146_
timestamp 1607194113
transform 1 0 87400 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_971
timestamp 1607194113
transform 1 0 90436 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_959
timestamp 1607194113
transform 1 0 89332 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_989
timestamp 1607194113
transform 1 0 92092 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_977
timestamp 1607194113
transform 1 0 90988 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_975
timestamp 1607194113
transform 1 0 90804 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607194113
transform 1 0 90896 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1001
timestamp 1607194113
transform 1 0 93196 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1025
timestamp 1607194113
transform 1 0 95404 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1013
timestamp 1607194113
transform 1 0 94300 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1050
timestamp 1607194113
transform 1 0 97704 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1038
timestamp 1607194113
transform 1 0 96600 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607194113
transform 1 0 96508 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1062
timestamp 1607194113
transform 1 0 98808 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1086
timestamp 1607194113
transform 1 0 101016 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1074
timestamp 1607194113
transform 1 0 99912 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1099
timestamp 1607194113
transform 1 0 102212 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607194113
transform 1 0 102120 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1123
timestamp 1607194113
transform 1 0 104420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1111
timestamp 1607194113
transform 1 0 103316 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1147
timestamp 1607194113
transform 1 0 106628 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1135
timestamp 1607194113
transform 1 0 105524 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607194113
transform -1 0 108008 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_951
timestamp 1607194113
transform 1 0 88596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_940
timestamp 1607194113
transform 1 0 87584 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1607194113
transform 1 0 87400 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607194113
transform 1 0 88136 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1607194113
transform 1 0 88228 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_963
timestamp 1607194113
transform 1 0 89700 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_987
timestamp 1607194113
transform 1 0 91908 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_975
timestamp 1607194113
transform 1 0 90804 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1008
timestamp 1607194113
transform 1 0 93840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_999
timestamp 1607194113
transform 1 0 93012 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607194113
transform 1 0 93748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1020
timestamp 1607194113
transform 1 0 94944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1044
timestamp 1607194113
transform 1 0 97152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1032
timestamp 1607194113
transform 1 0 96048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1069
timestamp 1607194113
transform 1 0 99452 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1056
timestamp 1607194113
transform 1 0 98256 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607194113
transform 1 0 99360 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1081
timestamp 1607194113
transform 1 0 100556 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1105
timestamp 1607194113
transform 1 0 102764 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1093
timestamp 1607194113
transform 1 0 101660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1130
timestamp 1607194113
transform 1 0 105064 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1117
timestamp 1607194113
transform 1 0 103868 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607194113
transform 1 0 104972 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1142
timestamp 1607194113
transform 1 0 106168 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1158
timestamp 1607194113
transform 1 0 107640 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_1154
timestamp 1607194113
transform 1 0 107272 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607194113
transform -1 0 108008 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_945
timestamp 1607194113
transform 1 0 88044 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_933
timestamp 1607194113
transform 1 0 86940 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_940
timestamp 1607194113
transform 1 0 87584 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607194113
transform 1 0 88136 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1132_
timestamp 1607194113
transform 1 0 88228 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_56_968
timestamp 1607194113
transform 1 0 90160 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_956
timestamp 1607194113
transform 1 0 89056 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_964
timestamp 1607194113
transform 1 0 89792 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_952
timestamp 1607194113
transform 1 0 88688 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1607194113
transform 1 0 88872 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_980
timestamp 1607194113
transform 1 0 91264 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_989
timestamp 1607194113
transform 1 0 92092 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_977
timestamp 1607194113
transform 1 0 90988 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607194113
transform 1 0 90896 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1008
timestamp 1607194113
transform 1 0 93840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_1004
timestamp 1607194113
transform 1 0 93472 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_992
timestamp 1607194113
transform 1 0 92368 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1001
timestamp 1607194113
transform 1 0 93196 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607194113
transform 1 0 93748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1020
timestamp 1607194113
transform 1 0 94944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1025
timestamp 1607194113
transform 1 0 95404 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1013
timestamp 1607194113
transform 1 0 94300 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1044
timestamp 1607194113
transform 1 0 97152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1032
timestamp 1607194113
transform 1 0 96048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1050
timestamp 1607194113
transform 1 0 97704 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1038
timestamp 1607194113
transform 1 0 96600 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607194113
transform 1 0 96508 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1069
timestamp 1607194113
transform 1 0 99452 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1056
timestamp 1607194113
transform 1 0 98256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1062
timestamp 1607194113
transform 1 0 98808 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607194113
transform 1 0 99360 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1081
timestamp 1607194113
transform 1 0 100556 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1086
timestamp 1607194113
transform 1 0 101016 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1074
timestamp 1607194113
transform 1 0 99912 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1105
timestamp 1607194113
transform 1 0 102764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1093
timestamp 1607194113
transform 1 0 101660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1099
timestamp 1607194113
transform 1 0 102212 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607194113
transform 1 0 102120 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1130
timestamp 1607194113
transform 1 0 105064 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1117
timestamp 1607194113
transform 1 0 103868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1123
timestamp 1607194113
transform 1 0 104420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1111
timestamp 1607194113
transform 1 0 103316 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607194113
transform 1 0 104972 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1142
timestamp 1607194113
transform 1 0 106168 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1147
timestamp 1607194113
transform 1 0 106628 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1135
timestamp 1607194113
transform 1 0 105524 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1158
timestamp 1607194113
transform 1 0 107640 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_1154
timestamp 1607194113
transform 1 0 107272 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607194113
transform -1 0 108008 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607194113
transform -1 0 108008 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_944
timestamp 1607194113
transform 1 0 87952 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_938
timestamp 1607194113
transform 1 0 87400 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__CLK
timestamp 1607194113
transform 1 0 88044 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1459_
timestamp 1607194113
transform 1 0 88228 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_966
timestamp 1607194113
transform 1 0 89976 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_989
timestamp 1607194113
transform 1 0 92092 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_977
timestamp 1607194113
transform 1 0 90988 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_974
timestamp 1607194113
transform 1 0 90712 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607194113
transform 1 0 90896 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1001
timestamp 1607194113
transform 1 0 93196 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1025
timestamp 1607194113
transform 1 0 95404 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1013
timestamp 1607194113
transform 1 0 94300 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1050
timestamp 1607194113
transform 1 0 97704 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1038
timestamp 1607194113
transform 1 0 96600 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607194113
transform 1 0 96508 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1062
timestamp 1607194113
transform 1 0 98808 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1086
timestamp 1607194113
transform 1 0 101016 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1074
timestamp 1607194113
transform 1 0 99912 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1099
timestamp 1607194113
transform 1 0 102212 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607194113
transform 1 0 102120 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1123
timestamp 1607194113
transform 1 0 104420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1111
timestamp 1607194113
transform 1 0 103316 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1147
timestamp 1607194113
transform 1 0 106628 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1135
timestamp 1607194113
transform 1 0 105524 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607194113
transform -1 0 108008 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_938
timestamp 1607194113
transform 1 0 87400 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_933
timestamp 1607194113
transform 1 0 86940 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1607194113
transform 1 0 87952 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607194113
transform 1 0 88136 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1134_
timestamp 1607194113
transform 1 0 88228 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1607194113
transform 1 0 87124 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_968
timestamp 1607194113
transform 1 0 90160 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_956
timestamp 1607194113
transform 1 0 89056 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0729_
timestamp 1607194113
transform 1 0 89792 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_980
timestamp 1607194113
transform 1 0 91264 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1008
timestamp 1607194113
transform 1 0 93840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_1004
timestamp 1607194113
transform 1 0 93472 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_992
timestamp 1607194113
transform 1 0 92368 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607194113
transform 1 0 93748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1020
timestamp 1607194113
transform 1 0 94944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1044
timestamp 1607194113
transform 1 0 97152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1032
timestamp 1607194113
transform 1 0 96048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1069
timestamp 1607194113
transform 1 0 99452 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1056
timestamp 1607194113
transform 1 0 98256 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607194113
transform 1 0 99360 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1081
timestamp 1607194113
transform 1 0 100556 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1105
timestamp 1607194113
transform 1 0 102764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1093
timestamp 1607194113
transform 1 0 101660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1130
timestamp 1607194113
transform 1 0 105064 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1117
timestamp 1607194113
transform 1 0 103868 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607194113
transform 1 0 104972 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1142
timestamp 1607194113
transform 1 0 106168 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1158
timestamp 1607194113
transform 1 0 107640 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1154
timestamp 1607194113
transform 1 0 107272 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607194113
transform -1 0 108008 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_951
timestamp 1607194113
transform 1 0 88596 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_943
timestamp 1607194113
transform 1 0 87860 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1133_
timestamp 1607194113
transform 1 0 87952 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_59_962
timestamp 1607194113
transform 1 0 89608 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1607194113
transform 1 0 89332 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_989
timestamp 1607194113
transform 1 0 92092 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_977
timestamp 1607194113
transform 1 0 90988 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_974
timestamp 1607194113
transform 1 0 90712 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607194113
transform 1 0 90896 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1001
timestamp 1607194113
transform 1 0 93196 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1025
timestamp 1607194113
transform 1 0 95404 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1013
timestamp 1607194113
transform 1 0 94300 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1050
timestamp 1607194113
transform 1 0 97704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1038
timestamp 1607194113
transform 1 0 96600 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607194113
transform 1 0 96508 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1062
timestamp 1607194113
transform 1 0 98808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1086
timestamp 1607194113
transform 1 0 101016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1074
timestamp 1607194113
transform 1 0 99912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1099
timestamp 1607194113
transform 1 0 102212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607194113
transform 1 0 102120 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1123
timestamp 1607194113
transform 1 0 104420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1111
timestamp 1607194113
transform 1 0 103316 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1147
timestamp 1607194113
transform 1 0 106628 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1135
timestamp 1607194113
transform 1 0 105524 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607194113
transform -1 0 108008 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_950
timestamp 1607194113
transform 1 0 88504 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_934
timestamp 1607194113
transform 1 0 87032 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1607194113
transform 1 0 88136 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1607194113
transform 1 0 88228 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_962
timestamp 1607194113
transform 1 0 89608 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_986
timestamp 1607194113
transform 1 0 91816 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_974
timestamp 1607194113
transform 1 0 90712 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1008
timestamp 1607194113
transform 1 0 93840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1006
timestamp 1607194113
transform 1 0 93656 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_998
timestamp 1607194113
transform 1 0 92920 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1607194113
transform 1 0 93748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1020
timestamp 1607194113
transform 1 0 94944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1044
timestamp 1607194113
transform 1 0 97152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1032
timestamp 1607194113
transform 1 0 96048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1069
timestamp 1607194113
transform 1 0 99452 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1056
timestamp 1607194113
transform 1 0 98256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1607194113
transform 1 0 99360 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1081
timestamp 1607194113
transform 1 0 100556 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1105
timestamp 1607194113
transform 1 0 102764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1093
timestamp 1607194113
transform 1 0 101660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1130
timestamp 1607194113
transform 1 0 105064 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1117
timestamp 1607194113
transform 1 0 103868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1607194113
transform 1 0 104972 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1142
timestamp 1607194113
transform 1 0 106168 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1158
timestamp 1607194113
transform 1 0 107640 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1154
timestamp 1607194113
transform 1 0 107272 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607194113
transform -1 0 108008 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_938
timestamp 1607194113
transform 1 0 87400 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_939
timestamp 1607194113
transform 1 0 87492 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__CLK
timestamp 1607194113
transform 1 0 88228 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1607194113
transform 1 0 88504 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1607194113
transform 1 0 88136 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1461_
timestamp 1607194113
transform 1 0 88412 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1125_
timestamp 1607194113
transform 1 0 87860 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_968
timestamp 1607194113
transform 1 0 90160 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_964
timestamp 1607194113
transform 1 0 89792 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_952
timestamp 1607194113
transform 1 0 88688 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_980
timestamp 1607194113
transform 1 0 91264 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_989
timestamp 1607194113
transform 1 0 92092 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_977
timestamp 1607194113
transform 1 0 90988 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1607194113
transform 1 0 90896 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1008
timestamp 1607194113
transform 1 0 93840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1004
timestamp 1607194113
transform 1 0 93472 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_992
timestamp 1607194113
transform 1 0 92368 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1001
timestamp 1607194113
transform 1 0 93196 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1607194113
transform 1 0 93748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1020
timestamp 1607194113
transform 1 0 94944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1025
timestamp 1607194113
transform 1 0 95404 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1013
timestamp 1607194113
transform 1 0 94300 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1044
timestamp 1607194113
transform 1 0 97152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1032
timestamp 1607194113
transform 1 0 96048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1050
timestamp 1607194113
transform 1 0 97704 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1038
timestamp 1607194113
transform 1 0 96600 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1607194113
transform 1 0 96508 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1069
timestamp 1607194113
transform 1 0 99452 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1056
timestamp 1607194113
transform 1 0 98256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1062
timestamp 1607194113
transform 1 0 98808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1607194113
transform 1 0 99360 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1081
timestamp 1607194113
transform 1 0 100556 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1086
timestamp 1607194113
transform 1 0 101016 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1074
timestamp 1607194113
transform 1 0 99912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1105
timestamp 1607194113
transform 1 0 102764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1093
timestamp 1607194113
transform 1 0 101660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1099
timestamp 1607194113
transform 1 0 102212 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1607194113
transform 1 0 102120 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1130
timestamp 1607194113
transform 1 0 105064 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1117
timestamp 1607194113
transform 1 0 103868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1123
timestamp 1607194113
transform 1 0 104420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1111
timestamp 1607194113
transform 1 0 103316 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1607194113
transform 1 0 104972 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1142
timestamp 1607194113
transform 1 0 106168 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1147
timestamp 1607194113
transform 1 0 106628 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1135
timestamp 1607194113
transform 1 0 105524 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1158
timestamp 1607194113
transform 1 0 107640 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1154
timestamp 1607194113
transform 1 0 107272 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607194113
transform -1 0 108008 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607194113
transform -1 0 108008 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_938
timestamp 1607194113
transform 1 0 87400 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1607194113
transform 1 0 87952 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1127_
timestamp 1607194113
transform 1 0 88136 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_967
timestamp 1607194113
transform 1 0 90068 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_955
timestamp 1607194113
transform 1 0 88964 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_989
timestamp 1607194113
transform 1 0 92092 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_977
timestamp 1607194113
transform 1 0 90988 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_975
timestamp 1607194113
transform 1 0 90804 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1607194113
transform 1 0 90896 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1001
timestamp 1607194113
transform 1 0 93196 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1025
timestamp 1607194113
transform 1 0 95404 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1013
timestamp 1607194113
transform 1 0 94300 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1050
timestamp 1607194113
transform 1 0 97704 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1038
timestamp 1607194113
transform 1 0 96600 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1607194113
transform 1 0 96508 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1062
timestamp 1607194113
transform 1 0 98808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1086
timestamp 1607194113
transform 1 0 101016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1074
timestamp 1607194113
transform 1 0 99912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1099
timestamp 1607194113
transform 1 0 102212 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1607194113
transform 1 0 102120 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1123
timestamp 1607194113
transform 1 0 104420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1111
timestamp 1607194113
transform 1 0 103316 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1147
timestamp 1607194113
transform 1 0 106628 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1135
timestamp 1607194113
transform 1 0 105524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607194113
transform -1 0 108008 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_942
timestamp 1607194113
transform 1 0 87768 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1607194113
transform 1 0 88136 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1126_
timestamp 1607194113
transform 1 0 88228 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_64_968
timestamp 1607194113
transform 1 0 90160 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_956
timestamp 1607194113
transform 1 0 89056 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1607194113
transform 1 0 88872 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_980
timestamp 1607194113
transform 1 0 91264 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1008
timestamp 1607194113
transform 1 0 93840 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1004
timestamp 1607194113
transform 1 0 93472 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_992
timestamp 1607194113
transform 1 0 92368 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1607194113
transform 1 0 93748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1020
timestamp 1607194113
transform 1 0 94944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1044
timestamp 1607194113
transform 1 0 97152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1032
timestamp 1607194113
transform 1 0 96048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1069
timestamp 1607194113
transform 1 0 99452 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1056
timestamp 1607194113
transform 1 0 98256 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1607194113
transform 1 0 99360 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1081
timestamp 1607194113
transform 1 0 100556 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1105
timestamp 1607194113
transform 1 0 102764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1093
timestamp 1607194113
transform 1 0 101660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1130
timestamp 1607194113
transform 1 0 105064 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1117
timestamp 1607194113
transform 1 0 103868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1607194113
transform 1 0 104972 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1142
timestamp 1607194113
transform 1 0 106168 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1158
timestamp 1607194113
transform 1 0 107640 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1154
timestamp 1607194113
transform 1 0 107272 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607194113
transform -1 0 108008 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_944
timestamp 1607194113
transform 1 0 87952 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_968
timestamp 1607194113
transform 1 0 90160 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_956
timestamp 1607194113
transform 1 0 89056 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_989
timestamp 1607194113
transform 1 0 92092 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_977
timestamp 1607194113
transform 1 0 90988 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1607194113
transform 1 0 90896 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1001
timestamp 1607194113
transform 1 0 93196 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1025
timestamp 1607194113
transform 1 0 95404 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1013
timestamp 1607194113
transform 1 0 94300 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1050
timestamp 1607194113
transform 1 0 97704 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1038
timestamp 1607194113
transform 1 0 96600 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1607194113
transform 1 0 96508 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1062
timestamp 1607194113
transform 1 0 98808 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1086
timestamp 1607194113
transform 1 0 101016 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1074
timestamp 1607194113
transform 1 0 99912 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1099
timestamp 1607194113
transform 1 0 102212 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1607194113
transform 1 0 102120 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1123
timestamp 1607194113
transform 1 0 104420 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1111
timestamp 1607194113
transform 1 0 103316 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1147
timestamp 1607194113
transform 1 0 106628 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1135
timestamp 1607194113
transform 1 0 105524 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607194113
transform -1 0 108008 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_947
timestamp 1607194113
transform 1 0 88228 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_943
timestamp 1607194113
transform 1 0 87860 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1607194113
transform 1 0 88136 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_971
timestamp 1607194113
transform 1 0 90436 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_959
timestamp 1607194113
transform 1 0 89332 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_983
timestamp 1607194113
transform 1 0 91540 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1008
timestamp 1607194113
transform 1 0 93840 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_995
timestamp 1607194113
transform 1 0 92644 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1607194113
transform 1 0 93748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1020
timestamp 1607194113
transform 1 0 94944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1044
timestamp 1607194113
transform 1 0 97152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1032
timestamp 1607194113
transform 1 0 96048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1069
timestamp 1607194113
transform 1 0 99452 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1056
timestamp 1607194113
transform 1 0 98256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1607194113
transform 1 0 99360 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1081
timestamp 1607194113
transform 1 0 100556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1105
timestamp 1607194113
transform 1 0 102764 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1093
timestamp 1607194113
transform 1 0 101660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1130
timestamp 1607194113
transform 1 0 105064 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1117
timestamp 1607194113
transform 1 0 103868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1607194113
transform 1 0 104972 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1142
timestamp 1607194113
transform 1 0 106168 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1158
timestamp 1607194113
transform 1 0 107640 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_1154
timestamp 1607194113
transform 1 0 107272 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607194113
transform -1 0 108008 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_947
timestamp 1607194113
transform 1 0 88228 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_971
timestamp 1607194113
transform 1 0 90436 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_959
timestamp 1607194113
transform 1 0 89332 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_989
timestamp 1607194113
transform 1 0 92092 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_977
timestamp 1607194113
transform 1 0 90988 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_975
timestamp 1607194113
transform 1 0 90804 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1607194113
transform 1 0 90896 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1001
timestamp 1607194113
transform 1 0 93196 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1025
timestamp 1607194113
transform 1 0 95404 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1013
timestamp 1607194113
transform 1 0 94300 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1050
timestamp 1607194113
transform 1 0 97704 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1038
timestamp 1607194113
transform 1 0 96600 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1607194113
transform 1 0 96508 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1062
timestamp 1607194113
transform 1 0 98808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1086
timestamp 1607194113
transform 1 0 101016 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1074
timestamp 1607194113
transform 1 0 99912 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1099
timestamp 1607194113
transform 1 0 102212 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1607194113
transform 1 0 102120 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1123
timestamp 1607194113
transform 1 0 104420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1111
timestamp 1607194113
transform 1 0 103316 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1147
timestamp 1607194113
transform 1 0 106628 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1135
timestamp 1607194113
transform 1 0 105524 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607194113
transform -1 0 108008 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_940
timestamp 1607194113
transform 1 0 87584 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_947
timestamp 1607194113
transform 1 0 88228 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_934
timestamp 1607194113
transform 1 0 87032 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1607194113
transform 1 0 88136 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_964
timestamp 1607194113
transform 1 0 89792 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_952
timestamp 1607194113
transform 1 0 88688 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_971
timestamp 1607194113
transform 1 0 90436 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_959
timestamp 1607194113
transform 1 0 89332 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_989
timestamp 1607194113
transform 1 0 92092 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_977
timestamp 1607194113
transform 1 0 90988 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_983
timestamp 1607194113
transform 1 0 91540 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1607194113
transform 1 0 90896 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1001
timestamp 1607194113
transform 1 0 93196 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1008
timestamp 1607194113
transform 1 0 93840 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_995
timestamp 1607194113
transform 1 0 92644 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1607194113
transform 1 0 93748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1025
timestamp 1607194113
transform 1 0 95404 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1013
timestamp 1607194113
transform 1 0 94300 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1020
timestamp 1607194113
transform 1 0 94944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1050
timestamp 1607194113
transform 1 0 97704 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1038
timestamp 1607194113
transform 1 0 96600 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1044
timestamp 1607194113
transform 1 0 97152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1032
timestamp 1607194113
transform 1 0 96048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1607194113
transform 1 0 96508 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1062
timestamp 1607194113
transform 1 0 98808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1069
timestamp 1607194113
transform 1 0 99452 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1056
timestamp 1607194113
transform 1 0 98256 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1607194113
transform 1 0 99360 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1086
timestamp 1607194113
transform 1 0 101016 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1074
timestamp 1607194113
transform 1 0 99912 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1081
timestamp 1607194113
transform 1 0 100556 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1099
timestamp 1607194113
transform 1 0 102212 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1105
timestamp 1607194113
transform 1 0 102764 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1093
timestamp 1607194113
transform 1 0 101660 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1607194113
transform 1 0 102120 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1123
timestamp 1607194113
transform 1 0 104420 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1111
timestamp 1607194113
transform 1 0 103316 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1130
timestamp 1607194113
transform 1 0 105064 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1117
timestamp 1607194113
transform 1 0 103868 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1607194113
transform 1 0 104972 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1147
timestamp 1607194113
transform 1 0 106628 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1135
timestamp 1607194113
transform 1 0 105524 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1142
timestamp 1607194113
transform 1 0 106168 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1158
timestamp 1607194113
transform 1 0 107640 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_1154
timestamp 1607194113
transform 1 0 107272 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607194113
transform -1 0 108008 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607194113
transform -1 0 108008 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_947
timestamp 1607194113
transform 1 0 88228 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_934
timestamp 1607194113
transform 1 0 87032 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1607194113
transform 1 0 88136 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_971
timestamp 1607194113
transform 1 0 90436 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_959
timestamp 1607194113
transform 1 0 89332 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_983
timestamp 1607194113
transform 1 0 91540 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1008
timestamp 1607194113
transform 1 0 93840 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_995
timestamp 1607194113
transform 1 0 92644 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1607194113
transform 1 0 93748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1020
timestamp 1607194113
transform 1 0 94944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1044
timestamp 1607194113
transform 1 0 97152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1032
timestamp 1607194113
transform 1 0 96048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1069
timestamp 1607194113
transform 1 0 99452 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1056
timestamp 1607194113
transform 1 0 98256 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1607194113
transform 1 0 99360 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1081
timestamp 1607194113
transform 1 0 100556 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1105
timestamp 1607194113
transform 1 0 102764 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1093
timestamp 1607194113
transform 1 0 101660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1130
timestamp 1607194113
transform 1 0 105064 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1117
timestamp 1607194113
transform 1 0 103868 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1607194113
transform 1 0 104972 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1142
timestamp 1607194113
transform 1 0 106168 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1158
timestamp 1607194113
transform 1 0 107640 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_1154
timestamp 1607194113
transform 1 0 107272 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607194113
transform -1 0 108008 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_940
timestamp 1607194113
transform 1 0 87584 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_964
timestamp 1607194113
transform 1 0 89792 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_952
timestamp 1607194113
transform 1 0 88688 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_989
timestamp 1607194113
transform 1 0 92092 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_977
timestamp 1607194113
transform 1 0 90988 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1607194113
transform 1 0 90896 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1001
timestamp 1607194113
transform 1 0 93196 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1025
timestamp 1607194113
transform 1 0 95404 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1013
timestamp 1607194113
transform 1 0 94300 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1050
timestamp 1607194113
transform 1 0 97704 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1038
timestamp 1607194113
transform 1 0 96600 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1607194113
transform 1 0 96508 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1062
timestamp 1607194113
transform 1 0 98808 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1086
timestamp 1607194113
transform 1 0 101016 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1074
timestamp 1607194113
transform 1 0 99912 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1099
timestamp 1607194113
transform 1 0 102212 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1607194113
transform 1 0 102120 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1123
timestamp 1607194113
transform 1 0 104420 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1111
timestamp 1607194113
transform 1 0 103316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1147
timestamp 1607194113
transform 1 0 106628 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1135
timestamp 1607194113
transform 1 0 105524 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607194113
transform -1 0 108008 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_947
timestamp 1607194113
transform 1 0 88228 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_945
timestamp 1607194113
transform 1 0 88044 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_937
timestamp 1607194113
transform 1 0 87308 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1607194113
transform 1 0 88136 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_971
timestamp 1607194113
transform 1 0 90436 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_959
timestamp 1607194113
transform 1 0 89332 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_983
timestamp 1607194113
transform 1 0 91540 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1008
timestamp 1607194113
transform 1 0 93840 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_995
timestamp 1607194113
transform 1 0 92644 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1607194113
transform 1 0 93748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1020
timestamp 1607194113
transform 1 0 94944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1044
timestamp 1607194113
transform 1 0 97152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1032
timestamp 1607194113
transform 1 0 96048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1069
timestamp 1607194113
transform 1 0 99452 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1056
timestamp 1607194113
transform 1 0 98256 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1607194113
transform 1 0 99360 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1081
timestamp 1607194113
transform 1 0 100556 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1105
timestamp 1607194113
transform 1 0 102764 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1093
timestamp 1607194113
transform 1 0 101660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1130
timestamp 1607194113
transform 1 0 105064 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1117
timestamp 1607194113
transform 1 0 103868 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1607194113
transform 1 0 104972 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1142
timestamp 1607194113
transform 1 0 106168 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1158
timestamp 1607194113
transform 1 0 107640 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_1154
timestamp 1607194113
transform 1 0 107272 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607194113
transform -1 0 108008 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_940
timestamp 1607194113
transform 1 0 87584 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_964
timestamp 1607194113
transform 1 0 89792 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_952
timestamp 1607194113
transform 1 0 88688 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_989
timestamp 1607194113
transform 1 0 92092 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_977
timestamp 1607194113
transform 1 0 90988 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1607194113
transform 1 0 90896 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1001
timestamp 1607194113
transform 1 0 93196 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1025
timestamp 1607194113
transform 1 0 95404 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1013
timestamp 1607194113
transform 1 0 94300 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1050
timestamp 1607194113
transform 1 0 97704 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1038
timestamp 1607194113
transform 1 0 96600 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1607194113
transform 1 0 96508 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1062
timestamp 1607194113
transform 1 0 98808 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1086
timestamp 1607194113
transform 1 0 101016 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1074
timestamp 1607194113
transform 1 0 99912 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1099
timestamp 1607194113
transform 1 0 102212 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1607194113
transform 1 0 102120 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1123
timestamp 1607194113
transform 1 0 104420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1111
timestamp 1607194113
transform 1 0 103316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1147
timestamp 1607194113
transform 1 0 106628 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1135
timestamp 1607194113
transform 1 0 105524 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607194113
transform -1 0 108008 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_940
timestamp 1607194113
transform 1 0 87584 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_947
timestamp 1607194113
transform 1 0 88228 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_934
timestamp 1607194113
transform 1 0 87032 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1607194113
transform 1 0 88136 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_964
timestamp 1607194113
transform 1 0 89792 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_952
timestamp 1607194113
transform 1 0 88688 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_971
timestamp 1607194113
transform 1 0 90436 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_959
timestamp 1607194113
transform 1 0 89332 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_989
timestamp 1607194113
transform 1 0 92092 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_977
timestamp 1607194113
transform 1 0 90988 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_983
timestamp 1607194113
transform 1 0 91540 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1607194113
transform 1 0 90896 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1001
timestamp 1607194113
transform 1 0 93196 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1008
timestamp 1607194113
transform 1 0 93840 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_995
timestamp 1607194113
transform 1 0 92644 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1607194113
transform 1 0 93748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1025
timestamp 1607194113
transform 1 0 95404 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1013
timestamp 1607194113
transform 1 0 94300 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1020
timestamp 1607194113
transform 1 0 94944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1050
timestamp 1607194113
transform 1 0 97704 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1038
timestamp 1607194113
transform 1 0 96600 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1044
timestamp 1607194113
transform 1 0 97152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1032
timestamp 1607194113
transform 1 0 96048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1607194113
transform 1 0 96508 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1062
timestamp 1607194113
transform 1 0 98808 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1069
timestamp 1607194113
transform 1 0 99452 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1056
timestamp 1607194113
transform 1 0 98256 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1607194113
transform 1 0 99360 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1086
timestamp 1607194113
transform 1 0 101016 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1074
timestamp 1607194113
transform 1 0 99912 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1081
timestamp 1607194113
transform 1 0 100556 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1099
timestamp 1607194113
transform 1 0 102212 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1105
timestamp 1607194113
transform 1 0 102764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1093
timestamp 1607194113
transform 1 0 101660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1607194113
transform 1 0 102120 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1123
timestamp 1607194113
transform 1 0 104420 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1111
timestamp 1607194113
transform 1 0 103316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1130
timestamp 1607194113
transform 1 0 105064 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1117
timestamp 1607194113
transform 1 0 103868 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1607194113
transform 1 0 104972 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1147
timestamp 1607194113
transform 1 0 106628 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1135
timestamp 1607194113
transform 1 0 105524 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1142
timestamp 1607194113
transform 1 0 106168 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1158
timestamp 1607194113
transform 1 0 107640 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_1154
timestamp 1607194113
transform 1 0 107272 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607194113
transform -1 0 108008 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607194113
transform -1 0 108008 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_947
timestamp 1607194113
transform 1 0 88228 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_934
timestamp 1607194113
transform 1 0 87032 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1607194113
transform 1 0 88136 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_971
timestamp 1607194113
transform 1 0 90436 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_959
timestamp 1607194113
transform 1 0 89332 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_983
timestamp 1607194113
transform 1 0 91540 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1008
timestamp 1607194113
transform 1 0 93840 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_995
timestamp 1607194113
transform 1 0 92644 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1607194113
transform 1 0 93748 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1020
timestamp 1607194113
transform 1 0 94944 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1044
timestamp 1607194113
transform 1 0 97152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1032
timestamp 1607194113
transform 1 0 96048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1069
timestamp 1607194113
transform 1 0 99452 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1056
timestamp 1607194113
transform 1 0 98256 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1607194113
transform 1 0 99360 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1081
timestamp 1607194113
transform 1 0 100556 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1105
timestamp 1607194113
transform 1 0 102764 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1093
timestamp 1607194113
transform 1 0 101660 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1130
timestamp 1607194113
transform 1 0 105064 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1117
timestamp 1607194113
transform 1 0 103868 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1607194113
transform 1 0 104972 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1142
timestamp 1607194113
transform 1 0 106168 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1158
timestamp 1607194113
transform 1 0 107640 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_1154
timestamp 1607194113
transform 1 0 107272 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607194113
transform -1 0 108008 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_940
timestamp 1607194113
transform 1 0 87584 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_964
timestamp 1607194113
transform 1 0 89792 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_952
timestamp 1607194113
transform 1 0 88688 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_989
timestamp 1607194113
transform 1 0 92092 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_977
timestamp 1607194113
transform 1 0 90988 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1607194113
transform 1 0 90896 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1001
timestamp 1607194113
transform 1 0 93196 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1025
timestamp 1607194113
transform 1 0 95404 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1013
timestamp 1607194113
transform 1 0 94300 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1050
timestamp 1607194113
transform 1 0 97704 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1038
timestamp 1607194113
transform 1 0 96600 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1607194113
transform 1 0 96508 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1062
timestamp 1607194113
transform 1 0 98808 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1086
timestamp 1607194113
transform 1 0 101016 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1074
timestamp 1607194113
transform 1 0 99912 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1099
timestamp 1607194113
transform 1 0 102212 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1607194113
transform 1 0 102120 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1123
timestamp 1607194113
transform 1 0 104420 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1111
timestamp 1607194113
transform 1 0 103316 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1147
timestamp 1607194113
transform 1 0 106628 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_1135
timestamp 1607194113
transform 1 0 105524 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607194113
transform -1 0 108008 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_947
timestamp 1607194113
transform 1 0 88228 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_934
timestamp 1607194113
transform 1 0 87032 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1607194113
transform 1 0 88136 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_971
timestamp 1607194113
transform 1 0 90436 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_959
timestamp 1607194113
transform 1 0 89332 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_983
timestamp 1607194113
transform 1 0 91540 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1008
timestamp 1607194113
transform 1 0 93840 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_995
timestamp 1607194113
transform 1 0 92644 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1607194113
transform 1 0 93748 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1020
timestamp 1607194113
transform 1 0 94944 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1044
timestamp 1607194113
transform 1 0 97152 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1032
timestamp 1607194113
transform 1 0 96048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1069
timestamp 1607194113
transform 1 0 99452 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1056
timestamp 1607194113
transform 1 0 98256 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1607194113
transform 1 0 99360 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1081
timestamp 1607194113
transform 1 0 100556 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1105
timestamp 1607194113
transform 1 0 102764 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1093
timestamp 1607194113
transform 1 0 101660 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1130
timestamp 1607194113
transform 1 0 105064 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1117
timestamp 1607194113
transform 1 0 103868 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1607194113
transform 1 0 104972 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_1142
timestamp 1607194113
transform 1 0 106168 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_1158
timestamp 1607194113
transform 1 0 107640 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_1154
timestamp 1607194113
transform 1 0 107272 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1607194113
transform -1 0 108008 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_940
timestamp 1607194113
transform 1 0 87584 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_964
timestamp 1607194113
transform 1 0 89792 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_952
timestamp 1607194113
transform 1 0 88688 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_989
timestamp 1607194113
transform 1 0 92092 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_977
timestamp 1607194113
transform 1 0 90988 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1607194113
transform 1 0 90896 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1001
timestamp 1607194113
transform 1 0 93196 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1025
timestamp 1607194113
transform 1 0 95404 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1013
timestamp 1607194113
transform 1 0 94300 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1050
timestamp 1607194113
transform 1 0 97704 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1038
timestamp 1607194113
transform 1 0 96600 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1607194113
transform 1 0 96508 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1062
timestamp 1607194113
transform 1 0 98808 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1086
timestamp 1607194113
transform 1 0 101016 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1074
timestamp 1607194113
transform 1 0 99912 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1099
timestamp 1607194113
transform 1 0 102212 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1607194113
transform 1 0 102120 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1123
timestamp 1607194113
transform 1 0 104420 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1111
timestamp 1607194113
transform 1 0 103316 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1147
timestamp 1607194113
transform 1 0 106628 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_1135
timestamp 1607194113
transform 1 0 105524 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1607194113
transform -1 0 108008 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1607194113
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1607194113
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1607194113
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_81_11
timestamp 1607194113
transform 1 0 2116 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_3
timestamp 1607194113
transform 1 0 1380 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__D
timestamp 1607194113
transform 1 0 2392 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1607194113
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1345_
timestamp 1607194113
transform 1 0 2576 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1607194113
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1607194113
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1607194113
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_32
timestamp 1607194113
transform 1 0 4048 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1607194113
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_37
timestamp 1607194113
transform 1 0 4508 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1607194113
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_27
timestamp 1607194113
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__CLK
timestamp 1607194113
transform 1 0 4324 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1607194113
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1607194113
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1512_
timestamp 1607194113
transform 1 0 4232 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_82_55
timestamp 1607194113
transform 1 0 6164 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_49
timestamp 1607194113
transform 1 0 5612 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1607194113
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1607194113
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__CLK
timestamp 1607194113
transform 1 0 5980 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1607194113
transform 1 0 7268 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_66
timestamp 1607194113
transform 1 0 7176 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_62
timestamp 1607194113
transform 1 0 6808 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_68
timestamp 1607194113
transform 1 0 7360 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1607194113
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1510_
timestamp 1607194113
transform 1 0 7268 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _0877_
timestamp 1607194113
transform 1 0 7912 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0875_
timestamp 1607194113
transform 1 0 7636 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_80_93
timestamp 1607194113
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_91
timestamp 1607194113
transform 1 0 9476 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_83
timestamp 1607194113
transform 1 0 8740 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1607194113
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_88
timestamp 1607194113
transform 1 0 9200 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__CLK
timestamp 1607194113
transform 1 0 9016 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1607194113
transform 1 0 9660 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_90
timestamp 1607194113
transform 1 0 9384 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_82
timestamp 1607194113
transform 1 0 8648 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B
timestamp 1607194113
transform 1 0 8464 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1607194113
transform 1 0 9568 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_117
timestamp 1607194113
transform 1 0 11868 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_105
timestamp 1607194113
transform 1 0 10764 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_112
timestamp 1607194113
transform 1 0 11408 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_100
timestamp 1607194113
transform 1 0 10304 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_117
timestamp 1607194113
transform 1 0 11868 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_105
timestamp 1607194113
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B1
timestamp 1607194113
transform 1 0 12052 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_120
timestamp 1607194113
transform 1 0 12144 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_137
timestamp 1607194113
transform 1 0 13708 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_129
timestamp 1607194113
transform 1 0 12972 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A1_N
timestamp 1607194113
transform 1 0 13708 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1607194113
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1395_
timestamp 1607194113
transform 1 0 12420 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1244_
timestamp 1607194113
transform 1 0 12236 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_154
timestamp 1607194113
transform 1 0 15272 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_150
timestamp 1607194113
transform 1 0 14904 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_142
timestamp 1607194113
transform 1 0 14168 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1607194113
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1607194113
transform 1 0 13892 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_156
timestamp 1607194113
transform 1 0 15456 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_144
timestamp 1607194113
transform 1 0 14352 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__CLK
timestamp 1607194113
transform 1 0 14168 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_154
timestamp 1607194113
transform 1 0 15272 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_151
timestamp 1607194113
transform 1 0 14996 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_143
timestamp 1607194113
transform 1 0 14260 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A2_N
timestamp 1607194113
transform 1 0 14076 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B2
timestamp 1607194113
transform 1 0 13892 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1607194113
transform 1 0 15180 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_166
timestamp 1607194113
transform 1 0 16376 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_168
timestamp 1607194113
transform 1 0 16560 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_166
timestamp 1607194113
transform 1 0 16376 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__CLK
timestamp 1607194113
transform 1 0 16928 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B1
timestamp 1607194113
transform 1 0 16652 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1396_
timestamp 1607194113
transform 1 0 17112 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1243_
timestamp 1607194113
transform 1 0 16836 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_193
timestamp 1607194113
transform 1 0 18860 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A2_N
timestamp 1607194113
transform 1 0 18676 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B2
timestamp 1607194113
transform 1 0 18492 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A1_N
timestamp 1607194113
transform 1 0 18308 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_198
timestamp 1607194113
transform 1 0 19320 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_187
timestamp 1607194113
transform 1 0 18308 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_180
timestamp 1607194113
transform 1 0 17664 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1607194113
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1607194113
transform 1 0 19044 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1607194113
transform 1 0 18032 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_193
timestamp 1607194113
transform 1 0 18860 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_211
timestamp 1607194113
transform 1 0 20516 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_205
timestamp 1607194113
transform 1 0 19964 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B1
timestamp 1607194113
transform 1 0 20608 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1607194113
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0876_
timestamp 1607194113
transform 1 0 20884 0 -1 46240
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1607194113
transform 1 0 19872 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0878_
timestamp 1607194113
transform 1 0 20056 0 1 46240
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_82_215
timestamp 1607194113
transform 1 0 20884 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_213
timestamp 1607194113
transform 1 0 20700 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_205
timestamp 1607194113
transform 1 0 19964 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1607194113
transform 1 0 20792 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_231
timestamp 1607194113
transform 1 0 22356 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_227
timestamp 1607194113
transform 1 0 21988 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_222
timestamp 1607194113
transform 1 0 21528 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_231
timestamp 1607194113
transform 1 0 22356 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1607194113
transform 1 0 21344 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A1
timestamp 1607194113
transform 1 0 22172 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B1
timestamp 1607194113
transform 1 0 22448 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1607194113
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1607194113
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1607194113
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_32
timestamp 1607194113
transform 1 0 4048 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_27
timestamp 1607194113
transform 1 0 3588 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1607194113
transform 1 0 3956 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_56
timestamp 1607194113
transform 1 0 6256 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_44
timestamp 1607194113
transform 1 0 5152 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_71
timestamp 1607194113
transform 1 0 7636 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_63
timestamp 1607194113
transform 1 0 6900 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1607194113
transform 1 0 6808 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0879_
timestamp 1607194113
transform 1 0 7912 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_83_94
timestamp 1607194113
transform 1 0 9752 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_91
timestamp 1607194113
transform 1 0 9476 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_83
timestamp 1607194113
transform 1 0 8740 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1607194113
transform 1 0 9660 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_118
timestamp 1607194113
transform 1 0 11960 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_106
timestamp 1607194113
transform 1 0 10856 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_137
timestamp 1607194113
transform 1 0 13708 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_125
timestamp 1607194113
transform 1 0 12604 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1607194113
transform 1 0 12512 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_156
timestamp 1607194113
transform 1 0 15456 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_149
timestamp 1607194113
transform 1 0 14812 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1607194113
transform 1 0 15364 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_168
timestamp 1607194113
transform 1 0 16560 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_187
timestamp 1607194113
transform 1 0 18308 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_180
timestamp 1607194113
transform 1 0 17664 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1607194113
transform 1 0 18216 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_218
timestamp 1607194113
transform 1 0 21160 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_211
timestamp 1607194113
transform 1 0 20516 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_199
timestamp 1607194113
transform 1 0 19412 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1607194113
transform 1 0 21068 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_230
timestamp 1607194113
transform 1 0 22264 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_243
timestamp 1607194113
transform 1 0 23460 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B1
timestamp 1607194113
transform 1 0 23552 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1179_
timestamp 1607194113
transform 1 0 23736 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_81_245
timestamp 1607194113
transform 1 0 23644 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_242
timestamp 1607194113
transform 1 0 23368 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_234
timestamp 1607194113
transform 1 0 22632 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__CLK
timestamp 1607194113
transform 1 0 23736 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1607194113
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1436_
timestamp 1607194113
transform 1 0 23920 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_82_252
timestamp 1607194113
transform 1 0 24288 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1_N
timestamp 1607194113
transform 1 0 24104 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1180_
timestamp 1607194113
transform 1 0 22632 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_82_267
timestamp 1607194113
transform 1 0 25668 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_81_267
timestamp 1607194113
transform 1 0 25668 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_80_272
timestamp 1607194113
transform 1 0 26128 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_264
timestamp 1607194113
transform 1 0 25392 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1_N
timestamp 1607194113
transform 1 0 25208 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1607194113
transform 1 0 25392 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_288
timestamp 1607194113
transform 1 0 27600 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_276
timestamp 1607194113
transform 1 0 26496 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_285
timestamp 1607194113
transform 1 0 27324 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_276
timestamp 1607194113
transform 1 0 26496 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__CLK
timestamp 1607194113
transform 1 0 26220 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1607194113
transform 1 0 26404 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1607194113
transform 1 0 26404 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1437_
timestamp 1607194113
transform 1 0 26404 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1607194113
transform 1 0 27048 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_311
timestamp 1607194113
transform 1 0 29716 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1607194113
transform 1 0 29532 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1607194113
transform 1 0 29348 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0874_
timestamp 1607194113
transform 1 0 28060 0 -1 46240
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_81_306
timestamp 1607194113
transform 1 0 29256 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_302
timestamp 1607194113
transform 1 0 28888 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_294
timestamp 1607194113
transform 1 0 28152 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1607194113
transform 1 0 29164 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_312
timestamp 1607194113
transform 1 0 29808 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_300
timestamp 1607194113
transform 1 0 28704 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_324
timestamp 1607194113
transform 1 0 30912 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_318
timestamp 1607194113
transform 1 0 30360 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_323
timestamp 1607194113
transform 1 0 30820 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B1
timestamp 1607194113
transform 1 0 30912 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1178_
timestamp 1607194113
transform 1 0 31096 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_80_337
timestamp 1607194113
transform 1 0 32108 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_335
timestamp 1607194113
transform 1 0 31924 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1607194113
transform 1 0 32016 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1438_
timestamp 1607194113
transform 1 0 32844 0 -1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_81_352
timestamp 1607194113
transform 1 0 33488 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_344
timestamp 1607194113
transform 1 0 32752 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A1_N
timestamp 1607194113
transform 1 0 32568 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_341
timestamp 1607194113
transform 1 0 32476 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_337
timestamp 1607194113
transform 1 0 32108 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1607194113
transform 1 0 32016 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1397_
timestamp 1607194113
transform 1 0 32568 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_82_363
timestamp 1607194113
transform 1 0 34500 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1607194113
transform 1 0 35144 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_358
timestamp 1607194113
transform 1 0 34040 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_366
timestamp 1607194113
transform 1 0 34776 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__CLK
timestamp 1607194113
transform 1 0 34592 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1607194113
transform 1 0 34316 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1607194113
transform 1 0 34776 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1607194113
transform 1 0 33764 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1607194113
transform 1 0 34868 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_387
timestamp 1607194113
transform 1 0 36708 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_375
timestamp 1607194113
transform 1 0 35604 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_390
timestamp 1607194113
transform 1 0 36984 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1607194113
transform 1 0 36248 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_390
timestamp 1607194113
transform 1 0 36984 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_378
timestamp 1607194113
transform 1 0 35880 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A1_N
timestamp 1607194113
transform 1 0 37260 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B1
timestamp 1607194113
transform 1 0 37444 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1607194113
transform 1 0 37628 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0718_
timestamp 1607194113
transform 1 0 37720 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1_N
timestamp 1607194113
transform 1 0 37260 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B1
timestamp 1607194113
transform 1 0 37444 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0813_
timestamp 1607194113
transform 1 0 37628 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_82_406
timestamp 1607194113
transform 1 0 38456 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_398
timestamp 1607194113
transform 1 0 37720 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_395
timestamp 1607194113
transform 1 0 37444 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__CLK
timestamp 1607194113
transform 1 0 38732 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1607194113
transform 1 0 37628 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1607194113
transform 1 0 38916 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_80_430
timestamp 1607194113
transform 1 0 40664 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_418
timestamp 1607194113
transform 1 0 39560 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A2_N
timestamp 1607194113
transform 1 0 39376 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B2
timestamp 1607194113
transform 1 0 39192 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_431
timestamp 1607194113
transform 1 0 40756 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_425
timestamp 1607194113
transform 1 0 40204 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_417
timestamp 1607194113
transform 1 0 39468 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A2_N
timestamp 1607194113
transform 1 0 39284 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B2
timestamp 1607194113
transform 1 0 39100 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1607194113
transform 1 0 40388 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1607194113
transform 1 0 40480 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_430
timestamp 1607194113
transform 1 0 40664 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_442
timestamp 1607194113
transform 1 0 41768 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_443
timestamp 1607194113
transform 1 0 41860 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_442
timestamp 1607194113
transform 1 0 41768 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__CLK
timestamp 1607194113
transform 1 0 42044 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1480_
timestamp 1607194113
transform 1 0 42228 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_82_462
timestamp 1607194113
transform 1 0 43608 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_454
timestamp 1607194113
transform 1 0 42872 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_466
timestamp 1607194113
transform 1 0 43976 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_459
timestamp 1607194113
transform 1 0 43332 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_454
timestamp 1607194113
transform 1 0 42872 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1607194113
transform 1 0 43240 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1607194113
transform 1 0 43240 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1607194113
transform 1 0 43332 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_249
timestamp 1607194113
transform 1 0 24012 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_242
timestamp 1607194113
transform 1 0 23368 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1607194113
transform 1 0 23920 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_261
timestamp 1607194113
transform 1 0 25116 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_292
timestamp 1607194113
transform 1 0 27968 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_280
timestamp 1607194113
transform 1 0 26864 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1607194113
transform 1 0 26220 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1607194113
transform 1 0 26772 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_311
timestamp 1607194113
transform 1 0 29716 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_304
timestamp 1607194113
transform 1 0 29072 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1607194113
transform 1 0 29624 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_323
timestamp 1607194113
transform 1 0 30820 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_342
timestamp 1607194113
transform 1 0 32568 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_335
timestamp 1607194113
transform 1 0 31924 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1607194113
transform 1 0 32476 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_366
timestamp 1607194113
transform 1 0 34776 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_354
timestamp 1607194113
transform 1 0 33672 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1607194113
transform 1 0 35328 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_385
timestamp 1607194113
transform 1 0 36524 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_373
timestamp 1607194113
transform 1 0 35420 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_404
timestamp 1607194113
transform 1 0 38272 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_397
timestamp 1607194113
transform 1 0 37628 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1607194113
transform 1 0 38180 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_428
timestamp 1607194113
transform 1 0 40480 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_416
timestamp 1607194113
transform 1 0 39376 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_447
timestamp 1607194113
transform 1 0 42228 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_435
timestamp 1607194113
transform 1 0 41124 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1607194113
transform 1 0 41032 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_466
timestamp 1607194113
transform 1 0 43976 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_459
timestamp 1607194113
transform 1 0 43332 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1607194113
transform 1 0 43884 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_474
timestamp 1607194113
transform 1 0 44712 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_478
timestamp 1607194113
transform 1 0 45080 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_467
timestamp 1607194113
transform 1 0 44068 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A1
timestamp 1607194113
transform 1 0 45632 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1066_
timestamp 1607194113
transform 1 0 44896 0 -1 47328
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _1059_
timestamp 1607194113
transform 1 0 44344 0 -1 46240
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_80_503
timestamp 1607194113
transform 1 0 47380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_488
timestamp 1607194113
transform 1 0 46000 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B1
timestamp 1607194113
transform 1 0 45816 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__C
timestamp 1607194113
transform 1 0 47196 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1051_
timestamp 1607194113
transform 1 0 46368 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_81_498
timestamp 1607194113
transform 1 0 46920 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_81_486
timestamp 1607194113
transform 1 0 45816 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1607194113
transform 1 0 46736 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1607194113
transform 1 0 46000 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1607194113
transform 1 0 47472 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1052_
timestamp 1607194113
transform 1 0 46092 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_82_494
timestamp 1607194113
transform 1 0 46552 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1607194113
transform 1 0 46368 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B
timestamp 1607194113
transform 1 0 47564 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A2
timestamp 1607194113
transform 1 0 46184 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1061_
timestamp 1607194113
transform 1 0 46920 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_80_520
timestamp 1607194113
transform 1 0 48944 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_515
timestamp 1607194113
transform 1 0 48484 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1607194113
transform 1 0 48852 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_522
timestamp 1607194113
transform 1 0 49128 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_507
timestamp 1607194113
transform 1 0 47748 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1064_
timestamp 1607194113
transform 1 0 48484 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_82_524
timestamp 1607194113
transform 1 0 49312 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_520
timestamp 1607194113
transform 1 0 48944 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_507
timestamp 1607194113
transform 1 0 47748 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1607194113
transform 1 0 48852 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1607194113
transform 1 0 49404 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_532
timestamp 1607194113
transform 1 0 50048 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1_N
timestamp 1607194113
transform 1 0 50600 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1607194113
transform 1 0 50784 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0767_
timestamp 1607194113
transform 1 0 50968 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_81_538
timestamp 1607194113
transform 1 0 50600 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_530
timestamp 1607194113
transform 1 0 49864 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1063_
timestamp 1607194113
transform 1 0 49956 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_82_536
timestamp 1607194113
transform 1 0 50416 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_528
timestamp 1607194113
transform 1 0 49680 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1065_
timestamp 1607194113
transform 1 0 50600 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_82_559
timestamp 1607194113
transform 1 0 52532 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_549
timestamp 1607194113
transform 1 0 51612 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_546
timestamp 1607194113
transform 1 0 51336 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_558
timestamp 1607194113
transform 1 0 52440 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__CLK
timestamp 1607194113
transform 1 0 51428 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1607194113
transform 1 0 51428 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1607194113
transform 1 0 51612 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1607194113
transform 1 0 51704 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0766_
timestamp 1607194113
transform 1 0 52164 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_581
timestamp 1607194113
transform 1 0 54556 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_578
timestamp 1607194113
transform 1 0 54280 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_570
timestamp 1607194113
transform 1 0 53544 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1607194113
transform 1 0 54464 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_581
timestamp 1607194113
transform 1 0 54556 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_569
timestamp 1607194113
transform 1 0 53452 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1607194113
transform 1 0 54832 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_581
timestamp 1607194113
transform 1 0 54556 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_579
timestamp 1607194113
transform 1 0 54372 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_571
timestamp 1607194113
transform 1 0 53636 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1607194113
transform 1 0 54464 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_601
timestamp 1607194113
transform 1 0 56396 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_593
timestamp 1607194113
transform 1 0 55660 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_81_604
timestamp 1607194113
transform 1 0 56672 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_587
timestamp 1607194113
transform 1 0 55108 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_600
timestamp 1607194113
transform 1 0 56304 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1607194113
transform 1 0 56488 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1056_
timestamp 1607194113
transform 1 0 56488 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1055_
timestamp 1607194113
transform 1 0 55660 0 -1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1054_
timestamp 1607194113
transform 1 0 55844 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_82_613
timestamp 1607194113
transform 1 0 57500 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_624
timestamp 1607194113
transform 1 0 58512 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_612
timestamp 1607194113
transform 1 0 57408 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1607194113
transform 1 0 57316 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1607194113
transform 1 0 57224 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1481_
timestamp 1607194113
transform 1 0 57316 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_80_642
timestamp 1607194113
transform 1 0 60168 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_640
timestamp 1607194113
transform 1 0 59984 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_636
timestamp 1607194113
transform 1 0 59616 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1607194113
transform 1 0 60076 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_644
timestamp 1607194113
transform 1 0 60352 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_632
timestamp 1607194113
transform 1 0 59248 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__CLK
timestamp 1607194113
transform 1 0 59064 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_642
timestamp 1607194113
transform 1 0 60168 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_637
timestamp 1607194113
transform 1 0 59708 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_625
timestamp 1607194113
transform 1 0 58604 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1607194113
transform 1 0 60076 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_650
timestamp 1607194113
transform 1 0 60904 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_664
timestamp 1607194113
transform 1 0 62192 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_81_656
timestamp 1607194113
transform 1 0 61456 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_658
timestamp 1607194113
transform 1 0 61640 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_654
timestamp 1607194113
transform 1 0 61272 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1607194113
transform 1 0 62008 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1477_
timestamp 1607194113
transform 1 0 61180 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1073_
timestamp 1607194113
transform 1 0 61732 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1607194113
transform 1 0 61732 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_674
timestamp 1607194113
transform 1 0 63112 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_684
timestamp 1607194113
transform 1 0 64032 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_672
timestamp 1607194113
transform 1 0 62928 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_670
timestamp 1607194113
transform 1 0 62744 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_683
timestamp 1607194113
transform 1 0 63940 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_671
timestamp 1607194113
transform 1 0 62836 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__CLK
timestamp 1607194113
transform 1 0 62928 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1607194113
transform 1 0 62836 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_698
timestamp 1607194113
transform 1 0 65320 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_686
timestamp 1607194113
transform 1 0 64216 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_696
timestamp 1607194113
transform 1 0 65136 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_695
timestamp 1607194113
transform 1 0 65044 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_478
timestamp 1607194113
transform 1 0 45080 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_497
timestamp 1607194113
transform 1 0 46828 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_490
timestamp 1607194113
transform 1 0 46184 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1607194113
transform 1 0 46736 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_521
timestamp 1607194113
transform 1 0 49036 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_509
timestamp 1607194113
transform 1 0 47932 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_540
timestamp 1607194113
transform 1 0 50784 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_528
timestamp 1607194113
transform 1 0 49680 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1607194113
transform 1 0 49588 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_559
timestamp 1607194113
transform 1 0 52532 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_552
timestamp 1607194113
transform 1 0 51888 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1607194113
transform 1 0 52440 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_583
timestamp 1607194113
transform 1 0 54740 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_571
timestamp 1607194113
transform 1 0 53636 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_602
timestamp 1607194113
transform 1 0 56488 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_590
timestamp 1607194113
transform 1 0 55384 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1607194113
transform 1 0 55292 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_621
timestamp 1607194113
transform 1 0 58236 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_614
timestamp 1607194113
transform 1 0 57592 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1607194113
transform 1 0 58144 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_633
timestamp 1607194113
transform 1 0 59340 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_664
timestamp 1607194113
transform 1 0 62192 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_652
timestamp 1607194113
transform 1 0 61088 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_645
timestamp 1607194113
transform 1 0 60444 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1607194113
transform 1 0 60996 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_683
timestamp 1607194113
transform 1 0 63940 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_676
timestamp 1607194113
transform 1 0 63296 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1607194113
transform 1 0 63848 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_695
timestamp 1607194113
transform 1 0 65044 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_715
timestamp 1607194113
transform 1 0 66884 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_703
timestamp 1607194113
transform 1 0 65780 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_701
timestamp 1607194113
transform 1 0 65596 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1607194113
transform 1 0 65688 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_720
timestamp 1607194113
transform 1 0 67344 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_708
timestamp 1607194113
transform 1 0 66240 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_715
timestamp 1607194113
transform 1 0 66884 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_703
timestamp 1607194113
transform 1 0 65780 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1607194113
transform 1 0 65688 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_714
timestamp 1607194113
transform 1 0 66792 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_707
timestamp 1607194113
transform 1 0 66148 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1607194113
transform 1 0 66700 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_739
timestamp 1607194113
transform 1 0 69092 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_727
timestamp 1607194113
transform 1 0 67988 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_745
timestamp 1607194113
transform 1 0 69644 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_733
timestamp 1607194113
transform 1 0 68540 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1607194113
transform 1 0 68448 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_739
timestamp 1607194113
transform 1 0 69092 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_727
timestamp 1607194113
transform 1 0 67988 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_745
timestamp 1607194113
transform 1 0 69644 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_738
timestamp 1607194113
transform 1 0 69000 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_726
timestamp 1607194113
transform 1 0 67896 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1607194113
transform 1 0 69552 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_757
timestamp 1607194113
transform 1 0 70748 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_764
timestamp 1607194113
transform 1 0 71392 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_751
timestamp 1607194113
transform 1 0 70196 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_757
timestamp 1607194113
transform 1 0 70748 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_764
timestamp 1607194113
transform 1 0 71392 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_751
timestamp 1607194113
transform 1 0 70196 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1607194113
transform 1 0 71300 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1607194113
transform 1 0 71300 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_788
timestamp 1607194113
transform 1 0 73600 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_776
timestamp 1607194113
transform 1 0 72496 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_781
timestamp 1607194113
transform 1 0 72956 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_769
timestamp 1607194113
transform 1 0 71852 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_788
timestamp 1607194113
transform 1 0 73600 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_776
timestamp 1607194113
transform 1 0 72496 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_788
timestamp 1607194113
transform 1 0 73600 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_776
timestamp 1607194113
transform 1 0 72496 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_769
timestamp 1607194113
transform 1 0 71852 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1607194113
transform 1 0 72404 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_812
timestamp 1607194113
transform 1 0 75808 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_800
timestamp 1607194113
transform 1 0 74704 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_806
timestamp 1607194113
transform 1 0 75256 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_794
timestamp 1607194113
transform 1 0 74152 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1607194113
transform 1 0 74060 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_812
timestamp 1607194113
transform 1 0 75808 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_800
timestamp 1607194113
transform 1 0 74704 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_807
timestamp 1607194113
transform 1 0 75348 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_800
timestamp 1607194113
transform 1 0 74704 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1607194113
transform 1 0 75256 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_837
timestamp 1607194113
transform 1 0 78108 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_825
timestamp 1607194113
transform 1 0 77004 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1607194113
transform 1 0 76912 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_830
timestamp 1607194113
transform 1 0 77464 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_818
timestamp 1607194113
transform 1 0 76360 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_837
timestamp 1607194113
transform 1 0 78108 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_825
timestamp 1607194113
transform 1 0 77004 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1607194113
transform 1 0 76912 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_838
timestamp 1607194113
transform 1 0 78200 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_831
timestamp 1607194113
transform 1 0 77556 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_819
timestamp 1607194113
transform 1 0 76452 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1607194113
transform 1 0 78108 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_850
timestamp 1607194113
transform 1 0 79304 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_861
timestamp 1607194113
transform 1 0 80316 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_849
timestamp 1607194113
transform 1 0 79212 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_855
timestamp 1607194113
transform 1 0 79764 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_842
timestamp 1607194113
transform 1 0 78568 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_861
timestamp 1607194113
transform 1 0 80316 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_849
timestamp 1607194113
transform 1 0 79212 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1607194113
transform 1 0 79672 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_873
timestamp 1607194113
transform 1 0 81420 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1607194113
transform 1 0 82524 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_879
timestamp 1607194113
transform 1 0 81972 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_867
timestamp 1607194113
transform 1 0 80868 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_873
timestamp 1607194113
transform 1 0 81420 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1607194113
transform 1 0 82524 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_881
timestamp 1607194113
transform 1 0 82156 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_869
timestamp 1607194113
transform 1 0 81052 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_862
timestamp 1607194113
transform 1 0 80408 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1607194113
transform 1 0 80960 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_900
timestamp 1607194113
transform 1 0 83904 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_893
timestamp 1607194113
transform 1 0 83260 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_898
timestamp 1607194113
transform 1 0 83720 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_886
timestamp 1607194113
transform 1 0 82616 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_903
timestamp 1607194113
transform 1 0 84180 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_891
timestamp 1607194113
transform 1 0 83076 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_898
timestamp 1607194113
transform 1 0 83720 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_886
timestamp 1607194113
transform 1 0 82616 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1607194113
transform 1 0 83812 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_922
timestamp 1607194113
transform 1 0 85928 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_910
timestamp 1607194113
transform 1 0 84824 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_928
timestamp 1607194113
transform 1 0 86480 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_916
timestamp 1607194113
transform 1 0 85376 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1607194113
transform 1 0 85284 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_922
timestamp 1607194113
transform 1 0 85928 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_910
timestamp 1607194113
transform 1 0 84824 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_931
timestamp 1607194113
transform 1 0 86756 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_924
timestamp 1607194113
transform 1 0 86112 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_912
timestamp 1607194113
transform 1 0 85008 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1607194113
transform 1 0 86664 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_947
timestamp 1607194113
transform 1 0 88228 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_934
timestamp 1607194113
transform 1 0 87032 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1607194113
transform 1 0 88136 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_952
timestamp 1607194113
transform 1 0 88688 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_940
timestamp 1607194113
transform 1 0 87584 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_947
timestamp 1607194113
transform 1 0 88228 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_934
timestamp 1607194113
transform 1 0 87032 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1607194113
transform 1 0 88136 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_955
timestamp 1607194113
transform 1 0 88964 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_943
timestamp 1607194113
transform 1 0 87860 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_971
timestamp 1607194113
transform 1 0 90436 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_959
timestamp 1607194113
transform 1 0 89332 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_977
timestamp 1607194113
transform 1 0 90988 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_964
timestamp 1607194113
transform 1 0 89792 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1607194113
transform 1 0 90896 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_971
timestamp 1607194113
transform 1 0 90436 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_959
timestamp 1607194113
transform 1 0 89332 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_974
timestamp 1607194113
transform 1 0 90712 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_962
timestamp 1607194113
transform 1 0 89608 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1607194113
transform 1 0 89516 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_993
timestamp 1607194113
transform 1 0 92460 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_986
timestamp 1607194113
transform 1 0 91816 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_995
timestamp 1607194113
transform 1 0 92644 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_983
timestamp 1607194113
transform 1 0 91540 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1001
timestamp 1607194113
transform 1 0 93196 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_989
timestamp 1607194113
transform 1 0 92092 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_995
timestamp 1607194113
transform 1 0 92644 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_983
timestamp 1607194113
transform 1 0 91540 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1607194113
transform 1 0 92368 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1020
timestamp 1607194113
transform 1 0 94944 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1008
timestamp 1607194113
transform 1 0 93840 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1607194113
transform 1 0 93748 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1013
timestamp 1607194113
transform 1 0 94300 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1020
timestamp 1607194113
transform 1 0 94944 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1008
timestamp 1607194113
transform 1 0 93840 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1607194113
transform 1 0 93748 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1024
timestamp 1607194113
transform 1 0 95312 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_1017
timestamp 1607194113
transform 1 0 94668 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1005
timestamp 1607194113
transform 1 0 93564 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1607194113
transform 1 0 95220 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1036
timestamp 1607194113
transform 1 0 96416 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1044
timestamp 1607194113
transform 1 0 97152 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1032
timestamp 1607194113
transform 1 0 96048 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1038
timestamp 1607194113
transform 1 0 96600 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1025
timestamp 1607194113
transform 1 0 95404 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1044
timestamp 1607194113
transform 1 0 97152 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1032
timestamp 1607194113
transform 1 0 96048 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1607194113
transform 1 0 96508 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1069
timestamp 1607194113
transform 1 0 99452 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1056
timestamp 1607194113
transform 1 0 98256 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1607194113
transform 1 0 99360 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1062
timestamp 1607194113
transform 1 0 98808 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1050
timestamp 1607194113
transform 1 0 97704 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1069
timestamp 1607194113
transform 1 0 99452 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1056
timestamp 1607194113
transform 1 0 98256 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1607194113
transform 1 0 99360 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1067
timestamp 1607194113
transform 1 0 99268 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1055
timestamp 1607194113
transform 1 0 98164 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_1048
timestamp 1607194113
transform 1 0 97520 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1607194113
transform 1 0 98072 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1086
timestamp 1607194113
transform 1 0 101016 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_1079
timestamp 1607194113
transform 1 0 100372 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1093
timestamp 1607194113
transform 1 0 101660 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1081
timestamp 1607194113
transform 1 0 100556 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1086
timestamp 1607194113
transform 1 0 101016 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1074
timestamp 1607194113
transform 1 0 99912 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1093
timestamp 1607194113
transform 1 0 101660 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1081
timestamp 1607194113
transform 1 0 100556 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1607194113
transform 1 0 100924 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1117
timestamp 1607194113
transform 1 0 103868 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1105
timestamp 1607194113
transform 1 0 102764 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1111
timestamp 1607194113
transform 1 0 103316 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1099
timestamp 1607194113
transform 1 0 102212 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1607194113
transform 1 0 102120 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1117
timestamp 1607194113
transform 1 0 103868 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1105
timestamp 1607194113
transform 1 0 102764 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1117
timestamp 1607194113
transform 1 0 103868 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_1110
timestamp 1607194113
transform 1 0 103224 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1098
timestamp 1607194113
transform 1 0 102120 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1607194113
transform 1 0 103776 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_1129
timestamp 1607194113
transform 1 0 104972 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1130
timestamp 1607194113
transform 1 0 105064 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1135
timestamp 1607194113
transform 1 0 105524 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1123
timestamp 1607194113
transform 1 0 104420 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1130
timestamp 1607194113
transform 1 0 105064 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1607194113
transform 1 0 104972 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1607194113
transform 1 0 104972 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1158
timestamp 1607194113
transform 1 0 107640 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_1154
timestamp 1607194113
transform 1 0 107272 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_1142
timestamp 1607194113
transform 1 0 106168 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1607194113
transform -1 0 108008 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_1147
timestamp 1607194113
transform 1 0 106628 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1607194113
transform -1 0 108008 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1158
timestamp 1607194113
transform 1 0 107640 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_1154
timestamp 1607194113
transform 1 0 107272 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_1142
timestamp 1607194113
transform 1 0 106168 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1607194113
transform -1 0 108008 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_83_1156
timestamp 1607194113
transform 1 0 107456 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_1148
timestamp 1607194113
transform 1 0 106720 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_83_1141
timestamp 1607194113
transform 1 0 106076 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1607194113
transform 1 0 106628 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1607194113
transform -1 0 108008 0 1 47328
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 280 800 400 6 bus_in[0]
port 0 nsew default input
rlabel metal3 s 0 13200 800 13320 6 bus_in[10]
port 1 nsew default input
rlabel metal3 s 0 14560 800 14680 6 bus_in[11]
port 2 nsew default input
rlabel metal3 s 0 15784 800 15904 6 bus_in[12]
port 3 nsew default input
rlabel metal3 s 0 17144 800 17264 6 bus_in[13]
port 4 nsew default input
rlabel metal3 s 0 18368 800 18488 6 bus_in[14]
port 5 nsew default input
rlabel metal3 s 0 19728 800 19848 6 bus_in[15]
port 6 nsew default input
rlabel metal3 s 0 20952 800 21072 6 bus_in[16]
port 7 nsew default input
rlabel metal3 s 0 22312 800 22432 6 bus_in[17]
port 8 nsew default input
rlabel metal3 s 0 23672 800 23792 6 bus_in[18]
port 9 nsew default input
rlabel metal3 s 0 24896 800 25016 6 bus_in[19]
port 10 nsew default input
rlabel metal3 s 0 1504 800 1624 6 bus_in[1]
port 11 nsew default input
rlabel metal3 s 0 26256 800 26376 6 bus_in[20]
port 12 nsew default input
rlabel metal3 s 0 27480 800 27600 6 bus_in[21]
port 13 nsew default input
rlabel metal3 s 0 28840 800 28960 6 bus_in[22]
port 14 nsew default input
rlabel metal3 s 0 30064 800 30184 6 bus_in[23]
port 15 nsew default input
rlabel metal3 s 0 31424 800 31544 6 bus_in[24]
port 16 nsew default input
rlabel metal3 s 0 32648 800 32768 6 bus_in[25]
port 17 nsew default input
rlabel metal3 s 0 34008 800 34128 6 bus_in[26]
port 18 nsew default input
rlabel metal3 s 0 35368 800 35488 6 bus_in[27]
port 19 nsew default input
rlabel metal3 s 0 36592 800 36712 6 bus_in[28]
port 20 nsew default input
rlabel metal3 s 0 37952 800 38072 6 bus_in[29]
port 21 nsew default input
rlabel metal3 s 0 2864 800 2984 6 bus_in[2]
port 22 nsew default input
rlabel metal3 s 0 39176 800 39296 6 bus_in[30]
port 23 nsew default input
rlabel metal3 s 0 40536 800 40656 6 bus_in[31]
port 24 nsew default input
rlabel metal3 s 0 41760 800 41880 6 bus_in[32]
port 25 nsew default input
rlabel metal3 s 0 43120 800 43240 6 bus_in[33]
port 26 nsew default input
rlabel metal3 s 0 44344 800 44464 6 bus_in[34]
port 27 nsew default input
rlabel metal3 s 0 45704 800 45824 6 bus_in[35]
port 28 nsew default input
rlabel metal3 s 0 46384 800 46504 6 bus_in[36]
port 29 nsew default input
rlabel metal3 s 0 47064 800 47184 6 bus_in[37]
port 30 nsew default input
rlabel metal3 s 0 47608 800 47728 6 bus_in[38]
port 31 nsew default input
rlabel metal3 s 0 48288 800 48408 6 bus_in[39]
port 32 nsew default input
rlabel metal3 s 0 4088 800 4208 6 bus_in[3]
port 33 nsew default input
rlabel metal3 s 0 48968 800 49088 6 bus_in[40]
port 34 nsew default input
rlabel metal3 s 0 49648 800 49768 6 bus_in[41]
port 35 nsew default input
rlabel metal3 s 0 5448 800 5568 6 bus_in[4]
port 36 nsew default input
rlabel metal3 s 0 6672 800 6792 6 bus_in[5]
port 37 nsew default input
rlabel metal3 s 0 8032 800 8152 6 bus_in[6]
port 38 nsew default input
rlabel metal3 s 0 9256 800 9376 6 bus_in[7]
port 39 nsew default input
rlabel metal3 s 0 10616 800 10736 6 bus_in[8]
port 40 nsew default input
rlabel metal3 s 0 11976 800 12096 6 bus_in[9]
port 41 nsew default input
rlabel metal3 s 0 824 800 944 6 bus_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 13880 800 14000 6 bus_out[10]
port 43 nsew default tristate
rlabel metal3 s 0 15104 800 15224 6 bus_out[11]
port 44 nsew default tristate
rlabel metal3 s 0 16464 800 16584 6 bus_out[12]
port 45 nsew default tristate
rlabel metal3 s 0 17824 800 17944 6 bus_out[13]
port 46 nsew default tristate
rlabel metal3 s 0 19048 800 19168 6 bus_out[14]
port 47 nsew default tristate
rlabel metal3 s 0 20408 800 20528 6 bus_out[15]
port 48 nsew default tristate
rlabel metal3 s 0 21632 800 21752 6 bus_out[16]
port 49 nsew default tristate
rlabel metal3 s 0 22992 800 23112 6 bus_out[17]
port 50 nsew default tristate
rlabel metal3 s 0 24216 800 24336 6 bus_out[18]
port 51 nsew default tristate
rlabel metal3 s 0 25576 800 25696 6 bus_out[19]
port 52 nsew default tristate
rlabel metal3 s 0 2184 800 2304 6 bus_out[1]
port 53 nsew default tristate
rlabel metal3 s 0 26800 800 26920 6 bus_out[20]
port 54 nsew default tristate
rlabel metal3 s 0 28160 800 28280 6 bus_out[21]
port 55 nsew default tristate
rlabel metal3 s 0 29520 800 29640 6 bus_out[22]
port 56 nsew default tristate
rlabel metal3 s 0 30744 800 30864 6 bus_out[23]
port 57 nsew default tristate
rlabel metal3 s 0 32104 800 32224 6 bus_out[24]
port 58 nsew default tristate
rlabel metal3 s 0 33328 800 33448 6 bus_out[25]
port 59 nsew default tristate
rlabel metal3 s 0 34688 800 34808 6 bus_out[26]
port 60 nsew default tristate
rlabel metal3 s 0 35912 800 36032 6 bus_out[27]
port 61 nsew default tristate
rlabel metal3 s 0 37272 800 37392 6 bus_out[28]
port 62 nsew default tristate
rlabel metal3 s 0 38496 800 38616 6 bus_out[29]
port 63 nsew default tristate
rlabel metal3 s 0 3408 800 3528 6 bus_out[2]
port 64 nsew default tristate
rlabel metal3 s 0 39856 800 39976 6 bus_out[30]
port 65 nsew default tristate
rlabel metal3 s 0 41216 800 41336 6 bus_out[31]
port 66 nsew default tristate
rlabel metal3 s 0 42440 800 42560 6 bus_out[32]
port 67 nsew default tristate
rlabel metal3 s 0 43800 800 43920 6 bus_out[33]
port 68 nsew default tristate
rlabel metal3 s 0 45024 800 45144 6 bus_out[34]
port 69 nsew default tristate
rlabel metal3 s 0 4768 800 4888 6 bus_out[3]
port 70 nsew default tristate
rlabel metal3 s 0 6128 800 6248 6 bus_out[4]
port 71 nsew default tristate
rlabel metal3 s 0 7352 800 7472 6 bus_out[5]
port 72 nsew default tristate
rlabel metal3 s 0 8712 800 8832 6 bus_out[6]
port 73 nsew default tristate
rlabel metal3 s 0 9936 800 10056 6 bus_out[7]
port 74 nsew default tristate
rlabel metal3 s 0 11296 800 11416 6 bus_out[8]
port 75 nsew default tristate
rlabel metal3 s 0 12520 800 12640 6 bus_out[9]
port 76 nsew default tristate
rlabel metal2 s 54574 0 54630 800 6 clk_i
port 77 nsew default input
rlabel metal2 s 54482 49248 54538 50048 6 out1_o
port 78 nsew default tristate
rlabel metal2 s 90822 49248 90878 50048 6 out2_o
port 79 nsew default tristate
rlabel metal2 s 18142 49248 18198 50048 6 rst_n_i
port 80 nsew default input
rlabel metal5 s 1104 6436 108008 7036 6 VPWR
port 81 nsew default input
rlabel metal5 s 1104 24436 108008 25036 6 VGND
port 82 nsew default input
<< properties >>
string FIXED_BBOX 0 0 108256 50048
<< end >>
