VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO delayline_9_hd_25_1
  CLASS BLOCK ;
  FOREIGN delayline_9_hd_25_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 108.010 BY 115.925 ;
  PIN inp_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 4.000 4.600 4.600 ;
    END
  END inp_i
  PIN out_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 4.000 110.080 4.600 110.680 ;
    END
  END out_o
  PIN en_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 44.800 4.600 45.400 ;
    END
  END en_i[8]
  PIN en_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 66.560 4.600 67.160 ;
    END
  END en_i[7]
  PIN en_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 77.440 4.600 78.040 ;
    END
  END en_i[6]
  PIN en_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 82.880 4.600 83.480 ;
    END
  END en_i[5]
  PIN en_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 88.320 4.600 88.920 ;
    END
  END en_i[4]
  PIN en_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 93.760 4.600 94.360 ;
    END
  END en_i[3]
  PIN en_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 99.200 4.600 99.800 ;
    END
  END en_i[2]
  PIN en_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 104.640 4.600 105.240 ;
    END
  END en_i[1]
  PIN en_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 4.000 107.360 4.600 107.960 ;
    END
  END en_i[0]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 9.520 12.800 103.820 14.400 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 9.520 102.800 103.820 104.400 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 9.520 4.555 103.820 110.805 ;
      LAYER met1 ;
        RECT 9.395 4.400 103.820 110.960 ;
      LAYER met2 ;
        RECT 9.610 4.400 101.420 111.925 ;
      LAYER met3 ;
        RECT 4.150 111.080 90.240 111.905 ;
        RECT 5.000 109.680 90.240 111.080 ;
        RECT 4.150 108.360 90.240 109.680 ;
        RECT 5.000 106.960 90.240 108.360 ;
        RECT 4.150 105.640 90.240 106.960 ;
        RECT 5.000 104.240 90.240 105.640 ;
        RECT 4.150 100.200 90.240 104.240 ;
        RECT 5.000 98.800 90.240 100.200 ;
        RECT 4.150 94.760 90.240 98.800 ;
        RECT 5.000 93.360 90.240 94.760 ;
        RECT 4.150 89.320 90.240 93.360 ;
        RECT 5.000 87.920 90.240 89.320 ;
        RECT 4.150 83.880 90.240 87.920 ;
        RECT 5.000 82.480 90.240 83.880 ;
        RECT 4.150 78.440 90.240 82.480 ;
        RECT 5.000 77.040 90.240 78.440 ;
        RECT 4.150 67.560 90.240 77.040 ;
        RECT 5.000 66.160 90.240 67.560 ;
        RECT 4.150 45.800 90.240 66.160 ;
        RECT 5.000 44.400 90.240 45.800 ;
        RECT 4.150 5.000 90.240 44.400 ;
        RECT 5.000 4.475 90.240 5.000 ;
      LAYER met4 ;
        RECT 22.040 4.400 90.240 110.960 ;
  END
END delayline_9_hd_25_1
END LIBRARY

