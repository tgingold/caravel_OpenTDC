magic
tech sky130A
magscale 1 2
timestamp 1607274881
<< viali >>
rect 1933 22025 1967 22059
rect 2301 21957 2335 21991
rect 2393 21889 2427 21923
rect 3773 21889 3807 21923
rect 2485 21821 2519 21855
rect 3129 21821 3163 21855
rect 1933 21481 1967 21515
rect 2485 21345 2519 21379
rect 3129 21345 3163 21379
rect 2393 21209 2427 21243
rect 3773 21209 3807 21243
rect 2301 21141 2335 21175
rect 3773 20937 3807 20971
rect 3129 20733 3163 20767
rect 1933 20393 1967 20427
rect 2485 20257 2519 20291
rect 3129 20257 3163 20291
rect 4969 20257 5003 20291
rect 2393 20189 2427 20223
rect 3773 20189 3807 20223
rect 4325 20189 4359 20223
rect 2301 20053 2335 20087
rect 4969 19849 5003 19883
rect 3129 19645 3163 19679
rect 3773 19645 3807 19679
rect 4325 19645 4359 19679
rect 1933 19305 1967 19339
rect 2485 19169 2519 19203
rect 3129 19169 3163 19203
rect 4969 19169 5003 19203
rect 5521 19169 5555 19203
rect 7361 19169 7395 19203
rect 2393 19101 2427 19135
rect 3773 19101 3807 19135
rect 4325 19101 4359 19135
rect 6165 19101 6199 19135
rect 6717 19101 6751 19135
rect 2301 18965 2335 18999
rect 7361 18761 7395 18795
rect 3129 18557 3163 18591
rect 3773 18557 3807 18591
rect 4325 18557 4359 18591
rect 4969 18557 5003 18591
rect 5521 18557 5555 18591
rect 6165 18557 6199 18591
rect 6717 18557 6751 18591
rect 1933 18217 1967 18251
rect 10949 18149 10983 18183
rect 2485 18081 2519 18115
rect 3129 18081 3163 18115
rect 4969 18081 5003 18115
rect 5521 18081 5555 18115
rect 7361 18081 7395 18115
rect 7913 18081 7947 18115
rect 9109 18081 9143 18115
rect 10305 18081 10339 18115
rect 12145 18081 12179 18115
rect 2393 18013 2427 18047
rect 3773 18013 3807 18047
rect 4325 18013 4359 18047
rect 6165 18013 6199 18047
rect 6717 18013 6751 18047
rect 8557 18013 8591 18047
rect 9753 18013 9787 18047
rect 11501 18013 11535 18047
rect 2301 17877 2335 17911
rect 12145 17673 12179 17707
rect 3129 17537 3163 17571
rect 3773 17537 3807 17571
rect 4325 17537 4359 17571
rect 4969 17537 5003 17571
rect 5521 17537 5555 17571
rect 6165 17537 6199 17571
rect 6717 17537 6751 17571
rect 7361 17537 7395 17571
rect 7913 17537 7947 17571
rect 8557 17537 8591 17571
rect 9109 17537 9143 17571
rect 9753 17537 9787 17571
rect 10305 17537 10339 17571
rect 10949 17537 10983 17571
rect 11501 17537 11535 17571
rect 1933 17129 1967 17163
rect 2485 16993 2519 17027
rect 3129 16993 3163 17027
rect 4969 16993 5003 17027
rect 5521 16993 5555 17027
rect 7361 16993 7395 17027
rect 7913 16993 7947 17027
rect 9109 16993 9143 17027
rect 10949 16993 10983 17027
rect 11501 16993 11535 17027
rect 13341 16993 13375 17027
rect 13893 16993 13927 17027
rect 15733 16993 15767 17027
rect 16285 16993 16319 17027
rect 18125 16993 18159 17027
rect 18677 16993 18711 17027
rect 20517 16993 20551 17027
rect 4325 16925 4359 16959
rect 6165 16925 6199 16959
rect 6717 16925 6751 16959
rect 8557 16925 8591 16959
rect 9753 16925 9787 16959
rect 10305 16925 10339 16959
rect 12145 16925 12179 16959
rect 12697 16925 12731 16959
rect 14537 16925 14571 16959
rect 15089 16925 15123 16959
rect 16929 16925 16963 16959
rect 17481 16925 17515 16959
rect 19321 16925 19355 16959
rect 19873 16925 19907 16959
rect 21069 16925 21103 16959
rect 2393 16857 2427 16891
rect 3773 16857 3807 16891
rect 2301 16789 2335 16823
rect 21713 16789 21747 16823
rect 21713 16585 21747 16619
rect 3129 16381 3163 16415
rect 3773 16381 3807 16415
rect 4325 16381 4359 16415
rect 4969 16381 5003 16415
rect 5521 16381 5555 16415
rect 6165 16381 6199 16415
rect 6717 16381 6751 16415
rect 7361 16381 7395 16415
rect 7913 16381 7947 16415
rect 8557 16381 8591 16415
rect 9109 16381 9143 16415
rect 9753 16381 9787 16415
rect 10305 16381 10339 16415
rect 10949 16381 10983 16415
rect 11501 16381 11535 16415
rect 12145 16381 12179 16415
rect 12697 16381 12731 16415
rect 13341 16381 13375 16415
rect 13893 16381 13927 16415
rect 14537 16381 14571 16415
rect 15089 16381 15123 16415
rect 15733 16381 15767 16415
rect 16285 16381 16319 16415
rect 16929 16381 16963 16415
rect 17481 16381 17515 16415
rect 18125 16381 18159 16415
rect 18677 16381 18711 16415
rect 19321 16381 19355 16415
rect 19873 16381 19907 16415
rect 20517 16381 20551 16415
rect 21069 16381 21103 16415
rect 1933 15973 1967 16007
rect 2485 15905 2519 15939
rect 3129 15905 3163 15939
rect 4969 15905 5003 15939
rect 5521 15905 5555 15939
rect 7361 15905 7395 15939
rect 7913 15905 7947 15939
rect 9109 15905 9143 15939
rect 10949 15905 10983 15939
rect 11501 15905 11535 15939
rect 13341 15905 13375 15939
rect 13893 15905 13927 15939
rect 15733 15905 15767 15939
rect 16285 15905 16319 15939
rect 18125 15905 18159 15939
rect 18677 15905 18711 15939
rect 20517 15905 20551 15939
rect 2393 15837 2427 15871
rect 3773 15837 3807 15871
rect 4325 15837 4359 15871
rect 6165 15837 6199 15871
rect 6717 15837 6751 15871
rect 8557 15837 8591 15871
rect 9753 15837 9787 15871
rect 10305 15837 10339 15871
rect 12145 15837 12179 15871
rect 12697 15837 12731 15871
rect 14537 15837 14571 15871
rect 15089 15837 15123 15871
rect 16929 15837 16963 15871
rect 17481 15837 17515 15871
rect 19321 15837 19355 15871
rect 19873 15837 19907 15871
rect 21069 15837 21103 15871
rect 2301 15701 2335 15735
rect 21713 15701 21747 15735
rect 21713 15497 21747 15531
rect 3129 15361 3163 15395
rect 3773 15293 3807 15327
rect 4325 15293 4359 15327
rect 4969 15293 5003 15327
rect 5521 15293 5555 15327
rect 6165 15293 6199 15327
rect 6717 15293 6751 15327
rect 7361 15293 7395 15327
rect 7913 15293 7947 15327
rect 8557 15293 8591 15327
rect 9109 15293 9143 15327
rect 9753 15293 9787 15327
rect 10305 15293 10339 15327
rect 10949 15293 10983 15327
rect 11501 15293 11535 15327
rect 12145 15293 12179 15327
rect 12697 15293 12731 15327
rect 13341 15293 13375 15327
rect 13893 15293 13927 15327
rect 14537 15293 14571 15327
rect 15089 15293 15123 15327
rect 15733 15293 15767 15327
rect 16285 15293 16319 15327
rect 16929 15293 16963 15327
rect 17481 15293 17515 15327
rect 18125 15293 18159 15327
rect 18677 15293 18711 15327
rect 19321 15293 19355 15327
rect 19873 15293 19907 15327
rect 20517 15293 20551 15327
rect 21069 15293 21103 15327
rect 3773 14953 3807 14987
rect 3129 14817 3163 14851
rect 4969 14817 5003 14851
rect 5521 14817 5555 14851
rect 7361 14817 7395 14851
rect 7913 14817 7947 14851
rect 9109 14817 9143 14851
rect 10949 14817 10983 14851
rect 11501 14817 11535 14851
rect 13341 14817 13375 14851
rect 13893 14817 13927 14851
rect 15733 14817 15767 14851
rect 16285 14817 16319 14851
rect 18125 14817 18159 14851
rect 18677 14817 18711 14851
rect 20517 14817 20551 14851
rect 4325 14749 4359 14783
rect 6165 14749 6199 14783
rect 6717 14749 6751 14783
rect 8557 14749 8591 14783
rect 9753 14749 9787 14783
rect 10305 14749 10339 14783
rect 12145 14749 12179 14783
rect 12697 14749 12731 14783
rect 14537 14749 14571 14783
rect 15089 14749 15123 14783
rect 16929 14749 16963 14783
rect 17481 14749 17515 14783
rect 19321 14749 19355 14783
rect 19873 14749 19907 14783
rect 21069 14749 21103 14783
rect 21713 14613 21747 14647
rect 21713 14409 21747 14443
rect 3129 14273 3163 14307
rect 3773 14205 3807 14239
rect 4325 14205 4359 14239
rect 4969 14205 5003 14239
rect 5521 14205 5555 14239
rect 6165 14205 6199 14239
rect 6717 14205 6751 14239
rect 7361 14205 7395 14239
rect 7913 14205 7947 14239
rect 8557 14205 8591 14239
rect 9109 14205 9143 14239
rect 9753 14205 9787 14239
rect 10305 14205 10339 14239
rect 10949 14205 10983 14239
rect 11501 14205 11535 14239
rect 12145 14205 12179 14239
rect 12697 14205 12731 14239
rect 13341 14205 13375 14239
rect 13893 14205 13927 14239
rect 14537 14205 14571 14239
rect 15089 14205 15123 14239
rect 15733 14205 15767 14239
rect 16285 14205 16319 14239
rect 16929 14205 16963 14239
rect 17481 14205 17515 14239
rect 18125 14205 18159 14239
rect 18677 14205 18711 14239
rect 19321 14205 19355 14239
rect 19873 14205 19907 14239
rect 20517 14205 20551 14239
rect 21069 14205 21103 14239
rect 1933 13797 1967 13831
rect 2485 13729 2519 13763
rect 3129 13729 3163 13763
rect 4969 13729 5003 13763
rect 5521 13729 5555 13763
rect 7361 13729 7395 13763
rect 7913 13729 7947 13763
rect 9109 13729 9143 13763
rect 10949 13729 10983 13763
rect 11501 13729 11535 13763
rect 13341 13729 13375 13763
rect 13893 13729 13927 13763
rect 15733 13729 15767 13763
rect 16285 13729 16319 13763
rect 18125 13729 18159 13763
rect 18677 13729 18711 13763
rect 20517 13729 20551 13763
rect 4325 13661 4359 13695
rect 6165 13661 6199 13695
rect 6717 13661 6751 13695
rect 8557 13661 8591 13695
rect 9753 13661 9787 13695
rect 10305 13661 10339 13695
rect 12145 13661 12179 13695
rect 12697 13661 12731 13695
rect 14537 13661 14571 13695
rect 15089 13661 15123 13695
rect 16929 13661 16963 13695
rect 17481 13661 17515 13695
rect 19321 13661 19355 13695
rect 19873 13661 19907 13695
rect 21069 13661 21103 13695
rect 2393 13593 2427 13627
rect 3773 13593 3807 13627
rect 2301 13525 2335 13559
rect 21713 13525 21747 13559
rect 21713 13321 21747 13355
rect 3129 13185 3163 13219
rect 3773 13117 3807 13151
rect 4325 13117 4359 13151
rect 4969 13117 5003 13151
rect 5521 13117 5555 13151
rect 6165 13117 6199 13151
rect 6717 13117 6751 13151
rect 7361 13117 7395 13151
rect 7913 13117 7947 13151
rect 8557 13117 8591 13151
rect 9109 13117 9143 13151
rect 9753 13117 9787 13151
rect 10305 13117 10339 13151
rect 10949 13117 10983 13151
rect 11501 13117 11535 13151
rect 12145 13117 12179 13151
rect 12697 13117 12731 13151
rect 13341 13117 13375 13151
rect 13893 13117 13927 13151
rect 14537 13117 14571 13151
rect 15089 13117 15123 13151
rect 15733 13117 15767 13151
rect 16285 13117 16319 13151
rect 16929 13117 16963 13151
rect 17481 13117 17515 13151
rect 18125 13117 18159 13151
rect 18677 13117 18711 13151
rect 19321 13117 19355 13151
rect 19873 13117 19907 13151
rect 20517 13117 20551 13151
rect 21069 13117 21103 13151
rect 3773 12777 3807 12811
rect 3129 12641 3163 12675
rect 4969 12641 5003 12675
rect 5521 12641 5555 12675
rect 7361 12641 7395 12675
rect 7913 12641 7947 12675
rect 9109 12641 9143 12675
rect 10949 12641 10983 12675
rect 11501 12641 11535 12675
rect 13341 12641 13375 12675
rect 13893 12641 13927 12675
rect 15733 12641 15767 12675
rect 16285 12641 16319 12675
rect 18125 12641 18159 12675
rect 18677 12641 18711 12675
rect 20517 12641 20551 12675
rect 4325 12573 4359 12607
rect 6165 12573 6199 12607
rect 6717 12573 6751 12607
rect 8557 12573 8591 12607
rect 9753 12573 9787 12607
rect 10305 12573 10339 12607
rect 12145 12573 12179 12607
rect 12697 12573 12731 12607
rect 14537 12573 14571 12607
rect 15089 12573 15123 12607
rect 16929 12573 16963 12607
rect 17481 12573 17515 12607
rect 19321 12573 19355 12607
rect 19873 12573 19907 12607
rect 21069 12573 21103 12607
rect 21713 12437 21747 12471
rect 21713 12233 21747 12267
rect 3129 12097 3163 12131
rect 3773 12029 3807 12063
rect 4325 12029 4359 12063
rect 4969 12029 5003 12063
rect 5521 12029 5555 12063
rect 6165 12029 6199 12063
rect 6717 12029 6751 12063
rect 7361 12029 7395 12063
rect 7913 12029 7947 12063
rect 8557 12029 8591 12063
rect 9109 12029 9143 12063
rect 9753 12029 9787 12063
rect 10305 12029 10339 12063
rect 10949 12029 10983 12063
rect 11501 12029 11535 12063
rect 12145 12029 12179 12063
rect 12697 12029 12731 12063
rect 13341 12029 13375 12063
rect 13893 12029 13927 12063
rect 14537 12029 14571 12063
rect 15089 12029 15123 12063
rect 15733 12029 15767 12063
rect 16285 12029 16319 12063
rect 16929 12029 16963 12063
rect 17481 12029 17515 12063
rect 18125 12029 18159 12063
rect 18677 12029 18711 12063
rect 19321 12029 19355 12063
rect 19873 12029 19907 12063
rect 20517 12029 20551 12063
rect 21069 12029 21103 12063
rect 3773 11553 3807 11587
rect 5521 11553 5555 11587
rect 7361 11553 7395 11587
rect 8557 11553 8591 11587
rect 9109 11553 9143 11587
rect 10949 11553 10983 11587
rect 11501 11553 11535 11587
rect 13341 11553 13375 11587
rect 13893 11553 13927 11587
rect 15733 11553 15767 11587
rect 16285 11553 16319 11587
rect 18125 11553 18159 11587
rect 18677 11553 18711 11587
rect 20517 11553 20551 11587
rect 3129 11485 3163 11519
rect 4325 11485 4359 11519
rect 6165 11485 6199 11519
rect 6717 11485 6751 11519
rect 7913 11485 7947 11519
rect 9753 11485 9787 11519
rect 10305 11485 10339 11519
rect 12145 11485 12179 11519
rect 12697 11485 12731 11519
rect 14537 11485 14571 11519
rect 15089 11485 15123 11519
rect 16929 11485 16963 11519
rect 17481 11485 17515 11519
rect 19321 11485 19355 11519
rect 19873 11485 19907 11519
rect 21069 11485 21103 11519
rect 4969 11417 5003 11451
rect 21713 11349 21747 11383
rect 21713 11145 21747 11179
rect 3129 11009 3163 11043
rect 3773 10941 3807 10975
rect 4325 10941 4359 10975
rect 4969 10941 5003 10975
rect 5521 10941 5555 10975
rect 6165 10941 6199 10975
rect 6717 10941 6751 10975
rect 7361 10941 7395 10975
rect 7913 10941 7947 10975
rect 8557 10941 8591 10975
rect 9109 10941 9143 10975
rect 9753 10941 9787 10975
rect 10305 10941 10339 10975
rect 10949 10941 10983 10975
rect 11501 10941 11535 10975
rect 12145 10941 12179 10975
rect 12697 10941 12731 10975
rect 13341 10941 13375 10975
rect 13893 10941 13927 10975
rect 14537 10941 14571 10975
rect 15089 10941 15123 10975
rect 15733 10941 15767 10975
rect 16285 10941 16319 10975
rect 16929 10941 16963 10975
rect 17481 10941 17515 10975
rect 18125 10941 18159 10975
rect 18677 10941 18711 10975
rect 19321 10941 19355 10975
rect 19873 10941 19907 10975
rect 20517 10941 20551 10975
rect 21069 10941 21103 10975
rect 3773 10601 3807 10635
rect 3129 10465 3163 10499
rect 4969 10465 5003 10499
rect 5521 10465 5555 10499
rect 7361 10465 7395 10499
rect 8557 10465 8591 10499
rect 9109 10465 9143 10499
rect 10949 10465 10983 10499
rect 11501 10465 11535 10499
rect 13341 10465 13375 10499
rect 13893 10465 13927 10499
rect 15733 10465 15767 10499
rect 16285 10465 16319 10499
rect 18125 10465 18159 10499
rect 18677 10465 18711 10499
rect 20517 10465 20551 10499
rect 4325 10397 4359 10431
rect 6165 10397 6199 10431
rect 6717 10397 6751 10431
rect 7913 10397 7947 10431
rect 9753 10397 9787 10431
rect 10305 10397 10339 10431
rect 12145 10397 12179 10431
rect 12697 10397 12731 10431
rect 14537 10397 14571 10431
rect 15089 10397 15123 10431
rect 16929 10397 16963 10431
rect 17481 10397 17515 10431
rect 19321 10397 19355 10431
rect 19873 10397 19907 10431
rect 21069 10397 21103 10431
rect 21713 10261 21747 10295
rect 21713 10057 21747 10091
rect 3129 9921 3163 9955
rect 3773 9853 3807 9887
rect 4325 9853 4359 9887
rect 4969 9853 5003 9887
rect 5521 9853 5555 9887
rect 6165 9853 6199 9887
rect 6717 9853 6751 9887
rect 7361 9853 7395 9887
rect 7913 9853 7947 9887
rect 8557 9853 8591 9887
rect 9109 9853 9143 9887
rect 9753 9853 9787 9887
rect 10305 9853 10339 9887
rect 10949 9853 10983 9887
rect 11501 9853 11535 9887
rect 12145 9853 12179 9887
rect 12697 9853 12731 9887
rect 13341 9853 13375 9887
rect 13893 9853 13927 9887
rect 14537 9853 14571 9887
rect 15089 9853 15123 9887
rect 15733 9853 15767 9887
rect 16285 9853 16319 9887
rect 16929 9853 16963 9887
rect 17481 9853 17515 9887
rect 18125 9853 18159 9887
rect 18677 9853 18711 9887
rect 19321 9853 19355 9887
rect 19873 9853 19907 9887
rect 20517 9853 20551 9887
rect 21069 9853 21103 9887
rect 2485 9377 2519 9411
rect 3129 9377 3163 9411
rect 4969 9377 5003 9411
rect 5521 9377 5555 9411
rect 7361 9377 7395 9411
rect 8557 9377 8591 9411
rect 9109 9377 9143 9411
rect 10949 9377 10983 9411
rect 11501 9377 11535 9411
rect 13341 9377 13375 9411
rect 13893 9377 13927 9411
rect 15733 9377 15767 9411
rect 16285 9377 16319 9411
rect 18125 9377 18159 9411
rect 18677 9377 18711 9411
rect 20517 9377 20551 9411
rect 4325 9309 4359 9343
rect 6165 9309 6199 9343
rect 6717 9309 6751 9343
rect 7913 9309 7947 9343
rect 9753 9309 9787 9343
rect 10305 9309 10339 9343
rect 12145 9309 12179 9343
rect 12697 9309 12731 9343
rect 14537 9309 14571 9343
rect 15089 9309 15123 9343
rect 16929 9309 16963 9343
rect 17481 9309 17515 9343
rect 19321 9309 19355 9343
rect 19873 9309 19907 9343
rect 21069 9309 21103 9343
rect 2393 9241 2427 9275
rect 3773 9241 3807 9275
rect 1933 9173 1967 9207
rect 2301 9173 2335 9207
rect 21713 9173 21747 9207
rect 21713 8969 21747 9003
rect 3129 8833 3163 8867
rect 3773 8765 3807 8799
rect 4325 8765 4359 8799
rect 4969 8765 5003 8799
rect 5521 8765 5555 8799
rect 6165 8765 6199 8799
rect 6717 8765 6751 8799
rect 7361 8765 7395 8799
rect 7913 8765 7947 8799
rect 8557 8765 8591 8799
rect 9109 8765 9143 8799
rect 9753 8765 9787 8799
rect 10305 8765 10339 8799
rect 10949 8765 10983 8799
rect 11501 8765 11535 8799
rect 12145 8765 12179 8799
rect 12697 8765 12731 8799
rect 13341 8765 13375 8799
rect 13893 8765 13927 8799
rect 14537 8765 14571 8799
rect 15089 8765 15123 8799
rect 15733 8765 15767 8799
rect 16285 8765 16319 8799
rect 16929 8765 16963 8799
rect 17481 8765 17515 8799
rect 18125 8765 18159 8799
rect 18677 8765 18711 8799
rect 19321 8765 19355 8799
rect 19873 8765 19907 8799
rect 20517 8765 20551 8799
rect 21069 8765 21103 8799
rect 3773 8425 3807 8459
rect 3129 8289 3163 8323
rect 4969 8289 5003 8323
rect 5521 8289 5555 8323
rect 7361 8289 7395 8323
rect 8557 8289 8591 8323
rect 9109 8289 9143 8323
rect 10949 8289 10983 8323
rect 11501 8289 11535 8323
rect 13341 8289 13375 8323
rect 13893 8289 13927 8323
rect 15733 8289 15767 8323
rect 16285 8289 16319 8323
rect 18125 8289 18159 8323
rect 18677 8289 18711 8323
rect 20517 8289 20551 8323
rect 4325 8221 4359 8255
rect 6165 8221 6199 8255
rect 6717 8221 6751 8255
rect 7913 8221 7947 8255
rect 9753 8221 9787 8255
rect 10305 8221 10339 8255
rect 12145 8221 12179 8255
rect 12697 8221 12731 8255
rect 14537 8221 14571 8255
rect 15089 8221 15123 8255
rect 16929 8221 16963 8255
rect 17481 8221 17515 8255
rect 19321 8221 19355 8255
rect 19873 8221 19907 8255
rect 21069 8221 21103 8255
rect 21713 8085 21747 8119
rect 21713 7881 21747 7915
rect 3129 7745 3163 7779
rect 3773 7677 3807 7711
rect 4325 7677 4359 7711
rect 4969 7677 5003 7711
rect 5521 7677 5555 7711
rect 6165 7677 6199 7711
rect 6717 7677 6751 7711
rect 7361 7677 7395 7711
rect 7913 7677 7947 7711
rect 8557 7677 8591 7711
rect 9109 7677 9143 7711
rect 9753 7677 9787 7711
rect 10305 7677 10339 7711
rect 10949 7677 10983 7711
rect 11501 7677 11535 7711
rect 12145 7677 12179 7711
rect 12697 7677 12731 7711
rect 13341 7677 13375 7711
rect 13893 7677 13927 7711
rect 14537 7677 14571 7711
rect 15089 7677 15123 7711
rect 15733 7677 15767 7711
rect 16285 7677 16319 7711
rect 16929 7677 16963 7711
rect 17481 7677 17515 7711
rect 18125 7677 18159 7711
rect 18677 7677 18711 7711
rect 19321 7677 19355 7711
rect 19873 7677 19907 7711
rect 20517 7677 20551 7711
rect 21069 7677 21103 7711
rect 11501 7201 11535 7235
rect 13893 7201 13927 7235
rect 3129 7133 3163 7167
rect 3773 7133 3807 7167
rect 4325 7133 4359 7167
rect 5521 7133 5555 7167
rect 6717 7133 6751 7167
rect 7913 7133 7947 7167
rect 9109 7133 9143 7167
rect 10305 7133 10339 7167
rect 12145 7133 12179 7167
rect 12697 7133 12731 7167
rect 14537 7133 14571 7167
rect 15089 7133 15123 7167
rect 16285 7133 16319 7167
rect 17481 7133 17515 7167
rect 18677 7133 18711 7167
rect 19873 7133 19907 7167
rect 21069 7133 21103 7167
rect 4969 7065 5003 7099
rect 7361 7065 7395 7099
rect 8557 7065 8591 7099
rect 9753 7065 9787 7099
rect 15733 7065 15767 7099
rect 18125 7065 18159 7099
rect 20517 7065 20551 7099
rect 6165 6997 6199 7031
rect 10949 6997 10983 7031
rect 13341 6997 13375 7031
rect 16929 6997 16963 7031
rect 19321 6997 19355 7031
rect 21713 6997 21747 7031
rect 21713 6793 21747 6827
rect 3129 6657 3163 6691
rect 3773 6589 3807 6623
rect 4325 6589 4359 6623
rect 4969 6589 5003 6623
rect 5521 6589 5555 6623
rect 6165 6589 6199 6623
rect 6717 6589 6751 6623
rect 7361 6589 7395 6623
rect 7913 6589 7947 6623
rect 8557 6589 8591 6623
rect 9109 6589 9143 6623
rect 9753 6589 9787 6623
rect 10305 6589 10339 6623
rect 10949 6589 10983 6623
rect 11501 6589 11535 6623
rect 12145 6589 12179 6623
rect 12697 6589 12731 6623
rect 13341 6589 13375 6623
rect 13893 6589 13927 6623
rect 14537 6589 14571 6623
rect 15089 6589 15123 6623
rect 15733 6589 15767 6623
rect 16285 6589 16319 6623
rect 16929 6589 16963 6623
rect 17481 6589 17515 6623
rect 18125 6589 18159 6623
rect 18677 6589 18711 6623
rect 19321 6589 19355 6623
rect 19873 6589 19907 6623
rect 20517 6589 20551 6623
rect 21069 6589 21103 6623
rect 3773 6249 3807 6283
rect 3129 6113 3163 6147
rect 4969 6113 5003 6147
rect 5521 6113 5555 6147
rect 7361 6113 7395 6147
rect 7913 6113 7947 6147
rect 9109 6113 9143 6147
rect 10949 6113 10983 6147
rect 11501 6113 11535 6147
rect 13341 6113 13375 6147
rect 13893 6113 13927 6147
rect 15733 6113 15767 6147
rect 16285 6113 16319 6147
rect 18125 6113 18159 6147
rect 19321 6113 19355 6147
rect 19873 6113 19907 6147
rect 21713 6113 21747 6147
rect 4325 6045 4359 6079
rect 6165 6045 6199 6079
rect 6717 6045 6751 6079
rect 8557 6045 8591 6079
rect 9753 6045 9787 6079
rect 10305 6045 10339 6079
rect 12145 6045 12179 6079
rect 12697 6045 12731 6079
rect 14537 6045 14571 6079
rect 15089 6045 15123 6079
rect 16929 6045 16963 6079
rect 17481 6045 17515 6079
rect 18677 6045 18711 6079
rect 20517 6045 20551 6079
rect 21069 6045 21103 6079
rect 21713 5705 21747 5739
rect 3129 5569 3163 5603
rect 3773 5501 3807 5535
rect 4325 5501 4359 5535
rect 4969 5501 5003 5535
rect 5521 5501 5555 5535
rect 6165 5501 6199 5535
rect 6717 5501 6751 5535
rect 7361 5501 7395 5535
rect 7913 5501 7947 5535
rect 8557 5501 8591 5535
rect 9109 5501 9143 5535
rect 9753 5501 9787 5535
rect 10305 5501 10339 5535
rect 10949 5501 10983 5535
rect 11501 5501 11535 5535
rect 12145 5501 12179 5535
rect 12697 5501 12731 5535
rect 13341 5501 13375 5535
rect 13893 5501 13927 5535
rect 14537 5501 14571 5535
rect 15089 5501 15123 5535
rect 15733 5501 15767 5535
rect 16285 5501 16319 5535
rect 16929 5501 16963 5535
rect 17481 5501 17515 5535
rect 18125 5501 18159 5535
rect 18677 5501 18711 5535
rect 19321 5501 19355 5535
rect 19873 5501 19907 5535
rect 20517 5501 20551 5535
rect 21069 5501 21103 5535
rect 12145 5161 12179 5195
rect 6165 5093 6199 5127
rect 9753 5093 9787 5127
rect 13341 5093 13375 5127
rect 15733 5093 15767 5127
rect 19321 5093 19355 5127
rect 3129 5025 3163 5059
rect 4325 5025 4359 5059
rect 5521 5025 5555 5059
rect 6717 5025 6751 5059
rect 7913 5025 7947 5059
rect 9109 5025 9143 5059
rect 10305 5025 10339 5059
rect 11501 5025 11535 5059
rect 12697 5025 12731 5059
rect 13893 5025 13927 5059
rect 15089 5025 15123 5059
rect 16285 5025 16319 5059
rect 18677 5025 18711 5059
rect 19873 5025 19907 5059
rect 21713 5025 21747 5059
rect 3773 4957 3807 4991
rect 4969 4957 5003 4991
rect 7361 4957 7395 4991
rect 8557 4957 8591 4991
rect 14537 4957 14571 4991
rect 16929 4957 16963 4991
rect 17481 4957 17515 4991
rect 18125 4957 18159 4991
rect 20517 4957 20551 4991
rect 21069 4957 21103 4991
rect 10949 4889 10983 4923
rect 21713 4617 21747 4651
rect 3129 4481 3163 4515
rect 3773 4413 3807 4447
rect 4325 4413 4359 4447
rect 4969 4413 5003 4447
rect 5521 4413 5555 4447
rect 6165 4413 6199 4447
rect 6717 4413 6751 4447
rect 7361 4413 7395 4447
rect 7913 4413 7947 4447
rect 8557 4413 8591 4447
rect 9109 4413 9143 4447
rect 9753 4413 9787 4447
rect 10305 4413 10339 4447
rect 10949 4413 10983 4447
rect 11501 4413 11535 4447
rect 12145 4413 12179 4447
rect 12697 4413 12731 4447
rect 13341 4413 13375 4447
rect 13893 4413 13927 4447
rect 14537 4413 14571 4447
rect 15089 4413 15123 4447
rect 15733 4413 15767 4447
rect 16285 4413 16319 4447
rect 16929 4413 16963 4447
rect 17481 4413 17515 4447
rect 18125 4413 18159 4447
rect 18677 4413 18711 4447
rect 19321 4413 19355 4447
rect 19873 4413 19907 4447
rect 20517 4413 20551 4447
rect 21069 4413 21103 4447
rect 3773 4073 3807 4107
rect 3129 3937 3163 3971
rect 4969 3937 5003 3971
rect 5521 3937 5555 3971
rect 7361 3937 7395 3971
rect 7913 3937 7947 3971
rect 9109 3937 9143 3971
rect 10949 3937 10983 3971
rect 11501 3937 11535 3971
rect 13341 3937 13375 3971
rect 13893 3937 13927 3971
rect 15733 3937 15767 3971
rect 16285 3937 16319 3971
rect 18125 3937 18159 3971
rect 19321 3937 19355 3971
rect 19873 3937 19907 3971
rect 21713 3937 21747 3971
rect 4325 3869 4359 3903
rect 6165 3869 6199 3903
rect 6717 3869 6751 3903
rect 8557 3869 8591 3903
rect 9753 3869 9787 3903
rect 10305 3869 10339 3903
rect 12145 3869 12179 3903
rect 12697 3869 12731 3903
rect 14537 3869 14571 3903
rect 15089 3869 15123 3903
rect 16929 3869 16963 3903
rect 17481 3869 17515 3903
rect 18677 3869 18711 3903
rect 20517 3869 20551 3903
rect 21069 3869 21103 3903
rect 21713 3461 21747 3495
rect 3129 3393 3163 3427
rect 3773 3325 3807 3359
rect 4325 3325 4359 3359
rect 4969 3325 5003 3359
rect 5521 3325 5555 3359
rect 6165 3325 6199 3359
rect 6717 3325 6751 3359
rect 7361 3325 7395 3359
rect 7913 3325 7947 3359
rect 8557 3325 8591 3359
rect 9109 3325 9143 3359
rect 9753 3325 9787 3359
rect 10305 3325 10339 3359
rect 10949 3325 10983 3359
rect 11501 3325 11535 3359
rect 12145 3325 12179 3359
rect 12697 3325 12731 3359
rect 13341 3325 13375 3359
rect 13893 3325 13927 3359
rect 14537 3325 14571 3359
rect 15089 3325 15123 3359
rect 15733 3325 15767 3359
rect 16285 3325 16319 3359
rect 16929 3325 16963 3359
rect 17481 3325 17515 3359
rect 18125 3325 18159 3359
rect 18677 3325 18711 3359
rect 19321 3325 19355 3359
rect 19873 3325 19907 3359
rect 20517 3325 20551 3359
rect 21069 3325 21103 3359
rect 3773 2985 3807 3019
rect 4325 2849 4359 2883
rect 6165 2849 6199 2883
rect 7913 2849 7947 2883
rect 9753 2849 9787 2883
rect 11501 2849 11535 2883
rect 13341 2849 13375 2883
rect 13893 2849 13927 2883
rect 15733 2849 15767 2883
rect 16285 2849 16319 2883
rect 17481 2849 17515 2883
rect 19321 2849 19355 2883
rect 19873 2849 19907 2883
rect 21713 2849 21747 2883
rect 3129 2781 3163 2815
rect 5521 2781 5555 2815
rect 6717 2781 6751 2815
rect 9109 2781 9143 2815
rect 10305 2781 10339 2815
rect 12145 2781 12179 2815
rect 12697 2781 12731 2815
rect 15089 2781 15123 2815
rect 18677 2781 18711 2815
rect 21069 2781 21103 2815
rect 4969 2713 5003 2747
rect 7361 2713 7395 2747
rect 8557 2713 8591 2747
rect 14537 2713 14571 2747
rect 16929 2713 16963 2747
rect 18125 2713 18159 2747
rect 20517 2713 20551 2747
rect 10949 2645 10983 2679
rect 21713 2441 21747 2475
rect 3129 2305 3163 2339
rect 3773 2237 3807 2271
rect 4325 2237 4359 2271
rect 4969 2237 5003 2271
rect 5521 2237 5555 2271
rect 6165 2237 6199 2271
rect 6717 2237 6751 2271
rect 7361 2237 7395 2271
rect 7913 2237 7947 2271
rect 8557 2237 8591 2271
rect 9109 2237 9143 2271
rect 9753 2237 9787 2271
rect 10305 2237 10339 2271
rect 10949 2237 10983 2271
rect 11501 2237 11535 2271
rect 12145 2237 12179 2271
rect 12697 2237 12731 2271
rect 13341 2237 13375 2271
rect 13893 2237 13927 2271
rect 14537 2237 14571 2271
rect 15089 2237 15123 2271
rect 15733 2237 15767 2271
rect 16285 2237 16319 2271
rect 16929 2237 16963 2271
rect 17481 2237 17515 2271
rect 18125 2237 18159 2271
rect 18677 2237 18711 2271
rect 19321 2237 19355 2271
rect 19873 2237 19907 2271
rect 20517 2237 20551 2271
rect 21069 2237 21103 2271
rect 3773 1897 3807 1931
rect 3129 1761 3163 1795
rect 4969 1761 5003 1795
rect 5521 1761 5555 1795
rect 7361 1761 7395 1795
rect 7913 1761 7947 1795
rect 9109 1761 9143 1795
rect 10949 1761 10983 1795
rect 11501 1761 11535 1795
rect 13341 1761 13375 1795
rect 13893 1761 13927 1795
rect 15733 1761 15767 1795
rect 16285 1761 16319 1795
rect 18125 1761 18159 1795
rect 19321 1761 19355 1795
rect 19873 1761 19907 1795
rect 21713 1761 21747 1795
rect 4325 1693 4359 1727
rect 6165 1693 6199 1727
rect 6717 1693 6751 1727
rect 8557 1693 8591 1727
rect 9753 1693 9787 1727
rect 10305 1693 10339 1727
rect 12145 1693 12179 1727
rect 12697 1693 12731 1727
rect 14537 1693 14571 1727
rect 15089 1693 15123 1727
rect 16929 1693 16963 1727
rect 17481 1693 17515 1727
rect 18677 1693 18711 1727
rect 20517 1693 20551 1727
rect 21069 1693 21103 1727
rect 21713 1285 21747 1319
rect 3129 1149 3163 1183
rect 3773 1149 3807 1183
rect 4325 1149 4359 1183
rect 4969 1149 5003 1183
rect 5521 1149 5555 1183
rect 6165 1149 6199 1183
rect 6717 1149 6751 1183
rect 7361 1149 7395 1183
rect 7913 1149 7947 1183
rect 8557 1149 8591 1183
rect 9109 1149 9143 1183
rect 9753 1149 9787 1183
rect 10305 1149 10339 1183
rect 10949 1149 10983 1183
rect 11501 1149 11535 1183
rect 12145 1149 12179 1183
rect 12697 1149 12731 1183
rect 13341 1149 13375 1183
rect 13893 1149 13927 1183
rect 14537 1149 14571 1183
rect 15089 1149 15123 1183
rect 15733 1149 15767 1183
rect 16285 1149 16319 1183
rect 16929 1149 16963 1183
rect 17481 1149 17515 1183
rect 18125 1149 18159 1183
rect 18677 1149 18711 1183
rect 19321 1149 19355 1183
rect 19873 1149 19907 1183
rect 20517 1149 20551 1183
rect 21069 1149 21103 1183
<< metal1 >>
rect 1904 22170 22236 22192
rect 1904 22118 4446 22170
rect 4498 22118 4510 22170
rect 4562 22118 4574 22170
rect 4626 22118 4638 22170
rect 4690 22118 9774 22170
rect 9826 22118 9838 22170
rect 9890 22118 9902 22170
rect 9954 22118 9966 22170
rect 10018 22118 15102 22170
rect 15154 22118 15166 22170
rect 15218 22118 15230 22170
rect 15282 22118 15294 22170
rect 15346 22118 20430 22170
rect 20482 22118 20494 22170
rect 20546 22118 20558 22170
rect 20610 22118 20622 22170
rect 20674 22118 22236 22170
rect 1904 22096 22236 22118
rect 1918 22056 1924 22068
rect 1879 22028 1924 22056
rect 1918 22016 1924 22028
rect 1976 22016 1982 22068
rect 2286 21988 2292 22000
rect 2247 21960 2292 21988
rect 2286 21948 2292 21960
rect 2344 21948 2350 22000
rect 2381 21923 2439 21929
rect 2381 21889 2393 21923
rect 2427 21920 2439 21923
rect 3761 21923 3819 21929
rect 3761 21920 3773 21923
rect 2427 21892 3773 21920
rect 2427 21889 2439 21892
rect 2381 21883 2439 21889
rect 3761 21889 3773 21892
rect 3807 21889 3819 21923
rect 3761 21883 3819 21889
rect 2470 21852 2476 21864
rect 2431 21824 2476 21852
rect 2470 21812 2476 21824
rect 2528 21812 2534 21864
rect 3117 21855 3175 21861
rect 3117 21821 3129 21855
rect 3163 21821 3175 21855
rect 3117 21815 3175 21821
rect 2286 21744 2292 21796
rect 2344 21784 2350 21796
rect 3132 21784 3160 21815
rect 2344 21756 3160 21784
rect 2344 21744 2350 21756
rect 1904 21626 22236 21648
rect 1904 21574 7110 21626
rect 7162 21574 7174 21626
rect 7226 21574 7238 21626
rect 7290 21574 7302 21626
rect 7354 21574 12438 21626
rect 12490 21574 12502 21626
rect 12554 21574 12566 21626
rect 12618 21574 12630 21626
rect 12682 21574 17766 21626
rect 17818 21574 17830 21626
rect 17882 21574 17894 21626
rect 17946 21574 17958 21626
rect 18010 21574 22236 21626
rect 1904 21552 22236 21574
rect 1921 21515 1979 21521
rect 1921 21481 1933 21515
rect 1967 21512 1979 21515
rect 2286 21512 2292 21524
rect 1967 21484 2292 21512
rect 1967 21481 1979 21484
rect 1921 21475 1979 21481
rect 2286 21472 2292 21484
rect 2344 21472 2350 21524
rect 2470 21376 2476 21388
rect 2431 21348 2476 21376
rect 2470 21336 2476 21348
rect 2528 21336 2534 21388
rect 3117 21379 3175 21385
rect 3117 21345 3129 21379
rect 3163 21376 3175 21379
rect 3758 21376 3764 21388
rect 3163 21348 3764 21376
rect 3163 21345 3175 21348
rect 3117 21339 3175 21345
rect 3758 21336 3764 21348
rect 3816 21336 3822 21388
rect 2381 21243 2439 21249
rect 2381 21209 2393 21243
rect 2427 21240 2439 21243
rect 3761 21243 3819 21249
rect 3761 21240 3773 21243
rect 2427 21212 3773 21240
rect 2427 21209 2439 21212
rect 2381 21203 2439 21209
rect 3761 21209 3773 21212
rect 3807 21209 3819 21243
rect 3761 21203 3819 21209
rect 2286 21132 2292 21184
rect 2344 21172 2350 21184
rect 2344 21144 2389 21172
rect 2344 21132 2350 21144
rect 1904 21082 22236 21104
rect 1904 21030 4446 21082
rect 4498 21030 4510 21082
rect 4562 21030 4574 21082
rect 4626 21030 4638 21082
rect 4690 21030 9774 21082
rect 9826 21030 9838 21082
rect 9890 21030 9902 21082
rect 9954 21030 9966 21082
rect 10018 21030 15102 21082
rect 15154 21030 15166 21082
rect 15218 21030 15230 21082
rect 15282 21030 15294 21082
rect 15346 21030 20430 21082
rect 20482 21030 20494 21082
rect 20546 21030 20558 21082
rect 20610 21030 20622 21082
rect 20674 21030 22236 21082
rect 1904 21008 22236 21030
rect 3758 20968 3764 20980
rect 3719 20940 3764 20968
rect 3758 20928 3764 20940
rect 3816 20928 3822 20980
rect 2286 20724 2292 20776
rect 2344 20764 2350 20776
rect 3117 20767 3175 20773
rect 3117 20764 3129 20767
rect 2344 20736 3129 20764
rect 2344 20724 2350 20736
rect 3117 20733 3129 20736
rect 3163 20733 3175 20767
rect 3117 20727 3175 20733
rect 1904 20538 22236 20560
rect 1904 20486 7110 20538
rect 7162 20486 7174 20538
rect 7226 20486 7238 20538
rect 7290 20486 7302 20538
rect 7354 20486 12438 20538
rect 12490 20486 12502 20538
rect 12554 20486 12566 20538
rect 12618 20486 12630 20538
rect 12682 20486 17766 20538
rect 17818 20486 17830 20538
rect 17882 20486 17894 20538
rect 17946 20486 17958 20538
rect 18010 20486 22236 20538
rect 1904 20464 22236 20486
rect 1921 20427 1979 20433
rect 1921 20393 1933 20427
rect 1967 20424 1979 20427
rect 2286 20424 2292 20436
rect 1967 20396 2292 20424
rect 1967 20393 1979 20396
rect 1921 20387 1979 20393
rect 2286 20384 2292 20396
rect 2344 20384 2350 20436
rect 2470 20288 2476 20300
rect 2431 20260 2476 20288
rect 2470 20248 2476 20260
rect 2528 20248 2534 20300
rect 3117 20291 3175 20297
rect 3117 20257 3129 20291
rect 3163 20288 3175 20291
rect 4957 20291 5015 20297
rect 4957 20288 4969 20291
rect 3163 20260 4969 20288
rect 3163 20257 3175 20260
rect 3117 20251 3175 20257
rect 4957 20257 4969 20260
rect 5003 20257 5015 20291
rect 4957 20251 5015 20257
rect 2381 20223 2439 20229
rect 2381 20189 2393 20223
rect 2427 20220 2439 20223
rect 3761 20223 3819 20229
rect 3761 20220 3773 20223
rect 2427 20192 3773 20220
rect 2427 20189 2439 20192
rect 2381 20183 2439 20189
rect 3761 20189 3773 20192
rect 3807 20189 3819 20223
rect 4310 20220 4316 20232
rect 4271 20192 4316 20220
rect 3761 20183 3819 20189
rect 4310 20180 4316 20192
rect 4368 20180 4374 20232
rect 2286 20044 2292 20096
rect 2344 20084 2350 20096
rect 2344 20056 2389 20084
rect 2344 20044 2350 20056
rect 1904 19994 22236 20016
rect 1904 19942 4446 19994
rect 4498 19942 4510 19994
rect 4562 19942 4574 19994
rect 4626 19942 4638 19994
rect 4690 19942 9774 19994
rect 9826 19942 9838 19994
rect 9890 19942 9902 19994
rect 9954 19942 9966 19994
rect 10018 19942 15102 19994
rect 15154 19942 15166 19994
rect 15218 19942 15230 19994
rect 15282 19942 15294 19994
rect 15346 19942 20430 19994
rect 20482 19942 20494 19994
rect 20546 19942 20558 19994
rect 20610 19942 20622 19994
rect 20674 19942 22236 19994
rect 1904 19920 22236 19942
rect 4310 19840 4316 19892
rect 4368 19880 4374 19892
rect 4957 19883 5015 19889
rect 4957 19880 4969 19883
rect 4368 19852 4969 19880
rect 4368 19840 4374 19852
rect 4957 19849 4969 19852
rect 5003 19849 5015 19883
rect 4957 19843 5015 19849
rect 2286 19636 2292 19688
rect 2344 19676 2350 19688
rect 3117 19679 3175 19685
rect 3117 19676 3129 19679
rect 2344 19648 3129 19676
rect 2344 19636 2350 19648
rect 3117 19645 3129 19648
rect 3163 19645 3175 19679
rect 3117 19639 3175 19645
rect 3761 19679 3819 19685
rect 3761 19645 3773 19679
rect 3807 19676 3819 19679
rect 4313 19679 4371 19685
rect 4313 19676 4325 19679
rect 3807 19648 4325 19676
rect 3807 19645 3819 19648
rect 3761 19639 3819 19645
rect 4313 19645 4325 19648
rect 4359 19645 4371 19679
rect 4313 19639 4371 19645
rect 1904 19450 22236 19472
rect 1904 19398 7110 19450
rect 7162 19398 7174 19450
rect 7226 19398 7238 19450
rect 7290 19398 7302 19450
rect 7354 19398 12438 19450
rect 12490 19398 12502 19450
rect 12554 19398 12566 19450
rect 12618 19398 12630 19450
rect 12682 19398 17766 19450
rect 17818 19398 17830 19450
rect 17882 19398 17894 19450
rect 17946 19398 17958 19450
rect 18010 19398 22236 19450
rect 1904 19376 22236 19398
rect 1921 19339 1979 19345
rect 1921 19305 1933 19339
rect 1967 19336 1979 19339
rect 2286 19336 2292 19348
rect 1967 19308 2292 19336
rect 1967 19305 1979 19308
rect 1921 19299 1979 19305
rect 2286 19296 2292 19308
rect 2344 19296 2350 19348
rect 2470 19200 2476 19212
rect 2431 19172 2476 19200
rect 2470 19160 2476 19172
rect 2528 19160 2534 19212
rect 3117 19203 3175 19209
rect 3117 19169 3129 19203
rect 3163 19200 3175 19203
rect 4957 19203 5015 19209
rect 4957 19200 4969 19203
rect 3163 19172 4969 19200
rect 3163 19169 3175 19172
rect 3117 19163 3175 19169
rect 4957 19169 4969 19172
rect 5003 19169 5015 19203
rect 4957 19163 5015 19169
rect 5509 19203 5567 19209
rect 5509 19169 5521 19203
rect 5555 19200 5567 19203
rect 7349 19203 7407 19209
rect 7349 19200 7361 19203
rect 5555 19172 7361 19200
rect 5555 19169 5567 19172
rect 5509 19163 5567 19169
rect 7349 19169 7361 19172
rect 7395 19169 7407 19203
rect 7349 19163 7407 19169
rect 2381 19135 2439 19141
rect 2381 19101 2393 19135
rect 2427 19132 2439 19135
rect 3761 19135 3819 19141
rect 3761 19132 3773 19135
rect 2427 19104 3773 19132
rect 2427 19101 2439 19104
rect 2381 19095 2439 19101
rect 3761 19101 3773 19104
rect 3807 19101 3819 19135
rect 3761 19095 3819 19101
rect 4313 19135 4371 19141
rect 4313 19101 4325 19135
rect 4359 19132 4371 19135
rect 6153 19135 6211 19141
rect 6153 19132 6165 19135
rect 4359 19104 6165 19132
rect 4359 19101 4371 19104
rect 4313 19095 4371 19101
rect 6153 19101 6165 19104
rect 6199 19101 6211 19135
rect 6702 19132 6708 19144
rect 6663 19104 6708 19132
rect 6153 19095 6211 19101
rect 6702 19092 6708 19104
rect 6760 19092 6766 19144
rect 2286 18956 2292 19008
rect 2344 18996 2350 19008
rect 2344 18968 2389 18996
rect 2344 18956 2350 18968
rect 1904 18906 22236 18928
rect 1904 18854 4446 18906
rect 4498 18854 4510 18906
rect 4562 18854 4574 18906
rect 4626 18854 4638 18906
rect 4690 18854 9774 18906
rect 9826 18854 9838 18906
rect 9890 18854 9902 18906
rect 9954 18854 9966 18906
rect 10018 18854 15102 18906
rect 15154 18854 15166 18906
rect 15218 18854 15230 18906
rect 15282 18854 15294 18906
rect 15346 18854 20430 18906
rect 20482 18854 20494 18906
rect 20546 18854 20558 18906
rect 20610 18854 20622 18906
rect 20674 18854 22236 18906
rect 1904 18832 22236 18854
rect 6702 18752 6708 18804
rect 6760 18792 6766 18804
rect 7349 18795 7407 18801
rect 7349 18792 7361 18795
rect 6760 18764 7361 18792
rect 6760 18752 6766 18764
rect 7349 18761 7361 18764
rect 7395 18761 7407 18795
rect 7349 18755 7407 18761
rect 2286 18548 2292 18600
rect 2344 18588 2350 18600
rect 3117 18591 3175 18597
rect 3117 18588 3129 18591
rect 2344 18560 3129 18588
rect 2344 18548 2350 18560
rect 3117 18557 3129 18560
rect 3163 18557 3175 18591
rect 3117 18551 3175 18557
rect 3761 18591 3819 18597
rect 3761 18557 3773 18591
rect 3807 18588 3819 18591
rect 4313 18591 4371 18597
rect 4313 18588 4325 18591
rect 3807 18560 4325 18588
rect 3807 18557 3819 18560
rect 3761 18551 3819 18557
rect 4313 18557 4325 18560
rect 4359 18557 4371 18591
rect 4313 18551 4371 18557
rect 4957 18591 5015 18597
rect 4957 18557 4969 18591
rect 5003 18588 5015 18591
rect 5509 18591 5567 18597
rect 5509 18588 5521 18591
rect 5003 18560 5521 18588
rect 5003 18557 5015 18560
rect 4957 18551 5015 18557
rect 5509 18557 5521 18560
rect 5555 18557 5567 18591
rect 5509 18551 5567 18557
rect 6153 18591 6211 18597
rect 6153 18557 6165 18591
rect 6199 18588 6211 18591
rect 6705 18591 6763 18597
rect 6705 18588 6717 18591
rect 6199 18560 6717 18588
rect 6199 18557 6211 18560
rect 6153 18551 6211 18557
rect 6705 18557 6717 18560
rect 6751 18557 6763 18591
rect 6705 18551 6763 18557
rect 1904 18362 22236 18384
rect 1904 18310 7110 18362
rect 7162 18310 7174 18362
rect 7226 18310 7238 18362
rect 7290 18310 7302 18362
rect 7354 18310 12438 18362
rect 12490 18310 12502 18362
rect 12554 18310 12566 18362
rect 12618 18310 12630 18362
rect 12682 18310 17766 18362
rect 17818 18310 17830 18362
rect 17882 18310 17894 18362
rect 17946 18310 17958 18362
rect 18010 18310 22236 18362
rect 1904 18288 22236 18310
rect 1921 18251 1979 18257
rect 1921 18217 1933 18251
rect 1967 18248 1979 18251
rect 2286 18248 2292 18260
rect 1967 18220 2292 18248
rect 1967 18217 1979 18220
rect 1921 18211 1979 18217
rect 2286 18208 2292 18220
rect 2344 18208 2350 18260
rect 10937 18183 10995 18189
rect 10937 18180 10949 18183
rect 10216 18152 10949 18180
rect 2470 18112 2476 18124
rect 2431 18084 2476 18112
rect 2470 18072 2476 18084
rect 2528 18072 2534 18124
rect 3117 18115 3175 18121
rect 3117 18081 3129 18115
rect 3163 18112 3175 18115
rect 4957 18115 5015 18121
rect 4957 18112 4969 18115
rect 3163 18084 4969 18112
rect 3163 18081 3175 18084
rect 3117 18075 3175 18081
rect 4957 18081 4969 18084
rect 5003 18081 5015 18115
rect 4957 18075 5015 18081
rect 5509 18115 5567 18121
rect 5509 18081 5521 18115
rect 5555 18112 5567 18115
rect 7349 18115 7407 18121
rect 7349 18112 7361 18115
rect 5555 18084 7361 18112
rect 5555 18081 5567 18084
rect 5509 18075 5567 18081
rect 7349 18081 7361 18084
rect 7395 18081 7407 18115
rect 7349 18075 7407 18081
rect 7901 18115 7959 18121
rect 7901 18081 7913 18115
rect 7947 18112 7959 18115
rect 9097 18115 9155 18121
rect 7947 18084 8772 18112
rect 7947 18081 7959 18084
rect 7901 18075 7959 18081
rect 2381 18047 2439 18053
rect 2381 18013 2393 18047
rect 2427 18044 2439 18047
rect 3761 18047 3819 18053
rect 3761 18044 3773 18047
rect 2427 18016 3773 18044
rect 2427 18013 2439 18016
rect 2381 18007 2439 18013
rect 3761 18013 3773 18016
rect 3807 18013 3819 18047
rect 3761 18007 3819 18013
rect 4313 18047 4371 18053
rect 4313 18013 4325 18047
rect 4359 18044 4371 18047
rect 6153 18047 6211 18053
rect 6153 18044 6165 18047
rect 4359 18016 6165 18044
rect 4359 18013 4371 18016
rect 4313 18007 4371 18013
rect 6153 18013 6165 18016
rect 6199 18013 6211 18047
rect 6153 18007 6211 18013
rect 6705 18047 6763 18053
rect 6705 18013 6717 18047
rect 6751 18044 6763 18047
rect 8545 18047 8603 18053
rect 8545 18044 8557 18047
rect 6751 18016 8557 18044
rect 6751 18013 6763 18016
rect 6705 18007 6763 18013
rect 8545 18013 8557 18016
rect 8591 18013 8603 18047
rect 8744 18044 8772 18084
rect 9097 18081 9109 18115
rect 9143 18112 9155 18115
rect 10216 18112 10244 18152
rect 10937 18149 10949 18152
rect 10983 18149 10995 18183
rect 10937 18143 10995 18149
rect 9143 18084 10244 18112
rect 10293 18115 10351 18121
rect 9143 18081 9155 18084
rect 9097 18075 9155 18081
rect 10293 18081 10305 18115
rect 10339 18112 10351 18115
rect 12133 18115 12191 18121
rect 12133 18112 12145 18115
rect 10339 18084 12145 18112
rect 10339 18081 10351 18084
rect 10293 18075 10351 18081
rect 12133 18081 12145 18084
rect 12179 18081 12191 18115
rect 12133 18075 12191 18081
rect 9741 18047 9799 18053
rect 9741 18044 9753 18047
rect 8744 18016 9753 18044
rect 8545 18007 8603 18013
rect 9741 18013 9753 18016
rect 9787 18013 9799 18047
rect 11486 18044 11492 18056
rect 11447 18016 11492 18044
rect 9741 18007 9799 18013
rect 11486 18004 11492 18016
rect 11544 18004 11550 18056
rect 2286 17868 2292 17920
rect 2344 17908 2350 17920
rect 2344 17880 2389 17908
rect 2344 17868 2350 17880
rect 1904 17818 22236 17840
rect 1904 17766 4446 17818
rect 4498 17766 4510 17818
rect 4562 17766 4574 17818
rect 4626 17766 4638 17818
rect 4690 17766 9774 17818
rect 9826 17766 9838 17818
rect 9890 17766 9902 17818
rect 9954 17766 9966 17818
rect 10018 17766 15102 17818
rect 15154 17766 15166 17818
rect 15218 17766 15230 17818
rect 15282 17766 15294 17818
rect 15346 17766 20430 17818
rect 20482 17766 20494 17818
rect 20546 17766 20558 17818
rect 20610 17766 20622 17818
rect 20674 17766 22236 17818
rect 1904 17744 22236 17766
rect 11486 17664 11492 17716
rect 11544 17704 11550 17716
rect 12133 17707 12191 17713
rect 12133 17704 12145 17707
rect 11544 17676 12145 17704
rect 11544 17664 11550 17676
rect 12133 17673 12145 17676
rect 12179 17673 12191 17707
rect 12133 17667 12191 17673
rect 2286 17528 2292 17580
rect 2344 17568 2350 17580
rect 3117 17571 3175 17577
rect 3117 17568 3129 17571
rect 2344 17540 3129 17568
rect 2344 17528 2350 17540
rect 3117 17537 3129 17540
rect 3163 17537 3175 17571
rect 3117 17531 3175 17537
rect 3761 17571 3819 17577
rect 3761 17537 3773 17571
rect 3807 17568 3819 17571
rect 4313 17571 4371 17577
rect 4313 17568 4325 17571
rect 3807 17540 4325 17568
rect 3807 17537 3819 17540
rect 3761 17531 3819 17537
rect 4313 17537 4325 17540
rect 4359 17537 4371 17571
rect 4313 17531 4371 17537
rect 4957 17571 5015 17577
rect 4957 17537 4969 17571
rect 5003 17568 5015 17571
rect 5509 17571 5567 17577
rect 5509 17568 5521 17571
rect 5003 17540 5521 17568
rect 5003 17537 5015 17540
rect 4957 17531 5015 17537
rect 5509 17537 5521 17540
rect 5555 17537 5567 17571
rect 5509 17531 5567 17537
rect 6153 17571 6211 17577
rect 6153 17537 6165 17571
rect 6199 17568 6211 17571
rect 6705 17571 6763 17577
rect 6705 17568 6717 17571
rect 6199 17540 6717 17568
rect 6199 17537 6211 17540
rect 6153 17531 6211 17537
rect 6705 17537 6717 17540
rect 6751 17537 6763 17571
rect 6705 17531 6763 17537
rect 7349 17571 7407 17577
rect 7349 17537 7361 17571
rect 7395 17568 7407 17571
rect 7901 17571 7959 17577
rect 7901 17568 7913 17571
rect 7395 17540 7913 17568
rect 7395 17537 7407 17540
rect 7349 17531 7407 17537
rect 7901 17537 7913 17540
rect 7947 17537 7959 17571
rect 7901 17531 7959 17537
rect 8545 17571 8603 17577
rect 8545 17537 8557 17571
rect 8591 17568 8603 17571
rect 9097 17571 9155 17577
rect 9097 17568 9109 17571
rect 8591 17540 9109 17568
rect 8591 17537 8603 17540
rect 8545 17531 8603 17537
rect 9097 17537 9109 17540
rect 9143 17537 9155 17571
rect 9097 17531 9155 17537
rect 9741 17571 9799 17577
rect 9741 17537 9753 17571
rect 9787 17568 9799 17571
rect 10293 17571 10351 17577
rect 10293 17568 10305 17571
rect 9787 17540 10305 17568
rect 9787 17537 9799 17540
rect 9741 17531 9799 17537
rect 10293 17537 10305 17540
rect 10339 17537 10351 17571
rect 10293 17531 10351 17537
rect 10937 17571 10995 17577
rect 10937 17537 10949 17571
rect 10983 17568 10995 17571
rect 11489 17571 11547 17577
rect 11489 17568 11501 17571
rect 10983 17540 11501 17568
rect 10983 17537 10995 17540
rect 10937 17531 10995 17537
rect 11489 17537 11501 17540
rect 11535 17537 11547 17571
rect 11489 17531 11547 17537
rect 1904 17274 22236 17296
rect 1904 17222 7110 17274
rect 7162 17222 7174 17274
rect 7226 17222 7238 17274
rect 7290 17222 7302 17274
rect 7354 17222 12438 17274
rect 12490 17222 12502 17274
rect 12554 17222 12566 17274
rect 12618 17222 12630 17274
rect 12682 17222 17766 17274
rect 17818 17222 17830 17274
rect 17882 17222 17894 17274
rect 17946 17222 17958 17274
rect 18010 17222 22236 17274
rect 1904 17200 22236 17222
rect 1921 17163 1979 17169
rect 1921 17129 1933 17163
rect 1967 17160 1979 17163
rect 2286 17160 2292 17172
rect 1967 17132 2292 17160
rect 1967 17129 1979 17132
rect 1921 17123 1979 17129
rect 2286 17120 2292 17132
rect 2344 17120 2350 17172
rect 2470 17024 2476 17036
rect 2431 16996 2476 17024
rect 2470 16984 2476 16996
rect 2528 16984 2534 17036
rect 3117 17027 3175 17033
rect 3117 16993 3129 17027
rect 3163 17024 3175 17027
rect 4957 17027 5015 17033
rect 4957 17024 4969 17027
rect 3163 16996 4969 17024
rect 3163 16993 3175 16996
rect 3117 16987 3175 16993
rect 4957 16993 4969 16996
rect 5003 16993 5015 17027
rect 4957 16987 5015 16993
rect 5509 17027 5567 17033
rect 5509 16993 5521 17027
rect 5555 17024 5567 17027
rect 7349 17027 7407 17033
rect 7349 17024 7361 17027
rect 5555 16996 7361 17024
rect 5555 16993 5567 16996
rect 5509 16987 5567 16993
rect 7349 16993 7361 16996
rect 7395 16993 7407 17027
rect 7349 16987 7407 16993
rect 7901 17027 7959 17033
rect 7901 16993 7913 17027
rect 7947 17024 7959 17027
rect 9097 17027 9155 17033
rect 7947 16996 8772 17024
rect 7947 16993 7959 16996
rect 7901 16987 7959 16993
rect 4313 16959 4371 16965
rect 4313 16925 4325 16959
rect 4359 16956 4371 16959
rect 6153 16959 6211 16965
rect 6153 16956 6165 16959
rect 4359 16928 6165 16956
rect 4359 16925 4371 16928
rect 4313 16919 4371 16925
rect 6153 16925 6165 16928
rect 6199 16925 6211 16959
rect 6153 16919 6211 16925
rect 6705 16959 6763 16965
rect 6705 16925 6717 16959
rect 6751 16956 6763 16959
rect 8545 16959 8603 16965
rect 8545 16956 8557 16959
rect 6751 16928 8557 16956
rect 6751 16925 6763 16928
rect 6705 16919 6763 16925
rect 8545 16925 8557 16928
rect 8591 16925 8603 16959
rect 8744 16956 8772 16996
rect 9097 16993 9109 17027
rect 9143 17024 9155 17027
rect 10937 17027 10995 17033
rect 10937 17024 10949 17027
rect 9143 16996 10949 17024
rect 9143 16993 9155 16996
rect 9097 16987 9155 16993
rect 10937 16993 10949 16996
rect 10983 16993 10995 17027
rect 10937 16987 10995 16993
rect 11489 17027 11547 17033
rect 11489 16993 11501 17027
rect 11535 17024 11547 17027
rect 13329 17027 13387 17033
rect 13329 17024 13341 17027
rect 11535 16996 13341 17024
rect 11535 16993 11547 16996
rect 11489 16987 11547 16993
rect 13329 16993 13341 16996
rect 13375 16993 13387 17027
rect 13329 16987 13387 16993
rect 13881 17027 13939 17033
rect 13881 16993 13893 17027
rect 13927 17024 13939 17027
rect 15721 17027 15779 17033
rect 15721 17024 15733 17027
rect 13927 16996 15733 17024
rect 13927 16993 13939 16996
rect 13881 16987 13939 16993
rect 15721 16993 15733 16996
rect 15767 16993 15779 17027
rect 15721 16987 15779 16993
rect 16273 17027 16331 17033
rect 16273 16993 16285 17027
rect 16319 17024 16331 17027
rect 18113 17027 18171 17033
rect 18113 17024 18125 17027
rect 16319 16996 18125 17024
rect 16319 16993 16331 16996
rect 16273 16987 16331 16993
rect 18113 16993 18125 16996
rect 18159 16993 18171 17027
rect 18113 16987 18171 16993
rect 18665 17027 18723 17033
rect 18665 16993 18677 17027
rect 18711 17024 18723 17027
rect 20505 17027 20563 17033
rect 20505 17024 20517 17027
rect 18711 16996 20517 17024
rect 18711 16993 18723 16996
rect 18665 16987 18723 16993
rect 20505 16993 20517 16996
rect 20551 16993 20563 17027
rect 20505 16987 20563 16993
rect 9741 16959 9799 16965
rect 9741 16956 9753 16959
rect 8744 16928 9753 16956
rect 8545 16919 8603 16925
rect 9741 16925 9753 16928
rect 9787 16925 9799 16959
rect 9741 16919 9799 16925
rect 10293 16959 10351 16965
rect 10293 16925 10305 16959
rect 10339 16956 10351 16959
rect 12133 16959 12191 16965
rect 12133 16956 12145 16959
rect 10339 16928 12145 16956
rect 10339 16925 10351 16928
rect 10293 16919 10351 16925
rect 12133 16925 12145 16928
rect 12179 16925 12191 16959
rect 12133 16919 12191 16925
rect 12685 16959 12743 16965
rect 12685 16925 12697 16959
rect 12731 16956 12743 16959
rect 14525 16959 14583 16965
rect 14525 16956 14537 16959
rect 12731 16928 14537 16956
rect 12731 16925 12743 16928
rect 12685 16919 12743 16925
rect 14525 16925 14537 16928
rect 14571 16925 14583 16959
rect 14525 16919 14583 16925
rect 15077 16959 15135 16965
rect 15077 16925 15089 16959
rect 15123 16956 15135 16959
rect 16917 16959 16975 16965
rect 16917 16956 16929 16959
rect 15123 16928 16929 16956
rect 15123 16925 15135 16928
rect 15077 16919 15135 16925
rect 16917 16925 16929 16928
rect 16963 16925 16975 16959
rect 16917 16919 16975 16925
rect 17469 16959 17527 16965
rect 17469 16925 17481 16959
rect 17515 16956 17527 16959
rect 19309 16959 19367 16965
rect 19309 16956 19321 16959
rect 17515 16928 19321 16956
rect 17515 16925 17527 16928
rect 17469 16919 17527 16925
rect 19309 16925 19321 16928
rect 19355 16925 19367 16959
rect 19309 16919 19367 16925
rect 19861 16959 19919 16965
rect 19861 16925 19873 16959
rect 19907 16925 19919 16959
rect 19861 16919 19919 16925
rect 21057 16959 21115 16965
rect 21057 16925 21069 16959
rect 21103 16956 21115 16959
rect 21606 16956 21612 16968
rect 21103 16928 21612 16956
rect 21103 16925 21115 16928
rect 21057 16919 21115 16925
rect 2381 16891 2439 16897
rect 2381 16857 2393 16891
rect 2427 16888 2439 16891
rect 3761 16891 3819 16897
rect 3761 16888 3773 16891
rect 2427 16860 3773 16888
rect 2427 16857 2439 16860
rect 2381 16851 2439 16857
rect 3761 16857 3773 16860
rect 3807 16857 3819 16891
rect 3761 16851 3819 16857
rect 2286 16780 2292 16832
rect 2344 16820 2350 16832
rect 19876 16820 19904 16919
rect 21606 16916 21612 16928
rect 21664 16916 21670 16968
rect 21701 16823 21759 16829
rect 21701 16820 21713 16823
rect 2344 16792 2389 16820
rect 19876 16792 21713 16820
rect 2344 16780 2350 16792
rect 21701 16789 21713 16792
rect 21747 16789 21759 16823
rect 21701 16783 21759 16789
rect 1904 16730 22236 16752
rect 1904 16678 4446 16730
rect 4498 16678 4510 16730
rect 4562 16678 4574 16730
rect 4626 16678 4638 16730
rect 4690 16678 9774 16730
rect 9826 16678 9838 16730
rect 9890 16678 9902 16730
rect 9954 16678 9966 16730
rect 10018 16678 15102 16730
rect 15154 16678 15166 16730
rect 15218 16678 15230 16730
rect 15282 16678 15294 16730
rect 15346 16678 20430 16730
rect 20482 16678 20494 16730
rect 20546 16678 20558 16730
rect 20610 16678 20622 16730
rect 20674 16678 22236 16730
rect 1904 16656 22236 16678
rect 21606 16576 21612 16628
rect 21664 16616 21670 16628
rect 21701 16619 21759 16625
rect 21701 16616 21713 16619
rect 21664 16588 21713 16616
rect 21664 16576 21670 16588
rect 21701 16585 21713 16588
rect 21747 16585 21759 16619
rect 21701 16579 21759 16585
rect 2378 16372 2384 16424
rect 2436 16412 2442 16424
rect 3117 16415 3175 16421
rect 3117 16412 3129 16415
rect 2436 16384 3129 16412
rect 2436 16372 2442 16384
rect 3117 16381 3129 16384
rect 3163 16381 3175 16415
rect 3117 16375 3175 16381
rect 3761 16415 3819 16421
rect 3761 16381 3773 16415
rect 3807 16412 3819 16415
rect 4313 16415 4371 16421
rect 4313 16412 4325 16415
rect 3807 16384 4325 16412
rect 3807 16381 3819 16384
rect 3761 16375 3819 16381
rect 4313 16381 4325 16384
rect 4359 16381 4371 16415
rect 4313 16375 4371 16381
rect 4957 16415 5015 16421
rect 4957 16381 4969 16415
rect 5003 16412 5015 16415
rect 5509 16415 5567 16421
rect 5509 16412 5521 16415
rect 5003 16384 5521 16412
rect 5003 16381 5015 16384
rect 4957 16375 5015 16381
rect 5509 16381 5521 16384
rect 5555 16381 5567 16415
rect 5509 16375 5567 16381
rect 6153 16415 6211 16421
rect 6153 16381 6165 16415
rect 6199 16412 6211 16415
rect 6705 16415 6763 16421
rect 6705 16412 6717 16415
rect 6199 16384 6717 16412
rect 6199 16381 6211 16384
rect 6153 16375 6211 16381
rect 6705 16381 6717 16384
rect 6751 16381 6763 16415
rect 6705 16375 6763 16381
rect 7349 16415 7407 16421
rect 7349 16381 7361 16415
rect 7395 16412 7407 16415
rect 7901 16415 7959 16421
rect 7901 16412 7913 16415
rect 7395 16384 7913 16412
rect 7395 16381 7407 16384
rect 7349 16375 7407 16381
rect 7901 16381 7913 16384
rect 7947 16381 7959 16415
rect 7901 16375 7959 16381
rect 8545 16415 8603 16421
rect 8545 16381 8557 16415
rect 8591 16412 8603 16415
rect 9097 16415 9155 16421
rect 9097 16412 9109 16415
rect 8591 16384 9109 16412
rect 8591 16381 8603 16384
rect 8545 16375 8603 16381
rect 9097 16381 9109 16384
rect 9143 16381 9155 16415
rect 9097 16375 9155 16381
rect 9741 16415 9799 16421
rect 9741 16381 9753 16415
rect 9787 16412 9799 16415
rect 10293 16415 10351 16421
rect 10293 16412 10305 16415
rect 9787 16384 10305 16412
rect 9787 16381 9799 16384
rect 9741 16375 9799 16381
rect 10293 16381 10305 16384
rect 10339 16381 10351 16415
rect 10293 16375 10351 16381
rect 10937 16415 10995 16421
rect 10937 16381 10949 16415
rect 10983 16412 10995 16415
rect 11489 16415 11547 16421
rect 11489 16412 11501 16415
rect 10983 16384 11501 16412
rect 10983 16381 10995 16384
rect 10937 16375 10995 16381
rect 11489 16381 11501 16384
rect 11535 16381 11547 16415
rect 11489 16375 11547 16381
rect 12133 16415 12191 16421
rect 12133 16381 12145 16415
rect 12179 16412 12191 16415
rect 12685 16415 12743 16421
rect 12685 16412 12697 16415
rect 12179 16384 12697 16412
rect 12179 16381 12191 16384
rect 12133 16375 12191 16381
rect 12685 16381 12697 16384
rect 12731 16381 12743 16415
rect 12685 16375 12743 16381
rect 13329 16415 13387 16421
rect 13329 16381 13341 16415
rect 13375 16412 13387 16415
rect 13881 16415 13939 16421
rect 13881 16412 13893 16415
rect 13375 16384 13893 16412
rect 13375 16381 13387 16384
rect 13329 16375 13387 16381
rect 13881 16381 13893 16384
rect 13927 16381 13939 16415
rect 13881 16375 13939 16381
rect 14525 16415 14583 16421
rect 14525 16381 14537 16415
rect 14571 16412 14583 16415
rect 15077 16415 15135 16421
rect 15077 16412 15089 16415
rect 14571 16384 15089 16412
rect 14571 16381 14583 16384
rect 14525 16375 14583 16381
rect 15077 16381 15089 16384
rect 15123 16381 15135 16415
rect 15077 16375 15135 16381
rect 15721 16415 15779 16421
rect 15721 16381 15733 16415
rect 15767 16412 15779 16415
rect 16273 16415 16331 16421
rect 16273 16412 16285 16415
rect 15767 16384 16285 16412
rect 15767 16381 15779 16384
rect 15721 16375 15779 16381
rect 16273 16381 16285 16384
rect 16319 16381 16331 16415
rect 16273 16375 16331 16381
rect 16917 16415 16975 16421
rect 16917 16381 16929 16415
rect 16963 16412 16975 16415
rect 17469 16415 17527 16421
rect 17469 16412 17481 16415
rect 16963 16384 17481 16412
rect 16963 16381 16975 16384
rect 16917 16375 16975 16381
rect 17469 16381 17481 16384
rect 17515 16381 17527 16415
rect 17469 16375 17527 16381
rect 18113 16415 18171 16421
rect 18113 16381 18125 16415
rect 18159 16412 18171 16415
rect 18665 16415 18723 16421
rect 18665 16412 18677 16415
rect 18159 16384 18677 16412
rect 18159 16381 18171 16384
rect 18113 16375 18171 16381
rect 18665 16381 18677 16384
rect 18711 16381 18723 16415
rect 18665 16375 18723 16381
rect 19309 16415 19367 16421
rect 19309 16381 19321 16415
rect 19355 16412 19367 16415
rect 19861 16415 19919 16421
rect 19861 16412 19873 16415
rect 19355 16384 19873 16412
rect 19355 16381 19367 16384
rect 19309 16375 19367 16381
rect 19861 16381 19873 16384
rect 19907 16381 19919 16415
rect 19861 16375 19919 16381
rect 20505 16415 20563 16421
rect 20505 16381 20517 16415
rect 20551 16412 20563 16415
rect 21057 16415 21115 16421
rect 21057 16412 21069 16415
rect 20551 16384 21069 16412
rect 20551 16381 20563 16384
rect 20505 16375 20563 16381
rect 21057 16381 21069 16384
rect 21103 16381 21115 16415
rect 21057 16375 21115 16381
rect 1904 16186 22236 16208
rect 1904 16134 7110 16186
rect 7162 16134 7174 16186
rect 7226 16134 7238 16186
rect 7290 16134 7302 16186
rect 7354 16134 12438 16186
rect 12490 16134 12502 16186
rect 12554 16134 12566 16186
rect 12618 16134 12630 16186
rect 12682 16134 17766 16186
rect 17818 16134 17830 16186
rect 17882 16134 17894 16186
rect 17946 16134 17958 16186
rect 18010 16134 22236 16186
rect 1904 16112 22236 16134
rect 1921 16007 1979 16013
rect 1921 15973 1933 16007
rect 1967 16004 1979 16007
rect 2378 16004 2384 16016
rect 1967 15976 2384 16004
rect 1967 15973 1979 15976
rect 1921 15967 1979 15973
rect 2378 15964 2384 15976
rect 2436 15964 2442 16016
rect 2470 15936 2476 15948
rect 2431 15908 2476 15936
rect 2470 15896 2476 15908
rect 2528 15896 2534 15948
rect 3117 15939 3175 15945
rect 3117 15905 3129 15939
rect 3163 15936 3175 15939
rect 4957 15939 5015 15945
rect 4957 15936 4969 15939
rect 3163 15908 4969 15936
rect 3163 15905 3175 15908
rect 3117 15899 3175 15905
rect 4957 15905 4969 15908
rect 5003 15905 5015 15939
rect 4957 15899 5015 15905
rect 5509 15939 5567 15945
rect 5509 15905 5521 15939
rect 5555 15936 5567 15939
rect 7349 15939 7407 15945
rect 7349 15936 7361 15939
rect 5555 15908 7361 15936
rect 5555 15905 5567 15908
rect 5509 15899 5567 15905
rect 7349 15905 7361 15908
rect 7395 15905 7407 15939
rect 7349 15899 7407 15905
rect 7901 15939 7959 15945
rect 7901 15905 7913 15939
rect 7947 15936 7959 15939
rect 9097 15939 9155 15945
rect 7947 15908 8772 15936
rect 7947 15905 7959 15908
rect 7901 15899 7959 15905
rect 2381 15871 2439 15877
rect 2381 15837 2393 15871
rect 2427 15868 2439 15871
rect 3761 15871 3819 15877
rect 3761 15868 3773 15871
rect 2427 15840 3773 15868
rect 2427 15837 2439 15840
rect 2381 15831 2439 15837
rect 3761 15837 3773 15840
rect 3807 15837 3819 15871
rect 3761 15831 3819 15837
rect 4313 15871 4371 15877
rect 4313 15837 4325 15871
rect 4359 15868 4371 15871
rect 6153 15871 6211 15877
rect 6153 15868 6165 15871
rect 4359 15840 6165 15868
rect 4359 15837 4371 15840
rect 4313 15831 4371 15837
rect 6153 15837 6165 15840
rect 6199 15837 6211 15871
rect 6153 15831 6211 15837
rect 6705 15871 6763 15877
rect 6705 15837 6717 15871
rect 6751 15868 6763 15871
rect 8545 15871 8603 15877
rect 8545 15868 8557 15871
rect 6751 15840 8557 15868
rect 6751 15837 6763 15840
rect 6705 15831 6763 15837
rect 8545 15837 8557 15840
rect 8591 15837 8603 15871
rect 8744 15868 8772 15908
rect 9097 15905 9109 15939
rect 9143 15936 9155 15939
rect 10937 15939 10995 15945
rect 10937 15936 10949 15939
rect 9143 15908 10949 15936
rect 9143 15905 9155 15908
rect 9097 15899 9155 15905
rect 10937 15905 10949 15908
rect 10983 15905 10995 15939
rect 10937 15899 10995 15905
rect 11489 15939 11547 15945
rect 11489 15905 11501 15939
rect 11535 15936 11547 15939
rect 13329 15939 13387 15945
rect 13329 15936 13341 15939
rect 11535 15908 13341 15936
rect 11535 15905 11547 15908
rect 11489 15899 11547 15905
rect 13329 15905 13341 15908
rect 13375 15905 13387 15939
rect 13329 15899 13387 15905
rect 13881 15939 13939 15945
rect 13881 15905 13893 15939
rect 13927 15936 13939 15939
rect 15721 15939 15779 15945
rect 15721 15936 15733 15939
rect 13927 15908 15733 15936
rect 13927 15905 13939 15908
rect 13881 15899 13939 15905
rect 15721 15905 15733 15908
rect 15767 15905 15779 15939
rect 15721 15899 15779 15905
rect 16273 15939 16331 15945
rect 16273 15905 16285 15939
rect 16319 15936 16331 15939
rect 18113 15939 18171 15945
rect 18113 15936 18125 15939
rect 16319 15908 18125 15936
rect 16319 15905 16331 15908
rect 16273 15899 16331 15905
rect 18113 15905 18125 15908
rect 18159 15905 18171 15939
rect 18113 15899 18171 15905
rect 18665 15939 18723 15945
rect 18665 15905 18677 15939
rect 18711 15936 18723 15939
rect 20505 15939 20563 15945
rect 20505 15936 20517 15939
rect 18711 15908 20517 15936
rect 18711 15905 18723 15908
rect 18665 15899 18723 15905
rect 20505 15905 20517 15908
rect 20551 15905 20563 15939
rect 20505 15899 20563 15905
rect 9741 15871 9799 15877
rect 9741 15868 9753 15871
rect 8744 15840 9753 15868
rect 8545 15831 8603 15837
rect 9741 15837 9753 15840
rect 9787 15837 9799 15871
rect 9741 15831 9799 15837
rect 10293 15871 10351 15877
rect 10293 15837 10305 15871
rect 10339 15868 10351 15871
rect 12133 15871 12191 15877
rect 12133 15868 12145 15871
rect 10339 15840 12145 15868
rect 10339 15837 10351 15840
rect 10293 15831 10351 15837
rect 12133 15837 12145 15840
rect 12179 15837 12191 15871
rect 12133 15831 12191 15837
rect 12685 15871 12743 15877
rect 12685 15837 12697 15871
rect 12731 15868 12743 15871
rect 14525 15871 14583 15877
rect 14525 15868 14537 15871
rect 12731 15840 14537 15868
rect 12731 15837 12743 15840
rect 12685 15831 12743 15837
rect 14525 15837 14537 15840
rect 14571 15837 14583 15871
rect 14525 15831 14583 15837
rect 15077 15871 15135 15877
rect 15077 15837 15089 15871
rect 15123 15868 15135 15871
rect 16917 15871 16975 15877
rect 16917 15868 16929 15871
rect 15123 15840 16929 15868
rect 15123 15837 15135 15840
rect 15077 15831 15135 15837
rect 16917 15837 16929 15840
rect 16963 15837 16975 15871
rect 16917 15831 16975 15837
rect 17469 15871 17527 15877
rect 17469 15837 17481 15871
rect 17515 15868 17527 15871
rect 19309 15871 19367 15877
rect 19309 15868 19321 15871
rect 17515 15840 19321 15868
rect 17515 15837 17527 15840
rect 17469 15831 17527 15837
rect 19309 15837 19321 15840
rect 19355 15837 19367 15871
rect 19309 15831 19367 15837
rect 19861 15871 19919 15877
rect 19861 15837 19873 15871
rect 19907 15837 19919 15871
rect 21054 15868 21060 15880
rect 21015 15840 21060 15868
rect 19861 15831 19919 15837
rect 2286 15692 2292 15744
rect 2344 15732 2350 15744
rect 19876 15732 19904 15831
rect 21054 15828 21060 15840
rect 21112 15828 21118 15880
rect 21701 15735 21759 15741
rect 21701 15732 21713 15735
rect 2344 15704 2389 15732
rect 19876 15704 21713 15732
rect 2344 15692 2350 15704
rect 21701 15701 21713 15704
rect 21747 15701 21759 15735
rect 21701 15695 21759 15701
rect 1904 15642 22236 15664
rect 1904 15590 4446 15642
rect 4498 15590 4510 15642
rect 4562 15590 4574 15642
rect 4626 15590 4638 15642
rect 4690 15590 9774 15642
rect 9826 15590 9838 15642
rect 9890 15590 9902 15642
rect 9954 15590 9966 15642
rect 10018 15590 15102 15642
rect 15154 15590 15166 15642
rect 15218 15590 15230 15642
rect 15282 15590 15294 15642
rect 15346 15590 20430 15642
rect 20482 15590 20494 15642
rect 20546 15590 20558 15642
rect 20610 15590 20622 15642
rect 20674 15590 22236 15642
rect 1904 15568 22236 15590
rect 21054 15488 21060 15540
rect 21112 15528 21118 15540
rect 21701 15531 21759 15537
rect 21701 15528 21713 15531
rect 21112 15500 21713 15528
rect 21112 15488 21118 15500
rect 21701 15497 21713 15500
rect 21747 15497 21759 15531
rect 21701 15491 21759 15497
rect 3117 15395 3175 15401
rect 3117 15361 3129 15395
rect 3163 15392 3175 15395
rect 3850 15392 3856 15404
rect 3163 15364 3856 15392
rect 3163 15361 3175 15364
rect 3117 15355 3175 15361
rect 3850 15352 3856 15364
rect 3908 15352 3914 15404
rect 3761 15327 3819 15333
rect 3761 15293 3773 15327
rect 3807 15324 3819 15327
rect 4313 15327 4371 15333
rect 4313 15324 4325 15327
rect 3807 15296 4325 15324
rect 3807 15293 3819 15296
rect 3761 15287 3819 15293
rect 4313 15293 4325 15296
rect 4359 15293 4371 15327
rect 4313 15287 4371 15293
rect 4957 15327 5015 15333
rect 4957 15293 4969 15327
rect 5003 15324 5015 15327
rect 5509 15327 5567 15333
rect 5509 15324 5521 15327
rect 5003 15296 5521 15324
rect 5003 15293 5015 15296
rect 4957 15287 5015 15293
rect 5509 15293 5521 15296
rect 5555 15293 5567 15327
rect 5509 15287 5567 15293
rect 6153 15327 6211 15333
rect 6153 15293 6165 15327
rect 6199 15324 6211 15327
rect 6705 15327 6763 15333
rect 6705 15324 6717 15327
rect 6199 15296 6717 15324
rect 6199 15293 6211 15296
rect 6153 15287 6211 15293
rect 6705 15293 6717 15296
rect 6751 15293 6763 15327
rect 6705 15287 6763 15293
rect 7349 15327 7407 15333
rect 7349 15293 7361 15327
rect 7395 15324 7407 15327
rect 7901 15327 7959 15333
rect 7901 15324 7913 15327
rect 7395 15296 7913 15324
rect 7395 15293 7407 15296
rect 7349 15287 7407 15293
rect 7901 15293 7913 15296
rect 7947 15293 7959 15327
rect 7901 15287 7959 15293
rect 8545 15327 8603 15333
rect 8545 15293 8557 15327
rect 8591 15324 8603 15327
rect 9097 15327 9155 15333
rect 9097 15324 9109 15327
rect 8591 15296 9109 15324
rect 8591 15293 8603 15296
rect 8545 15287 8603 15293
rect 9097 15293 9109 15296
rect 9143 15293 9155 15327
rect 9097 15287 9155 15293
rect 9741 15327 9799 15333
rect 9741 15293 9753 15327
rect 9787 15324 9799 15327
rect 10293 15327 10351 15333
rect 10293 15324 10305 15327
rect 9787 15296 10305 15324
rect 9787 15293 9799 15296
rect 9741 15287 9799 15293
rect 10293 15293 10305 15296
rect 10339 15293 10351 15327
rect 10293 15287 10351 15293
rect 10937 15327 10995 15333
rect 10937 15293 10949 15327
rect 10983 15324 10995 15327
rect 11489 15327 11547 15333
rect 11489 15324 11501 15327
rect 10983 15296 11501 15324
rect 10983 15293 10995 15296
rect 10937 15287 10995 15293
rect 11489 15293 11501 15296
rect 11535 15293 11547 15327
rect 11489 15287 11547 15293
rect 12133 15327 12191 15333
rect 12133 15293 12145 15327
rect 12179 15324 12191 15327
rect 12685 15327 12743 15333
rect 12685 15324 12697 15327
rect 12179 15296 12697 15324
rect 12179 15293 12191 15296
rect 12133 15287 12191 15293
rect 12685 15293 12697 15296
rect 12731 15293 12743 15327
rect 12685 15287 12743 15293
rect 13329 15327 13387 15333
rect 13329 15293 13341 15327
rect 13375 15324 13387 15327
rect 13881 15327 13939 15333
rect 13881 15324 13893 15327
rect 13375 15296 13893 15324
rect 13375 15293 13387 15296
rect 13329 15287 13387 15293
rect 13881 15293 13893 15296
rect 13927 15293 13939 15327
rect 13881 15287 13939 15293
rect 14525 15327 14583 15333
rect 14525 15293 14537 15327
rect 14571 15324 14583 15327
rect 15077 15327 15135 15333
rect 15077 15324 15089 15327
rect 14571 15296 15089 15324
rect 14571 15293 14583 15296
rect 14525 15287 14583 15293
rect 15077 15293 15089 15296
rect 15123 15293 15135 15327
rect 15077 15287 15135 15293
rect 15721 15327 15779 15333
rect 15721 15293 15733 15327
rect 15767 15324 15779 15327
rect 16273 15327 16331 15333
rect 16273 15324 16285 15327
rect 15767 15296 16285 15324
rect 15767 15293 15779 15296
rect 15721 15287 15779 15293
rect 16273 15293 16285 15296
rect 16319 15293 16331 15327
rect 16273 15287 16331 15293
rect 16917 15327 16975 15333
rect 16917 15293 16929 15327
rect 16963 15324 16975 15327
rect 17469 15327 17527 15333
rect 17469 15324 17481 15327
rect 16963 15296 17481 15324
rect 16963 15293 16975 15296
rect 16917 15287 16975 15293
rect 17469 15293 17481 15296
rect 17515 15293 17527 15327
rect 17469 15287 17527 15293
rect 18113 15327 18171 15333
rect 18113 15293 18125 15327
rect 18159 15324 18171 15327
rect 18665 15327 18723 15333
rect 18665 15324 18677 15327
rect 18159 15296 18677 15324
rect 18159 15293 18171 15296
rect 18113 15287 18171 15293
rect 18665 15293 18677 15296
rect 18711 15293 18723 15327
rect 18665 15287 18723 15293
rect 19309 15327 19367 15333
rect 19309 15293 19321 15327
rect 19355 15324 19367 15327
rect 19861 15327 19919 15333
rect 19861 15324 19873 15327
rect 19355 15296 19873 15324
rect 19355 15293 19367 15296
rect 19309 15287 19367 15293
rect 19861 15293 19873 15296
rect 19907 15293 19919 15327
rect 19861 15287 19919 15293
rect 20505 15327 20563 15333
rect 20505 15293 20517 15327
rect 20551 15324 20563 15327
rect 21057 15327 21115 15333
rect 21057 15324 21069 15327
rect 20551 15296 21069 15324
rect 20551 15293 20563 15296
rect 20505 15287 20563 15293
rect 21057 15293 21069 15296
rect 21103 15293 21115 15327
rect 21057 15287 21115 15293
rect 1904 15098 22236 15120
rect 1904 15046 7110 15098
rect 7162 15046 7174 15098
rect 7226 15046 7238 15098
rect 7290 15046 7302 15098
rect 7354 15046 12438 15098
rect 12490 15046 12502 15098
rect 12554 15046 12566 15098
rect 12618 15046 12630 15098
rect 12682 15046 17766 15098
rect 17818 15046 17830 15098
rect 17882 15046 17894 15098
rect 17946 15046 17958 15098
rect 18010 15046 22236 15098
rect 1904 15024 22236 15046
rect 3761 14987 3819 14993
rect 3761 14953 3773 14987
rect 3807 14984 3819 14987
rect 3850 14984 3856 14996
rect 3807 14956 3856 14984
rect 3807 14953 3819 14956
rect 3761 14947 3819 14953
rect 3850 14944 3856 14956
rect 3908 14944 3914 14996
rect 3117 14851 3175 14857
rect 3117 14817 3129 14851
rect 3163 14848 3175 14851
rect 4957 14851 5015 14857
rect 4957 14848 4969 14851
rect 3163 14820 4969 14848
rect 3163 14817 3175 14820
rect 3117 14811 3175 14817
rect 4957 14817 4969 14820
rect 5003 14817 5015 14851
rect 4957 14811 5015 14817
rect 5509 14851 5567 14857
rect 5509 14817 5521 14851
rect 5555 14848 5567 14851
rect 7349 14851 7407 14857
rect 7349 14848 7361 14851
rect 5555 14820 7361 14848
rect 5555 14817 5567 14820
rect 5509 14811 5567 14817
rect 7349 14817 7361 14820
rect 7395 14817 7407 14851
rect 7349 14811 7407 14817
rect 7901 14851 7959 14857
rect 7901 14817 7913 14851
rect 7947 14848 7959 14851
rect 9097 14851 9155 14857
rect 7947 14820 8772 14848
rect 7947 14817 7959 14820
rect 7901 14811 7959 14817
rect 4313 14783 4371 14789
rect 4313 14749 4325 14783
rect 4359 14780 4371 14783
rect 6153 14783 6211 14789
rect 6153 14780 6165 14783
rect 4359 14752 6165 14780
rect 4359 14749 4371 14752
rect 4313 14743 4371 14749
rect 6153 14749 6165 14752
rect 6199 14749 6211 14783
rect 6153 14743 6211 14749
rect 6705 14783 6763 14789
rect 6705 14749 6717 14783
rect 6751 14780 6763 14783
rect 8545 14783 8603 14789
rect 8545 14780 8557 14783
rect 6751 14752 8557 14780
rect 6751 14749 6763 14752
rect 6705 14743 6763 14749
rect 8545 14749 8557 14752
rect 8591 14749 8603 14783
rect 8744 14780 8772 14820
rect 9097 14817 9109 14851
rect 9143 14848 9155 14851
rect 10937 14851 10995 14857
rect 10937 14848 10949 14851
rect 9143 14820 10949 14848
rect 9143 14817 9155 14820
rect 9097 14811 9155 14817
rect 10937 14817 10949 14820
rect 10983 14817 10995 14851
rect 10937 14811 10995 14817
rect 11489 14851 11547 14857
rect 11489 14817 11501 14851
rect 11535 14848 11547 14851
rect 13329 14851 13387 14857
rect 13329 14848 13341 14851
rect 11535 14820 13341 14848
rect 11535 14817 11547 14820
rect 11489 14811 11547 14817
rect 13329 14817 13341 14820
rect 13375 14817 13387 14851
rect 13329 14811 13387 14817
rect 13881 14851 13939 14857
rect 13881 14817 13893 14851
rect 13927 14848 13939 14851
rect 15721 14851 15779 14857
rect 15721 14848 15733 14851
rect 13927 14820 15733 14848
rect 13927 14817 13939 14820
rect 13881 14811 13939 14817
rect 15721 14817 15733 14820
rect 15767 14817 15779 14851
rect 15721 14811 15779 14817
rect 16273 14851 16331 14857
rect 16273 14817 16285 14851
rect 16319 14848 16331 14851
rect 18113 14851 18171 14857
rect 18113 14848 18125 14851
rect 16319 14820 18125 14848
rect 16319 14817 16331 14820
rect 16273 14811 16331 14817
rect 18113 14817 18125 14820
rect 18159 14817 18171 14851
rect 18113 14811 18171 14817
rect 18665 14851 18723 14857
rect 18665 14817 18677 14851
rect 18711 14848 18723 14851
rect 20505 14851 20563 14857
rect 20505 14848 20517 14851
rect 18711 14820 20517 14848
rect 18711 14817 18723 14820
rect 18665 14811 18723 14817
rect 20505 14817 20517 14820
rect 20551 14817 20563 14851
rect 20505 14811 20563 14817
rect 9741 14783 9799 14789
rect 9741 14780 9753 14783
rect 8744 14752 9753 14780
rect 8545 14743 8603 14749
rect 9741 14749 9753 14752
rect 9787 14749 9799 14783
rect 9741 14743 9799 14749
rect 10293 14783 10351 14789
rect 10293 14749 10305 14783
rect 10339 14780 10351 14783
rect 12133 14783 12191 14789
rect 12133 14780 12145 14783
rect 10339 14752 12145 14780
rect 10339 14749 10351 14752
rect 10293 14743 10351 14749
rect 12133 14749 12145 14752
rect 12179 14749 12191 14783
rect 12133 14743 12191 14749
rect 12685 14783 12743 14789
rect 12685 14749 12697 14783
rect 12731 14780 12743 14783
rect 14525 14783 14583 14789
rect 14525 14780 14537 14783
rect 12731 14752 14537 14780
rect 12731 14749 12743 14752
rect 12685 14743 12743 14749
rect 14525 14749 14537 14752
rect 14571 14749 14583 14783
rect 14525 14743 14583 14749
rect 15077 14783 15135 14789
rect 15077 14749 15089 14783
rect 15123 14780 15135 14783
rect 16917 14783 16975 14789
rect 16917 14780 16929 14783
rect 15123 14752 16929 14780
rect 15123 14749 15135 14752
rect 15077 14743 15135 14749
rect 16917 14749 16929 14752
rect 16963 14749 16975 14783
rect 16917 14743 16975 14749
rect 17469 14783 17527 14789
rect 17469 14749 17481 14783
rect 17515 14780 17527 14783
rect 19309 14783 19367 14789
rect 19309 14780 19321 14783
rect 17515 14752 19321 14780
rect 17515 14749 17527 14752
rect 17469 14743 17527 14749
rect 19309 14749 19321 14752
rect 19355 14749 19367 14783
rect 19309 14743 19367 14749
rect 19861 14783 19919 14789
rect 19861 14749 19873 14783
rect 19907 14749 19919 14783
rect 19861 14743 19919 14749
rect 21057 14783 21115 14789
rect 21057 14749 21069 14783
rect 21103 14780 21115 14783
rect 21606 14780 21612 14792
rect 21103 14752 21612 14780
rect 21103 14749 21115 14752
rect 21057 14743 21115 14749
rect 19876 14644 19904 14743
rect 21606 14740 21612 14752
rect 21664 14740 21670 14792
rect 21701 14647 21759 14653
rect 21701 14644 21713 14647
rect 19876 14616 21713 14644
rect 21701 14613 21713 14616
rect 21747 14613 21759 14647
rect 21701 14607 21759 14613
rect 1904 14554 22236 14576
rect 1904 14502 4446 14554
rect 4498 14502 4510 14554
rect 4562 14502 4574 14554
rect 4626 14502 4638 14554
rect 4690 14502 9774 14554
rect 9826 14502 9838 14554
rect 9890 14502 9902 14554
rect 9954 14502 9966 14554
rect 10018 14502 15102 14554
rect 15154 14502 15166 14554
rect 15218 14502 15230 14554
rect 15282 14502 15294 14554
rect 15346 14502 20430 14554
rect 20482 14502 20494 14554
rect 20546 14502 20558 14554
rect 20610 14502 20622 14554
rect 20674 14502 22236 14554
rect 1904 14480 22236 14502
rect 21606 14400 21612 14452
rect 21664 14440 21670 14452
rect 21701 14443 21759 14449
rect 21701 14440 21713 14443
rect 21664 14412 21713 14440
rect 21664 14400 21670 14412
rect 21701 14409 21713 14412
rect 21747 14409 21759 14443
rect 21701 14403 21759 14409
rect 2286 14264 2292 14316
rect 2344 14304 2350 14316
rect 3117 14307 3175 14313
rect 3117 14304 3129 14307
rect 2344 14276 3129 14304
rect 2344 14264 2350 14276
rect 3117 14273 3129 14276
rect 3163 14273 3175 14307
rect 3117 14267 3175 14273
rect 3761 14239 3819 14245
rect 3761 14205 3773 14239
rect 3807 14236 3819 14239
rect 4313 14239 4371 14245
rect 4313 14236 4325 14239
rect 3807 14208 4325 14236
rect 3807 14205 3819 14208
rect 3761 14199 3819 14205
rect 4313 14205 4325 14208
rect 4359 14205 4371 14239
rect 4313 14199 4371 14205
rect 4957 14239 5015 14245
rect 4957 14205 4969 14239
rect 5003 14236 5015 14239
rect 5509 14239 5567 14245
rect 5509 14236 5521 14239
rect 5003 14208 5521 14236
rect 5003 14205 5015 14208
rect 4957 14199 5015 14205
rect 5509 14205 5521 14208
rect 5555 14205 5567 14239
rect 5509 14199 5567 14205
rect 6153 14239 6211 14245
rect 6153 14205 6165 14239
rect 6199 14236 6211 14239
rect 6705 14239 6763 14245
rect 6705 14236 6717 14239
rect 6199 14208 6717 14236
rect 6199 14205 6211 14208
rect 6153 14199 6211 14205
rect 6705 14205 6717 14208
rect 6751 14205 6763 14239
rect 6705 14199 6763 14205
rect 7349 14239 7407 14245
rect 7349 14205 7361 14239
rect 7395 14236 7407 14239
rect 7901 14239 7959 14245
rect 7901 14236 7913 14239
rect 7395 14208 7913 14236
rect 7395 14205 7407 14208
rect 7349 14199 7407 14205
rect 7901 14205 7913 14208
rect 7947 14205 7959 14239
rect 7901 14199 7959 14205
rect 8545 14239 8603 14245
rect 8545 14205 8557 14239
rect 8591 14236 8603 14239
rect 9097 14239 9155 14245
rect 9097 14236 9109 14239
rect 8591 14208 9109 14236
rect 8591 14205 8603 14208
rect 8545 14199 8603 14205
rect 9097 14205 9109 14208
rect 9143 14205 9155 14239
rect 9097 14199 9155 14205
rect 9741 14239 9799 14245
rect 9741 14205 9753 14239
rect 9787 14236 9799 14239
rect 10293 14239 10351 14245
rect 10293 14236 10305 14239
rect 9787 14208 10305 14236
rect 9787 14205 9799 14208
rect 9741 14199 9799 14205
rect 10293 14205 10305 14208
rect 10339 14205 10351 14239
rect 10293 14199 10351 14205
rect 10937 14239 10995 14245
rect 10937 14205 10949 14239
rect 10983 14236 10995 14239
rect 11489 14239 11547 14245
rect 11489 14236 11501 14239
rect 10983 14208 11501 14236
rect 10983 14205 10995 14208
rect 10937 14199 10995 14205
rect 11489 14205 11501 14208
rect 11535 14205 11547 14239
rect 11489 14199 11547 14205
rect 12133 14239 12191 14245
rect 12133 14205 12145 14239
rect 12179 14236 12191 14239
rect 12685 14239 12743 14245
rect 12685 14236 12697 14239
rect 12179 14208 12697 14236
rect 12179 14205 12191 14208
rect 12133 14199 12191 14205
rect 12685 14205 12697 14208
rect 12731 14205 12743 14239
rect 12685 14199 12743 14205
rect 13329 14239 13387 14245
rect 13329 14205 13341 14239
rect 13375 14236 13387 14239
rect 13881 14239 13939 14245
rect 13881 14236 13893 14239
rect 13375 14208 13893 14236
rect 13375 14205 13387 14208
rect 13329 14199 13387 14205
rect 13881 14205 13893 14208
rect 13927 14205 13939 14239
rect 13881 14199 13939 14205
rect 14525 14239 14583 14245
rect 14525 14205 14537 14239
rect 14571 14236 14583 14239
rect 15077 14239 15135 14245
rect 15077 14236 15089 14239
rect 14571 14208 15089 14236
rect 14571 14205 14583 14208
rect 14525 14199 14583 14205
rect 15077 14205 15089 14208
rect 15123 14205 15135 14239
rect 15077 14199 15135 14205
rect 15721 14239 15779 14245
rect 15721 14205 15733 14239
rect 15767 14236 15779 14239
rect 16273 14239 16331 14245
rect 16273 14236 16285 14239
rect 15767 14208 16285 14236
rect 15767 14205 15779 14208
rect 15721 14199 15779 14205
rect 16273 14205 16285 14208
rect 16319 14205 16331 14239
rect 16273 14199 16331 14205
rect 16917 14239 16975 14245
rect 16917 14205 16929 14239
rect 16963 14236 16975 14239
rect 17469 14239 17527 14245
rect 17469 14236 17481 14239
rect 16963 14208 17481 14236
rect 16963 14205 16975 14208
rect 16917 14199 16975 14205
rect 17469 14205 17481 14208
rect 17515 14205 17527 14239
rect 17469 14199 17527 14205
rect 18113 14239 18171 14245
rect 18113 14205 18125 14239
rect 18159 14236 18171 14239
rect 18665 14239 18723 14245
rect 18665 14236 18677 14239
rect 18159 14208 18677 14236
rect 18159 14205 18171 14208
rect 18113 14199 18171 14205
rect 18665 14205 18677 14208
rect 18711 14205 18723 14239
rect 18665 14199 18723 14205
rect 19309 14239 19367 14245
rect 19309 14205 19321 14239
rect 19355 14236 19367 14239
rect 19861 14239 19919 14245
rect 19861 14236 19873 14239
rect 19355 14208 19873 14236
rect 19355 14205 19367 14208
rect 19309 14199 19367 14205
rect 19861 14205 19873 14208
rect 19907 14205 19919 14239
rect 19861 14199 19919 14205
rect 20505 14239 20563 14245
rect 20505 14205 20517 14239
rect 20551 14236 20563 14239
rect 21057 14239 21115 14245
rect 21057 14236 21069 14239
rect 20551 14208 21069 14236
rect 20551 14205 20563 14208
rect 20505 14199 20563 14205
rect 21057 14205 21069 14208
rect 21103 14205 21115 14239
rect 21057 14199 21115 14205
rect 1904 14010 22236 14032
rect 1904 13958 7110 14010
rect 7162 13958 7174 14010
rect 7226 13958 7238 14010
rect 7290 13958 7302 14010
rect 7354 13958 12438 14010
rect 12490 13958 12502 14010
rect 12554 13958 12566 14010
rect 12618 13958 12630 14010
rect 12682 13958 17766 14010
rect 17818 13958 17830 14010
rect 17882 13958 17894 14010
rect 17946 13958 17958 14010
rect 18010 13958 22236 14010
rect 1904 13936 22236 13958
rect 1921 13831 1979 13837
rect 1921 13797 1933 13831
rect 1967 13828 1979 13831
rect 2286 13828 2292 13840
rect 1967 13800 2292 13828
rect 1967 13797 1979 13800
rect 1921 13791 1979 13797
rect 2286 13788 2292 13800
rect 2344 13788 2350 13840
rect 2470 13760 2476 13772
rect 2431 13732 2476 13760
rect 2470 13720 2476 13732
rect 2528 13720 2534 13772
rect 3117 13763 3175 13769
rect 3117 13729 3129 13763
rect 3163 13760 3175 13763
rect 4957 13763 5015 13769
rect 4957 13760 4969 13763
rect 3163 13732 4969 13760
rect 3163 13729 3175 13732
rect 3117 13723 3175 13729
rect 4957 13729 4969 13732
rect 5003 13729 5015 13763
rect 4957 13723 5015 13729
rect 5509 13763 5567 13769
rect 5509 13729 5521 13763
rect 5555 13760 5567 13763
rect 7349 13763 7407 13769
rect 7349 13760 7361 13763
rect 5555 13732 7361 13760
rect 5555 13729 5567 13732
rect 5509 13723 5567 13729
rect 7349 13729 7361 13732
rect 7395 13729 7407 13763
rect 7349 13723 7407 13729
rect 7901 13763 7959 13769
rect 7901 13729 7913 13763
rect 7947 13760 7959 13763
rect 9097 13763 9155 13769
rect 7947 13732 8772 13760
rect 7947 13729 7959 13732
rect 7901 13723 7959 13729
rect 4313 13695 4371 13701
rect 4313 13661 4325 13695
rect 4359 13692 4371 13695
rect 6153 13695 6211 13701
rect 6153 13692 6165 13695
rect 4359 13664 6165 13692
rect 4359 13661 4371 13664
rect 4313 13655 4371 13661
rect 6153 13661 6165 13664
rect 6199 13661 6211 13695
rect 6153 13655 6211 13661
rect 6705 13695 6763 13701
rect 6705 13661 6717 13695
rect 6751 13692 6763 13695
rect 8545 13695 8603 13701
rect 8545 13692 8557 13695
rect 6751 13664 8557 13692
rect 6751 13661 6763 13664
rect 6705 13655 6763 13661
rect 8545 13661 8557 13664
rect 8591 13661 8603 13695
rect 8744 13692 8772 13732
rect 9097 13729 9109 13763
rect 9143 13760 9155 13763
rect 10937 13763 10995 13769
rect 10937 13760 10949 13763
rect 9143 13732 10949 13760
rect 9143 13729 9155 13732
rect 9097 13723 9155 13729
rect 10937 13729 10949 13732
rect 10983 13729 10995 13763
rect 10937 13723 10995 13729
rect 11489 13763 11547 13769
rect 11489 13729 11501 13763
rect 11535 13760 11547 13763
rect 13329 13763 13387 13769
rect 13329 13760 13341 13763
rect 11535 13732 13341 13760
rect 11535 13729 11547 13732
rect 11489 13723 11547 13729
rect 13329 13729 13341 13732
rect 13375 13729 13387 13763
rect 13329 13723 13387 13729
rect 13881 13763 13939 13769
rect 13881 13729 13893 13763
rect 13927 13760 13939 13763
rect 15721 13763 15779 13769
rect 15721 13760 15733 13763
rect 13927 13732 15733 13760
rect 13927 13729 13939 13732
rect 13881 13723 13939 13729
rect 15721 13729 15733 13732
rect 15767 13729 15779 13763
rect 15721 13723 15779 13729
rect 16273 13763 16331 13769
rect 16273 13729 16285 13763
rect 16319 13760 16331 13763
rect 18113 13763 18171 13769
rect 18113 13760 18125 13763
rect 16319 13732 18125 13760
rect 16319 13729 16331 13732
rect 16273 13723 16331 13729
rect 18113 13729 18125 13732
rect 18159 13729 18171 13763
rect 18113 13723 18171 13729
rect 18665 13763 18723 13769
rect 18665 13729 18677 13763
rect 18711 13760 18723 13763
rect 20505 13763 20563 13769
rect 20505 13760 20517 13763
rect 18711 13732 20517 13760
rect 18711 13729 18723 13732
rect 18665 13723 18723 13729
rect 20505 13729 20517 13732
rect 20551 13729 20563 13763
rect 20505 13723 20563 13729
rect 9741 13695 9799 13701
rect 9741 13692 9753 13695
rect 8744 13664 9753 13692
rect 8545 13655 8603 13661
rect 9741 13661 9753 13664
rect 9787 13661 9799 13695
rect 9741 13655 9799 13661
rect 10293 13695 10351 13701
rect 10293 13661 10305 13695
rect 10339 13692 10351 13695
rect 12133 13695 12191 13701
rect 12133 13692 12145 13695
rect 10339 13664 12145 13692
rect 10339 13661 10351 13664
rect 10293 13655 10351 13661
rect 12133 13661 12145 13664
rect 12179 13661 12191 13695
rect 12133 13655 12191 13661
rect 12685 13695 12743 13701
rect 12685 13661 12697 13695
rect 12731 13692 12743 13695
rect 14525 13695 14583 13701
rect 14525 13692 14537 13695
rect 12731 13664 14537 13692
rect 12731 13661 12743 13664
rect 12685 13655 12743 13661
rect 14525 13661 14537 13664
rect 14571 13661 14583 13695
rect 14525 13655 14583 13661
rect 15077 13695 15135 13701
rect 15077 13661 15089 13695
rect 15123 13692 15135 13695
rect 16917 13695 16975 13701
rect 16917 13692 16929 13695
rect 15123 13664 16929 13692
rect 15123 13661 15135 13664
rect 15077 13655 15135 13661
rect 16917 13661 16929 13664
rect 16963 13661 16975 13695
rect 16917 13655 16975 13661
rect 17469 13695 17527 13701
rect 17469 13661 17481 13695
rect 17515 13692 17527 13695
rect 19309 13695 19367 13701
rect 19309 13692 19321 13695
rect 17515 13664 19321 13692
rect 17515 13661 17527 13664
rect 17469 13655 17527 13661
rect 19309 13661 19321 13664
rect 19355 13661 19367 13695
rect 19309 13655 19367 13661
rect 19861 13695 19919 13701
rect 19861 13661 19873 13695
rect 19907 13661 19919 13695
rect 21054 13692 21060 13704
rect 21015 13664 21060 13692
rect 19861 13655 19919 13661
rect 2381 13627 2439 13633
rect 2381 13593 2393 13627
rect 2427 13624 2439 13627
rect 3761 13627 3819 13633
rect 3761 13624 3773 13627
rect 2427 13596 3773 13624
rect 2427 13593 2439 13596
rect 2381 13587 2439 13593
rect 3761 13593 3773 13596
rect 3807 13593 3819 13627
rect 3761 13587 3819 13593
rect 2286 13516 2292 13568
rect 2344 13556 2350 13568
rect 19876 13556 19904 13655
rect 21054 13652 21060 13664
rect 21112 13652 21118 13704
rect 21701 13559 21759 13565
rect 21701 13556 21713 13559
rect 2344 13528 2389 13556
rect 19876 13528 21713 13556
rect 2344 13516 2350 13528
rect 21701 13525 21713 13528
rect 21747 13525 21759 13559
rect 21701 13519 21759 13525
rect 1904 13466 22236 13488
rect 1904 13414 4446 13466
rect 4498 13414 4510 13466
rect 4562 13414 4574 13466
rect 4626 13414 4638 13466
rect 4690 13414 9774 13466
rect 9826 13414 9838 13466
rect 9890 13414 9902 13466
rect 9954 13414 9966 13466
rect 10018 13414 15102 13466
rect 15154 13414 15166 13466
rect 15218 13414 15230 13466
rect 15282 13414 15294 13466
rect 15346 13414 20430 13466
rect 20482 13414 20494 13466
rect 20546 13414 20558 13466
rect 20610 13414 20622 13466
rect 20674 13414 22236 13466
rect 1904 13392 22236 13414
rect 21054 13312 21060 13364
rect 21112 13352 21118 13364
rect 21701 13355 21759 13361
rect 21701 13352 21713 13355
rect 21112 13324 21713 13352
rect 21112 13312 21118 13324
rect 21701 13321 21713 13324
rect 21747 13321 21759 13355
rect 21701 13315 21759 13321
rect 3117 13219 3175 13225
rect 3117 13185 3129 13219
rect 3163 13216 3175 13219
rect 3850 13216 3856 13228
rect 3163 13188 3856 13216
rect 3163 13185 3175 13188
rect 3117 13179 3175 13185
rect 3850 13176 3856 13188
rect 3908 13176 3914 13228
rect 3761 13151 3819 13157
rect 3761 13117 3773 13151
rect 3807 13148 3819 13151
rect 4313 13151 4371 13157
rect 4313 13148 4325 13151
rect 3807 13120 4325 13148
rect 3807 13117 3819 13120
rect 3761 13111 3819 13117
rect 4313 13117 4325 13120
rect 4359 13117 4371 13151
rect 4313 13111 4371 13117
rect 4957 13151 5015 13157
rect 4957 13117 4969 13151
rect 5003 13148 5015 13151
rect 5509 13151 5567 13157
rect 5509 13148 5521 13151
rect 5003 13120 5521 13148
rect 5003 13117 5015 13120
rect 4957 13111 5015 13117
rect 5509 13117 5521 13120
rect 5555 13117 5567 13151
rect 5509 13111 5567 13117
rect 6153 13151 6211 13157
rect 6153 13117 6165 13151
rect 6199 13148 6211 13151
rect 6705 13151 6763 13157
rect 6705 13148 6717 13151
rect 6199 13120 6717 13148
rect 6199 13117 6211 13120
rect 6153 13111 6211 13117
rect 6705 13117 6717 13120
rect 6751 13117 6763 13151
rect 6705 13111 6763 13117
rect 7349 13151 7407 13157
rect 7349 13117 7361 13151
rect 7395 13148 7407 13151
rect 7901 13151 7959 13157
rect 7901 13148 7913 13151
rect 7395 13120 7913 13148
rect 7395 13117 7407 13120
rect 7349 13111 7407 13117
rect 7901 13117 7913 13120
rect 7947 13117 7959 13151
rect 7901 13111 7959 13117
rect 8545 13151 8603 13157
rect 8545 13117 8557 13151
rect 8591 13148 8603 13151
rect 9097 13151 9155 13157
rect 9097 13148 9109 13151
rect 8591 13120 9109 13148
rect 8591 13117 8603 13120
rect 8545 13111 8603 13117
rect 9097 13117 9109 13120
rect 9143 13117 9155 13151
rect 9097 13111 9155 13117
rect 9741 13151 9799 13157
rect 9741 13117 9753 13151
rect 9787 13148 9799 13151
rect 10293 13151 10351 13157
rect 10293 13148 10305 13151
rect 9787 13120 10305 13148
rect 9787 13117 9799 13120
rect 9741 13111 9799 13117
rect 10293 13117 10305 13120
rect 10339 13117 10351 13151
rect 10293 13111 10351 13117
rect 10937 13151 10995 13157
rect 10937 13117 10949 13151
rect 10983 13148 10995 13151
rect 11489 13151 11547 13157
rect 11489 13148 11501 13151
rect 10983 13120 11501 13148
rect 10983 13117 10995 13120
rect 10937 13111 10995 13117
rect 11489 13117 11501 13120
rect 11535 13117 11547 13151
rect 11489 13111 11547 13117
rect 12133 13151 12191 13157
rect 12133 13117 12145 13151
rect 12179 13148 12191 13151
rect 12685 13151 12743 13157
rect 12685 13148 12697 13151
rect 12179 13120 12697 13148
rect 12179 13117 12191 13120
rect 12133 13111 12191 13117
rect 12685 13117 12697 13120
rect 12731 13117 12743 13151
rect 12685 13111 12743 13117
rect 13329 13151 13387 13157
rect 13329 13117 13341 13151
rect 13375 13148 13387 13151
rect 13881 13151 13939 13157
rect 13881 13148 13893 13151
rect 13375 13120 13893 13148
rect 13375 13117 13387 13120
rect 13329 13111 13387 13117
rect 13881 13117 13893 13120
rect 13927 13117 13939 13151
rect 13881 13111 13939 13117
rect 14525 13151 14583 13157
rect 14525 13117 14537 13151
rect 14571 13148 14583 13151
rect 15077 13151 15135 13157
rect 15077 13148 15089 13151
rect 14571 13120 15089 13148
rect 14571 13117 14583 13120
rect 14525 13111 14583 13117
rect 15077 13117 15089 13120
rect 15123 13117 15135 13151
rect 15077 13111 15135 13117
rect 15721 13151 15779 13157
rect 15721 13117 15733 13151
rect 15767 13148 15779 13151
rect 16273 13151 16331 13157
rect 16273 13148 16285 13151
rect 15767 13120 16285 13148
rect 15767 13117 15779 13120
rect 15721 13111 15779 13117
rect 16273 13117 16285 13120
rect 16319 13117 16331 13151
rect 16273 13111 16331 13117
rect 16917 13151 16975 13157
rect 16917 13117 16929 13151
rect 16963 13148 16975 13151
rect 17469 13151 17527 13157
rect 17469 13148 17481 13151
rect 16963 13120 17481 13148
rect 16963 13117 16975 13120
rect 16917 13111 16975 13117
rect 17469 13117 17481 13120
rect 17515 13117 17527 13151
rect 17469 13111 17527 13117
rect 18113 13151 18171 13157
rect 18113 13117 18125 13151
rect 18159 13148 18171 13151
rect 18665 13151 18723 13157
rect 18665 13148 18677 13151
rect 18159 13120 18677 13148
rect 18159 13117 18171 13120
rect 18113 13111 18171 13117
rect 18665 13117 18677 13120
rect 18711 13117 18723 13151
rect 18665 13111 18723 13117
rect 19309 13151 19367 13157
rect 19309 13117 19321 13151
rect 19355 13148 19367 13151
rect 19861 13151 19919 13157
rect 19861 13148 19873 13151
rect 19355 13120 19873 13148
rect 19355 13117 19367 13120
rect 19309 13111 19367 13117
rect 19861 13117 19873 13120
rect 19907 13117 19919 13151
rect 19861 13111 19919 13117
rect 20505 13151 20563 13157
rect 20505 13117 20517 13151
rect 20551 13148 20563 13151
rect 21057 13151 21115 13157
rect 21057 13148 21069 13151
rect 20551 13120 21069 13148
rect 20551 13117 20563 13120
rect 20505 13111 20563 13117
rect 21057 13117 21069 13120
rect 21103 13117 21115 13151
rect 21057 13111 21115 13117
rect 1904 12922 22236 12944
rect 1904 12870 7110 12922
rect 7162 12870 7174 12922
rect 7226 12870 7238 12922
rect 7290 12870 7302 12922
rect 7354 12870 12438 12922
rect 12490 12870 12502 12922
rect 12554 12870 12566 12922
rect 12618 12870 12630 12922
rect 12682 12870 17766 12922
rect 17818 12870 17830 12922
rect 17882 12870 17894 12922
rect 17946 12870 17958 12922
rect 18010 12870 22236 12922
rect 1904 12848 22236 12870
rect 3761 12811 3819 12817
rect 3761 12777 3773 12811
rect 3807 12808 3819 12811
rect 3850 12808 3856 12820
rect 3807 12780 3856 12808
rect 3807 12777 3819 12780
rect 3761 12771 3819 12777
rect 3850 12768 3856 12780
rect 3908 12768 3914 12820
rect 3117 12675 3175 12681
rect 3117 12641 3129 12675
rect 3163 12672 3175 12675
rect 4957 12675 5015 12681
rect 4957 12672 4969 12675
rect 3163 12644 4969 12672
rect 3163 12641 3175 12644
rect 3117 12635 3175 12641
rect 4957 12641 4969 12644
rect 5003 12641 5015 12675
rect 4957 12635 5015 12641
rect 5509 12675 5567 12681
rect 5509 12641 5521 12675
rect 5555 12672 5567 12675
rect 7349 12675 7407 12681
rect 7349 12672 7361 12675
rect 5555 12644 7361 12672
rect 5555 12641 5567 12644
rect 5509 12635 5567 12641
rect 7349 12641 7361 12644
rect 7395 12641 7407 12675
rect 7349 12635 7407 12641
rect 7901 12675 7959 12681
rect 7901 12641 7913 12675
rect 7947 12672 7959 12675
rect 9097 12675 9155 12681
rect 7947 12644 8772 12672
rect 7947 12641 7959 12644
rect 7901 12635 7959 12641
rect 4313 12607 4371 12613
rect 4313 12573 4325 12607
rect 4359 12604 4371 12607
rect 6153 12607 6211 12613
rect 6153 12604 6165 12607
rect 4359 12576 6165 12604
rect 4359 12573 4371 12576
rect 4313 12567 4371 12573
rect 6153 12573 6165 12576
rect 6199 12573 6211 12607
rect 6153 12567 6211 12573
rect 6705 12607 6763 12613
rect 6705 12573 6717 12607
rect 6751 12604 6763 12607
rect 8545 12607 8603 12613
rect 8545 12604 8557 12607
rect 6751 12576 8557 12604
rect 6751 12573 6763 12576
rect 6705 12567 6763 12573
rect 8545 12573 8557 12576
rect 8591 12573 8603 12607
rect 8744 12604 8772 12644
rect 9097 12641 9109 12675
rect 9143 12672 9155 12675
rect 10937 12675 10995 12681
rect 10937 12672 10949 12675
rect 9143 12644 10949 12672
rect 9143 12641 9155 12644
rect 9097 12635 9155 12641
rect 10937 12641 10949 12644
rect 10983 12641 10995 12675
rect 10937 12635 10995 12641
rect 11489 12675 11547 12681
rect 11489 12641 11501 12675
rect 11535 12672 11547 12675
rect 13329 12675 13387 12681
rect 13329 12672 13341 12675
rect 11535 12644 13341 12672
rect 11535 12641 11547 12644
rect 11489 12635 11547 12641
rect 13329 12641 13341 12644
rect 13375 12641 13387 12675
rect 13329 12635 13387 12641
rect 13881 12675 13939 12681
rect 13881 12641 13893 12675
rect 13927 12672 13939 12675
rect 15721 12675 15779 12681
rect 15721 12672 15733 12675
rect 13927 12644 15733 12672
rect 13927 12641 13939 12644
rect 13881 12635 13939 12641
rect 15721 12641 15733 12644
rect 15767 12641 15779 12675
rect 15721 12635 15779 12641
rect 16273 12675 16331 12681
rect 16273 12641 16285 12675
rect 16319 12672 16331 12675
rect 18113 12675 18171 12681
rect 18113 12672 18125 12675
rect 16319 12644 18125 12672
rect 16319 12641 16331 12644
rect 16273 12635 16331 12641
rect 18113 12641 18125 12644
rect 18159 12641 18171 12675
rect 18113 12635 18171 12641
rect 18665 12675 18723 12681
rect 18665 12641 18677 12675
rect 18711 12672 18723 12675
rect 20505 12675 20563 12681
rect 20505 12672 20517 12675
rect 18711 12644 20517 12672
rect 18711 12641 18723 12644
rect 18665 12635 18723 12641
rect 20505 12641 20517 12644
rect 20551 12641 20563 12675
rect 20505 12635 20563 12641
rect 9741 12607 9799 12613
rect 9741 12604 9753 12607
rect 8744 12576 9753 12604
rect 8545 12567 8603 12573
rect 9741 12573 9753 12576
rect 9787 12573 9799 12607
rect 9741 12567 9799 12573
rect 10293 12607 10351 12613
rect 10293 12573 10305 12607
rect 10339 12604 10351 12607
rect 12133 12607 12191 12613
rect 12133 12604 12145 12607
rect 10339 12576 12145 12604
rect 10339 12573 10351 12576
rect 10293 12567 10351 12573
rect 12133 12573 12145 12576
rect 12179 12573 12191 12607
rect 12133 12567 12191 12573
rect 12685 12607 12743 12613
rect 12685 12573 12697 12607
rect 12731 12604 12743 12607
rect 14525 12607 14583 12613
rect 14525 12604 14537 12607
rect 12731 12576 14537 12604
rect 12731 12573 12743 12576
rect 12685 12567 12743 12573
rect 14525 12573 14537 12576
rect 14571 12573 14583 12607
rect 14525 12567 14583 12573
rect 15077 12607 15135 12613
rect 15077 12573 15089 12607
rect 15123 12604 15135 12607
rect 16917 12607 16975 12613
rect 16917 12604 16929 12607
rect 15123 12576 16929 12604
rect 15123 12573 15135 12576
rect 15077 12567 15135 12573
rect 16917 12573 16929 12576
rect 16963 12573 16975 12607
rect 16917 12567 16975 12573
rect 17469 12607 17527 12613
rect 17469 12573 17481 12607
rect 17515 12604 17527 12607
rect 19309 12607 19367 12613
rect 19309 12604 19321 12607
rect 17515 12576 19321 12604
rect 17515 12573 17527 12576
rect 17469 12567 17527 12573
rect 19309 12573 19321 12576
rect 19355 12573 19367 12607
rect 19309 12567 19367 12573
rect 19861 12607 19919 12613
rect 19861 12573 19873 12607
rect 19907 12573 19919 12607
rect 19861 12567 19919 12573
rect 21057 12607 21115 12613
rect 21057 12573 21069 12607
rect 21103 12604 21115 12607
rect 21606 12604 21612 12616
rect 21103 12576 21612 12604
rect 21103 12573 21115 12576
rect 21057 12567 21115 12573
rect 19876 12468 19904 12567
rect 21606 12564 21612 12576
rect 21664 12564 21670 12616
rect 21701 12471 21759 12477
rect 21701 12468 21713 12471
rect 19876 12440 21713 12468
rect 21701 12437 21713 12440
rect 21747 12437 21759 12471
rect 21701 12431 21759 12437
rect 1904 12378 22236 12400
rect 1904 12326 4446 12378
rect 4498 12326 4510 12378
rect 4562 12326 4574 12378
rect 4626 12326 4638 12378
rect 4690 12326 9774 12378
rect 9826 12326 9838 12378
rect 9890 12326 9902 12378
rect 9954 12326 9966 12378
rect 10018 12326 15102 12378
rect 15154 12326 15166 12378
rect 15218 12326 15230 12378
rect 15282 12326 15294 12378
rect 15346 12326 20430 12378
rect 20482 12326 20494 12378
rect 20546 12326 20558 12378
rect 20610 12326 20622 12378
rect 20674 12326 22236 12378
rect 1904 12304 22236 12326
rect 21606 12224 21612 12276
rect 21664 12264 21670 12276
rect 21701 12267 21759 12273
rect 21701 12264 21713 12267
rect 21664 12236 21713 12264
rect 21664 12224 21670 12236
rect 21701 12233 21713 12236
rect 21747 12233 21759 12267
rect 21701 12227 21759 12233
rect 3117 12131 3175 12137
rect 3117 12097 3129 12131
rect 3163 12128 3175 12131
rect 3850 12128 3856 12140
rect 3163 12100 3856 12128
rect 3163 12097 3175 12100
rect 3117 12091 3175 12097
rect 3850 12088 3856 12100
rect 3908 12088 3914 12140
rect 3761 12063 3819 12069
rect 3761 12029 3773 12063
rect 3807 12060 3819 12063
rect 4313 12063 4371 12069
rect 4313 12060 4325 12063
rect 3807 12032 4325 12060
rect 3807 12029 3819 12032
rect 3761 12023 3819 12029
rect 4313 12029 4325 12032
rect 4359 12029 4371 12063
rect 4313 12023 4371 12029
rect 4957 12063 5015 12069
rect 4957 12029 4969 12063
rect 5003 12060 5015 12063
rect 5509 12063 5567 12069
rect 5509 12060 5521 12063
rect 5003 12032 5521 12060
rect 5003 12029 5015 12032
rect 4957 12023 5015 12029
rect 5509 12029 5521 12032
rect 5555 12029 5567 12063
rect 5509 12023 5567 12029
rect 6153 12063 6211 12069
rect 6153 12029 6165 12063
rect 6199 12060 6211 12063
rect 6705 12063 6763 12069
rect 6705 12060 6717 12063
rect 6199 12032 6717 12060
rect 6199 12029 6211 12032
rect 6153 12023 6211 12029
rect 6705 12029 6717 12032
rect 6751 12029 6763 12063
rect 6705 12023 6763 12029
rect 7349 12063 7407 12069
rect 7349 12029 7361 12063
rect 7395 12060 7407 12063
rect 7901 12063 7959 12069
rect 7901 12060 7913 12063
rect 7395 12032 7913 12060
rect 7395 12029 7407 12032
rect 7349 12023 7407 12029
rect 7901 12029 7913 12032
rect 7947 12029 7959 12063
rect 7901 12023 7959 12029
rect 8545 12063 8603 12069
rect 8545 12029 8557 12063
rect 8591 12060 8603 12063
rect 9097 12063 9155 12069
rect 9097 12060 9109 12063
rect 8591 12032 9109 12060
rect 8591 12029 8603 12032
rect 8545 12023 8603 12029
rect 9097 12029 9109 12032
rect 9143 12029 9155 12063
rect 9097 12023 9155 12029
rect 9741 12063 9799 12069
rect 9741 12029 9753 12063
rect 9787 12060 9799 12063
rect 10293 12063 10351 12069
rect 10293 12060 10305 12063
rect 9787 12032 10305 12060
rect 9787 12029 9799 12032
rect 9741 12023 9799 12029
rect 10293 12029 10305 12032
rect 10339 12029 10351 12063
rect 10293 12023 10351 12029
rect 10937 12063 10995 12069
rect 10937 12029 10949 12063
rect 10983 12060 10995 12063
rect 11489 12063 11547 12069
rect 11489 12060 11501 12063
rect 10983 12032 11501 12060
rect 10983 12029 10995 12032
rect 10937 12023 10995 12029
rect 11489 12029 11501 12032
rect 11535 12029 11547 12063
rect 11489 12023 11547 12029
rect 12133 12063 12191 12069
rect 12133 12029 12145 12063
rect 12179 12060 12191 12063
rect 12685 12063 12743 12069
rect 12685 12060 12697 12063
rect 12179 12032 12697 12060
rect 12179 12029 12191 12032
rect 12133 12023 12191 12029
rect 12685 12029 12697 12032
rect 12731 12029 12743 12063
rect 12685 12023 12743 12029
rect 13329 12063 13387 12069
rect 13329 12029 13341 12063
rect 13375 12060 13387 12063
rect 13881 12063 13939 12069
rect 13881 12060 13893 12063
rect 13375 12032 13893 12060
rect 13375 12029 13387 12032
rect 13329 12023 13387 12029
rect 13881 12029 13893 12032
rect 13927 12029 13939 12063
rect 13881 12023 13939 12029
rect 14525 12063 14583 12069
rect 14525 12029 14537 12063
rect 14571 12060 14583 12063
rect 15077 12063 15135 12069
rect 15077 12060 15089 12063
rect 14571 12032 15089 12060
rect 14571 12029 14583 12032
rect 14525 12023 14583 12029
rect 15077 12029 15089 12032
rect 15123 12029 15135 12063
rect 15077 12023 15135 12029
rect 15721 12063 15779 12069
rect 15721 12029 15733 12063
rect 15767 12060 15779 12063
rect 16273 12063 16331 12069
rect 16273 12060 16285 12063
rect 15767 12032 16285 12060
rect 15767 12029 15779 12032
rect 15721 12023 15779 12029
rect 16273 12029 16285 12032
rect 16319 12029 16331 12063
rect 16273 12023 16331 12029
rect 16917 12063 16975 12069
rect 16917 12029 16929 12063
rect 16963 12060 16975 12063
rect 17469 12063 17527 12069
rect 17469 12060 17481 12063
rect 16963 12032 17481 12060
rect 16963 12029 16975 12032
rect 16917 12023 16975 12029
rect 17469 12029 17481 12032
rect 17515 12029 17527 12063
rect 17469 12023 17527 12029
rect 18113 12063 18171 12069
rect 18113 12029 18125 12063
rect 18159 12060 18171 12063
rect 18665 12063 18723 12069
rect 18665 12060 18677 12063
rect 18159 12032 18677 12060
rect 18159 12029 18171 12032
rect 18113 12023 18171 12029
rect 18665 12029 18677 12032
rect 18711 12029 18723 12063
rect 18665 12023 18723 12029
rect 19309 12063 19367 12069
rect 19309 12029 19321 12063
rect 19355 12060 19367 12063
rect 19861 12063 19919 12069
rect 19861 12060 19873 12063
rect 19355 12032 19873 12060
rect 19355 12029 19367 12032
rect 19309 12023 19367 12029
rect 19861 12029 19873 12032
rect 19907 12029 19919 12063
rect 19861 12023 19919 12029
rect 20505 12063 20563 12069
rect 20505 12029 20517 12063
rect 20551 12060 20563 12063
rect 21057 12063 21115 12069
rect 21057 12060 21069 12063
rect 20551 12032 21069 12060
rect 20551 12029 20563 12032
rect 20505 12023 20563 12029
rect 21057 12029 21069 12032
rect 21103 12029 21115 12063
rect 21057 12023 21115 12029
rect 1904 11834 22236 11856
rect 1904 11782 7110 11834
rect 7162 11782 7174 11834
rect 7226 11782 7238 11834
rect 7290 11782 7302 11834
rect 7354 11782 12438 11834
rect 12490 11782 12502 11834
rect 12554 11782 12566 11834
rect 12618 11782 12630 11834
rect 12682 11782 17766 11834
rect 17818 11782 17830 11834
rect 17882 11782 17894 11834
rect 17946 11782 17958 11834
rect 18010 11782 22236 11834
rect 1904 11760 22236 11782
rect 9112 11624 9324 11652
rect 3761 11587 3819 11593
rect 3761 11553 3773 11587
rect 3807 11584 3819 11587
rect 3850 11584 3856 11596
rect 3807 11556 3856 11584
rect 3807 11553 3819 11556
rect 3761 11547 3819 11553
rect 3850 11544 3856 11556
rect 3908 11544 3914 11596
rect 9112 11593 9140 11624
rect 5509 11587 5567 11593
rect 5509 11553 5521 11587
rect 5555 11584 5567 11587
rect 7349 11587 7407 11593
rect 7349 11584 7361 11587
rect 5555 11556 7361 11584
rect 5555 11553 5567 11556
rect 5509 11547 5567 11553
rect 7349 11553 7361 11556
rect 7395 11553 7407 11587
rect 8545 11587 8603 11593
rect 8545 11584 8557 11587
rect 7349 11547 7407 11553
rect 7824 11556 8557 11584
rect 3117 11519 3175 11525
rect 3117 11485 3129 11519
rect 3163 11485 3175 11519
rect 3117 11479 3175 11485
rect 4313 11519 4371 11525
rect 4313 11485 4325 11519
rect 4359 11516 4371 11519
rect 6153 11519 6211 11525
rect 6153 11516 6165 11519
rect 4359 11488 6165 11516
rect 4359 11485 4371 11488
rect 4313 11479 4371 11485
rect 6153 11485 6165 11488
rect 6199 11485 6211 11519
rect 6153 11479 6211 11485
rect 6705 11519 6763 11525
rect 6705 11485 6717 11519
rect 6751 11516 6763 11519
rect 7824 11516 7852 11556
rect 8545 11553 8557 11556
rect 8591 11553 8603 11587
rect 8545 11547 8603 11553
rect 9097 11587 9155 11593
rect 9097 11553 9109 11587
rect 9143 11584 9155 11587
rect 9296 11584 9324 11624
rect 10937 11587 10995 11593
rect 10937 11584 10949 11587
rect 9143 11556 9177 11584
rect 9296 11556 10949 11584
rect 9143 11553 9155 11556
rect 9097 11547 9155 11553
rect 10937 11553 10949 11556
rect 10983 11553 10995 11587
rect 10937 11547 10995 11553
rect 11489 11587 11547 11593
rect 11489 11553 11501 11587
rect 11535 11584 11547 11587
rect 13329 11587 13387 11593
rect 13329 11584 13341 11587
rect 11535 11556 13341 11584
rect 11535 11553 11547 11556
rect 11489 11547 11547 11553
rect 13329 11553 13341 11556
rect 13375 11553 13387 11587
rect 13329 11547 13387 11553
rect 13881 11587 13939 11593
rect 13881 11553 13893 11587
rect 13927 11584 13939 11587
rect 15721 11587 15779 11593
rect 15721 11584 15733 11587
rect 13927 11556 15733 11584
rect 13927 11553 13939 11556
rect 13881 11547 13939 11553
rect 15721 11553 15733 11556
rect 15767 11553 15779 11587
rect 15721 11547 15779 11553
rect 16273 11587 16331 11593
rect 16273 11553 16285 11587
rect 16319 11584 16331 11587
rect 18113 11587 18171 11593
rect 18113 11584 18125 11587
rect 16319 11556 18125 11584
rect 16319 11553 16331 11556
rect 16273 11547 16331 11553
rect 18113 11553 18125 11556
rect 18159 11553 18171 11587
rect 18113 11547 18171 11553
rect 18665 11587 18723 11593
rect 18665 11553 18677 11587
rect 18711 11584 18723 11587
rect 20505 11587 20563 11593
rect 20505 11584 20517 11587
rect 18711 11556 20517 11584
rect 18711 11553 18723 11556
rect 18665 11547 18723 11553
rect 20505 11553 20517 11556
rect 20551 11553 20563 11587
rect 20505 11547 20563 11553
rect 6751 11488 7852 11516
rect 7901 11519 7959 11525
rect 6751 11485 6763 11488
rect 6705 11479 6763 11485
rect 7901 11485 7913 11519
rect 7947 11516 7959 11519
rect 9741 11519 9799 11525
rect 9741 11516 9753 11519
rect 7947 11488 9753 11516
rect 7947 11485 7959 11488
rect 7901 11479 7959 11485
rect 9741 11485 9753 11488
rect 9787 11485 9799 11519
rect 9741 11479 9799 11485
rect 10293 11519 10351 11525
rect 10293 11485 10305 11519
rect 10339 11516 10351 11519
rect 12133 11519 12191 11525
rect 12133 11516 12145 11519
rect 10339 11488 12145 11516
rect 10339 11485 10351 11488
rect 10293 11479 10351 11485
rect 12133 11485 12145 11488
rect 12179 11485 12191 11519
rect 12133 11479 12191 11485
rect 12685 11519 12743 11525
rect 12685 11485 12697 11519
rect 12731 11516 12743 11519
rect 14525 11519 14583 11525
rect 14525 11516 14537 11519
rect 12731 11488 14537 11516
rect 12731 11485 12743 11488
rect 12685 11479 12743 11485
rect 14525 11485 14537 11488
rect 14571 11485 14583 11519
rect 14525 11479 14583 11485
rect 15077 11519 15135 11525
rect 15077 11485 15089 11519
rect 15123 11516 15135 11519
rect 16917 11519 16975 11525
rect 16917 11516 16929 11519
rect 15123 11488 16929 11516
rect 15123 11485 15135 11488
rect 15077 11479 15135 11485
rect 16917 11485 16929 11488
rect 16963 11485 16975 11519
rect 16917 11479 16975 11485
rect 17469 11519 17527 11525
rect 17469 11485 17481 11519
rect 17515 11516 17527 11519
rect 19309 11519 19367 11525
rect 19309 11516 19321 11519
rect 17515 11488 19321 11516
rect 17515 11485 17527 11488
rect 17469 11479 17527 11485
rect 19309 11485 19321 11488
rect 19355 11485 19367 11519
rect 19309 11479 19367 11485
rect 19861 11519 19919 11525
rect 19861 11485 19873 11519
rect 19907 11485 19919 11519
rect 21054 11516 21060 11528
rect 21015 11488 21060 11516
rect 19861 11479 19919 11485
rect 3132 11448 3160 11479
rect 4957 11451 5015 11457
rect 4957 11448 4969 11451
rect 3132 11420 4969 11448
rect 4957 11417 4969 11420
rect 5003 11417 5015 11451
rect 4957 11411 5015 11417
rect 19876 11380 19904 11479
rect 21054 11476 21060 11488
rect 21112 11476 21118 11528
rect 21701 11383 21759 11389
rect 21701 11380 21713 11383
rect 19876 11352 21713 11380
rect 21701 11349 21713 11352
rect 21747 11349 21759 11383
rect 21701 11343 21759 11349
rect 1904 11290 22236 11312
rect 1904 11238 4446 11290
rect 4498 11238 4510 11290
rect 4562 11238 4574 11290
rect 4626 11238 4638 11290
rect 4690 11238 9774 11290
rect 9826 11238 9838 11290
rect 9890 11238 9902 11290
rect 9954 11238 9966 11290
rect 10018 11238 15102 11290
rect 15154 11238 15166 11290
rect 15218 11238 15230 11290
rect 15282 11238 15294 11290
rect 15346 11238 20430 11290
rect 20482 11238 20494 11290
rect 20546 11238 20558 11290
rect 20610 11238 20622 11290
rect 20674 11238 22236 11290
rect 1904 11216 22236 11238
rect 21054 11136 21060 11188
rect 21112 11176 21118 11188
rect 21701 11179 21759 11185
rect 21701 11176 21713 11179
rect 21112 11148 21713 11176
rect 21112 11136 21118 11148
rect 21701 11145 21713 11148
rect 21747 11145 21759 11179
rect 21701 11139 21759 11145
rect 3117 11043 3175 11049
rect 3117 11009 3129 11043
rect 3163 11040 3175 11043
rect 3850 11040 3856 11052
rect 3163 11012 3856 11040
rect 3163 11009 3175 11012
rect 3117 11003 3175 11009
rect 3850 11000 3856 11012
rect 3908 11000 3914 11052
rect 3761 10975 3819 10981
rect 3761 10941 3773 10975
rect 3807 10972 3819 10975
rect 4313 10975 4371 10981
rect 4313 10972 4325 10975
rect 3807 10944 4325 10972
rect 3807 10941 3819 10944
rect 3761 10935 3819 10941
rect 4313 10941 4325 10944
rect 4359 10941 4371 10975
rect 4313 10935 4371 10941
rect 4957 10975 5015 10981
rect 4957 10941 4969 10975
rect 5003 10972 5015 10975
rect 5509 10975 5567 10981
rect 5509 10972 5521 10975
rect 5003 10944 5521 10972
rect 5003 10941 5015 10944
rect 4957 10935 5015 10941
rect 5509 10941 5521 10944
rect 5555 10941 5567 10975
rect 5509 10935 5567 10941
rect 6153 10975 6211 10981
rect 6153 10941 6165 10975
rect 6199 10972 6211 10975
rect 6705 10975 6763 10981
rect 6705 10972 6717 10975
rect 6199 10944 6717 10972
rect 6199 10941 6211 10944
rect 6153 10935 6211 10941
rect 6705 10941 6717 10944
rect 6751 10941 6763 10975
rect 6705 10935 6763 10941
rect 7349 10975 7407 10981
rect 7349 10941 7361 10975
rect 7395 10972 7407 10975
rect 7901 10975 7959 10981
rect 7901 10972 7913 10975
rect 7395 10944 7913 10972
rect 7395 10941 7407 10944
rect 7349 10935 7407 10941
rect 7901 10941 7913 10944
rect 7947 10941 7959 10975
rect 7901 10935 7959 10941
rect 8545 10975 8603 10981
rect 8545 10941 8557 10975
rect 8591 10972 8603 10975
rect 9097 10975 9155 10981
rect 9097 10972 9109 10975
rect 8591 10944 9109 10972
rect 8591 10941 8603 10944
rect 8545 10935 8603 10941
rect 9097 10941 9109 10944
rect 9143 10941 9155 10975
rect 9097 10935 9155 10941
rect 9741 10975 9799 10981
rect 9741 10941 9753 10975
rect 9787 10972 9799 10975
rect 10293 10975 10351 10981
rect 10293 10972 10305 10975
rect 9787 10944 10305 10972
rect 9787 10941 9799 10944
rect 9741 10935 9799 10941
rect 10293 10941 10305 10944
rect 10339 10941 10351 10975
rect 10293 10935 10351 10941
rect 10937 10975 10995 10981
rect 10937 10941 10949 10975
rect 10983 10972 10995 10975
rect 11489 10975 11547 10981
rect 11489 10972 11501 10975
rect 10983 10944 11501 10972
rect 10983 10941 10995 10944
rect 10937 10935 10995 10941
rect 11489 10941 11501 10944
rect 11535 10941 11547 10975
rect 11489 10935 11547 10941
rect 12133 10975 12191 10981
rect 12133 10941 12145 10975
rect 12179 10972 12191 10975
rect 12685 10975 12743 10981
rect 12685 10972 12697 10975
rect 12179 10944 12697 10972
rect 12179 10941 12191 10944
rect 12133 10935 12191 10941
rect 12685 10941 12697 10944
rect 12731 10941 12743 10975
rect 12685 10935 12743 10941
rect 13329 10975 13387 10981
rect 13329 10941 13341 10975
rect 13375 10972 13387 10975
rect 13881 10975 13939 10981
rect 13881 10972 13893 10975
rect 13375 10944 13893 10972
rect 13375 10941 13387 10944
rect 13329 10935 13387 10941
rect 13881 10941 13893 10944
rect 13927 10941 13939 10975
rect 13881 10935 13939 10941
rect 14525 10975 14583 10981
rect 14525 10941 14537 10975
rect 14571 10972 14583 10975
rect 15077 10975 15135 10981
rect 15077 10972 15089 10975
rect 14571 10944 15089 10972
rect 14571 10941 14583 10944
rect 14525 10935 14583 10941
rect 15077 10941 15089 10944
rect 15123 10941 15135 10975
rect 15077 10935 15135 10941
rect 15721 10975 15779 10981
rect 15721 10941 15733 10975
rect 15767 10972 15779 10975
rect 16273 10975 16331 10981
rect 16273 10972 16285 10975
rect 15767 10944 16285 10972
rect 15767 10941 15779 10944
rect 15721 10935 15779 10941
rect 16273 10941 16285 10944
rect 16319 10941 16331 10975
rect 16273 10935 16331 10941
rect 16917 10975 16975 10981
rect 16917 10941 16929 10975
rect 16963 10972 16975 10975
rect 17469 10975 17527 10981
rect 17469 10972 17481 10975
rect 16963 10944 17481 10972
rect 16963 10941 16975 10944
rect 16917 10935 16975 10941
rect 17469 10941 17481 10944
rect 17515 10941 17527 10975
rect 17469 10935 17527 10941
rect 18113 10975 18171 10981
rect 18113 10941 18125 10975
rect 18159 10972 18171 10975
rect 18665 10975 18723 10981
rect 18665 10972 18677 10975
rect 18159 10944 18677 10972
rect 18159 10941 18171 10944
rect 18113 10935 18171 10941
rect 18665 10941 18677 10944
rect 18711 10941 18723 10975
rect 18665 10935 18723 10941
rect 19309 10975 19367 10981
rect 19309 10941 19321 10975
rect 19355 10972 19367 10975
rect 19861 10975 19919 10981
rect 19861 10972 19873 10975
rect 19355 10944 19873 10972
rect 19355 10941 19367 10944
rect 19309 10935 19367 10941
rect 19861 10941 19873 10944
rect 19907 10941 19919 10975
rect 19861 10935 19919 10941
rect 20505 10975 20563 10981
rect 20505 10941 20517 10975
rect 20551 10972 20563 10975
rect 21057 10975 21115 10981
rect 21057 10972 21069 10975
rect 20551 10944 21069 10972
rect 20551 10941 20563 10944
rect 20505 10935 20563 10941
rect 21057 10941 21069 10944
rect 21103 10941 21115 10975
rect 21057 10935 21115 10941
rect 1904 10746 22236 10768
rect 1904 10694 7110 10746
rect 7162 10694 7174 10746
rect 7226 10694 7238 10746
rect 7290 10694 7302 10746
rect 7354 10694 12438 10746
rect 12490 10694 12502 10746
rect 12554 10694 12566 10746
rect 12618 10694 12630 10746
rect 12682 10694 17766 10746
rect 17818 10694 17830 10746
rect 17882 10694 17894 10746
rect 17946 10694 17958 10746
rect 18010 10694 22236 10746
rect 1904 10672 22236 10694
rect 3761 10635 3819 10641
rect 3761 10601 3773 10635
rect 3807 10632 3819 10635
rect 3850 10632 3856 10644
rect 3807 10604 3856 10632
rect 3807 10601 3819 10604
rect 3761 10595 3819 10601
rect 3850 10592 3856 10604
rect 3908 10592 3914 10644
rect 3117 10499 3175 10505
rect 3117 10465 3129 10499
rect 3163 10496 3175 10499
rect 4957 10499 5015 10505
rect 4957 10496 4969 10499
rect 3163 10468 4969 10496
rect 3163 10465 3175 10468
rect 3117 10459 3175 10465
rect 4957 10465 4969 10468
rect 5003 10465 5015 10499
rect 4957 10459 5015 10465
rect 5509 10499 5567 10505
rect 5509 10465 5521 10499
rect 5555 10496 5567 10499
rect 7349 10499 7407 10505
rect 7349 10496 7361 10499
rect 5555 10468 7361 10496
rect 5555 10465 5567 10468
rect 5509 10459 5567 10465
rect 7349 10465 7361 10468
rect 7395 10465 7407 10499
rect 8545 10499 8603 10505
rect 8545 10496 8557 10499
rect 7349 10459 7407 10465
rect 7824 10468 8557 10496
rect 4313 10431 4371 10437
rect 4313 10397 4325 10431
rect 4359 10428 4371 10431
rect 6153 10431 6211 10437
rect 6153 10428 6165 10431
rect 4359 10400 6165 10428
rect 4359 10397 4371 10400
rect 4313 10391 4371 10397
rect 6153 10397 6165 10400
rect 6199 10397 6211 10431
rect 6153 10391 6211 10397
rect 6705 10431 6763 10437
rect 6705 10397 6717 10431
rect 6751 10428 6763 10431
rect 7824 10428 7852 10468
rect 8545 10465 8557 10468
rect 8591 10465 8603 10499
rect 8545 10459 8603 10465
rect 9097 10499 9155 10505
rect 9097 10465 9109 10499
rect 9143 10496 9155 10499
rect 10937 10499 10995 10505
rect 10937 10496 10949 10499
rect 9143 10468 10949 10496
rect 9143 10465 9155 10468
rect 9097 10459 9155 10465
rect 10937 10465 10949 10468
rect 10983 10465 10995 10499
rect 10937 10459 10995 10465
rect 11489 10499 11547 10505
rect 11489 10465 11501 10499
rect 11535 10496 11547 10499
rect 13329 10499 13387 10505
rect 13329 10496 13341 10499
rect 11535 10468 13341 10496
rect 11535 10465 11547 10468
rect 11489 10459 11547 10465
rect 13329 10465 13341 10468
rect 13375 10465 13387 10499
rect 13329 10459 13387 10465
rect 13881 10499 13939 10505
rect 13881 10465 13893 10499
rect 13927 10496 13939 10499
rect 15721 10499 15779 10505
rect 15721 10496 15733 10499
rect 13927 10468 15733 10496
rect 13927 10465 13939 10468
rect 13881 10459 13939 10465
rect 15721 10465 15733 10468
rect 15767 10465 15779 10499
rect 15721 10459 15779 10465
rect 16273 10499 16331 10505
rect 16273 10465 16285 10499
rect 16319 10496 16331 10499
rect 18113 10499 18171 10505
rect 18113 10496 18125 10499
rect 16319 10468 18125 10496
rect 16319 10465 16331 10468
rect 16273 10459 16331 10465
rect 18113 10465 18125 10468
rect 18159 10465 18171 10499
rect 18113 10459 18171 10465
rect 18665 10499 18723 10505
rect 18665 10465 18677 10499
rect 18711 10496 18723 10499
rect 20505 10499 20563 10505
rect 20505 10496 20517 10499
rect 18711 10468 20517 10496
rect 18711 10465 18723 10468
rect 18665 10459 18723 10465
rect 20505 10465 20517 10468
rect 20551 10465 20563 10499
rect 20505 10459 20563 10465
rect 6751 10400 7852 10428
rect 7901 10431 7959 10437
rect 6751 10397 6763 10400
rect 6705 10391 6763 10397
rect 7901 10397 7913 10431
rect 7947 10428 7959 10431
rect 9741 10431 9799 10437
rect 9741 10428 9753 10431
rect 7947 10400 9753 10428
rect 7947 10397 7959 10400
rect 7901 10391 7959 10397
rect 9741 10397 9753 10400
rect 9787 10397 9799 10431
rect 9741 10391 9799 10397
rect 10293 10431 10351 10437
rect 10293 10397 10305 10431
rect 10339 10428 10351 10431
rect 12133 10431 12191 10437
rect 12133 10428 12145 10431
rect 10339 10400 12145 10428
rect 10339 10397 10351 10400
rect 10293 10391 10351 10397
rect 12133 10397 12145 10400
rect 12179 10397 12191 10431
rect 12133 10391 12191 10397
rect 12685 10431 12743 10437
rect 12685 10397 12697 10431
rect 12731 10428 12743 10431
rect 14525 10431 14583 10437
rect 14525 10428 14537 10431
rect 12731 10400 14537 10428
rect 12731 10397 12743 10400
rect 12685 10391 12743 10397
rect 14525 10397 14537 10400
rect 14571 10397 14583 10431
rect 14525 10391 14583 10397
rect 15077 10431 15135 10437
rect 15077 10397 15089 10431
rect 15123 10428 15135 10431
rect 16917 10431 16975 10437
rect 16917 10428 16929 10431
rect 15123 10400 16929 10428
rect 15123 10397 15135 10400
rect 15077 10391 15135 10397
rect 16917 10397 16929 10400
rect 16963 10397 16975 10431
rect 16917 10391 16975 10397
rect 17469 10431 17527 10437
rect 17469 10397 17481 10431
rect 17515 10428 17527 10431
rect 19309 10431 19367 10437
rect 19309 10428 19321 10431
rect 17515 10400 19321 10428
rect 17515 10397 17527 10400
rect 17469 10391 17527 10397
rect 19309 10397 19321 10400
rect 19355 10397 19367 10431
rect 19309 10391 19367 10397
rect 19861 10431 19919 10437
rect 19861 10397 19873 10431
rect 19907 10397 19919 10431
rect 19861 10391 19919 10397
rect 21057 10431 21115 10437
rect 21057 10397 21069 10431
rect 21103 10428 21115 10431
rect 21606 10428 21612 10440
rect 21103 10400 21612 10428
rect 21103 10397 21115 10400
rect 21057 10391 21115 10397
rect 19876 10292 19904 10391
rect 21606 10388 21612 10400
rect 21664 10388 21670 10440
rect 21701 10295 21759 10301
rect 21701 10292 21713 10295
rect 19876 10264 21713 10292
rect 21701 10261 21713 10264
rect 21747 10261 21759 10295
rect 21701 10255 21759 10261
rect 1904 10202 22236 10224
rect 1904 10150 4446 10202
rect 4498 10150 4510 10202
rect 4562 10150 4574 10202
rect 4626 10150 4638 10202
rect 4690 10150 9774 10202
rect 9826 10150 9838 10202
rect 9890 10150 9902 10202
rect 9954 10150 9966 10202
rect 10018 10150 15102 10202
rect 15154 10150 15166 10202
rect 15218 10150 15230 10202
rect 15282 10150 15294 10202
rect 15346 10150 20430 10202
rect 20482 10150 20494 10202
rect 20546 10150 20558 10202
rect 20610 10150 20622 10202
rect 20674 10150 22236 10202
rect 1904 10128 22236 10150
rect 21606 10048 21612 10100
rect 21664 10088 21670 10100
rect 21701 10091 21759 10097
rect 21701 10088 21713 10091
rect 21664 10060 21713 10088
rect 21664 10048 21670 10060
rect 21701 10057 21713 10060
rect 21747 10057 21759 10091
rect 21701 10051 21759 10057
rect 2286 9912 2292 9964
rect 2344 9952 2350 9964
rect 3117 9955 3175 9961
rect 3117 9952 3129 9955
rect 2344 9924 3129 9952
rect 2344 9912 2350 9924
rect 3117 9921 3129 9924
rect 3163 9921 3175 9955
rect 3117 9915 3175 9921
rect 3761 9887 3819 9893
rect 3761 9853 3773 9887
rect 3807 9884 3819 9887
rect 4313 9887 4371 9893
rect 4313 9884 4325 9887
rect 3807 9856 4325 9884
rect 3807 9853 3819 9856
rect 3761 9847 3819 9853
rect 4313 9853 4325 9856
rect 4359 9853 4371 9887
rect 4313 9847 4371 9853
rect 4957 9887 5015 9893
rect 4957 9853 4969 9887
rect 5003 9884 5015 9887
rect 5509 9887 5567 9893
rect 5509 9884 5521 9887
rect 5003 9856 5521 9884
rect 5003 9853 5015 9856
rect 4957 9847 5015 9853
rect 5509 9853 5521 9856
rect 5555 9853 5567 9887
rect 5509 9847 5567 9853
rect 6153 9887 6211 9893
rect 6153 9853 6165 9887
rect 6199 9884 6211 9887
rect 6705 9887 6763 9893
rect 6705 9884 6717 9887
rect 6199 9856 6717 9884
rect 6199 9853 6211 9856
rect 6153 9847 6211 9853
rect 6705 9853 6717 9856
rect 6751 9853 6763 9887
rect 6705 9847 6763 9853
rect 7349 9887 7407 9893
rect 7349 9853 7361 9887
rect 7395 9884 7407 9887
rect 7901 9887 7959 9893
rect 7901 9884 7913 9887
rect 7395 9856 7913 9884
rect 7395 9853 7407 9856
rect 7349 9847 7407 9853
rect 7901 9853 7913 9856
rect 7947 9853 7959 9887
rect 7901 9847 7959 9853
rect 8545 9887 8603 9893
rect 8545 9853 8557 9887
rect 8591 9884 8603 9887
rect 9097 9887 9155 9893
rect 9097 9884 9109 9887
rect 8591 9856 9109 9884
rect 8591 9853 8603 9856
rect 8545 9847 8603 9853
rect 9097 9853 9109 9856
rect 9143 9853 9155 9887
rect 9097 9847 9155 9853
rect 9741 9887 9799 9893
rect 9741 9853 9753 9887
rect 9787 9884 9799 9887
rect 10293 9887 10351 9893
rect 10293 9884 10305 9887
rect 9787 9856 10305 9884
rect 9787 9853 9799 9856
rect 9741 9847 9799 9853
rect 10293 9853 10305 9856
rect 10339 9853 10351 9887
rect 10293 9847 10351 9853
rect 10937 9887 10995 9893
rect 10937 9853 10949 9887
rect 10983 9884 10995 9887
rect 11489 9887 11547 9893
rect 11489 9884 11501 9887
rect 10983 9856 11501 9884
rect 10983 9853 10995 9856
rect 10937 9847 10995 9853
rect 11489 9853 11501 9856
rect 11535 9853 11547 9887
rect 11489 9847 11547 9853
rect 12133 9887 12191 9893
rect 12133 9853 12145 9887
rect 12179 9884 12191 9887
rect 12685 9887 12743 9893
rect 12685 9884 12697 9887
rect 12179 9856 12697 9884
rect 12179 9853 12191 9856
rect 12133 9847 12191 9853
rect 12685 9853 12697 9856
rect 12731 9853 12743 9887
rect 12685 9847 12743 9853
rect 13329 9887 13387 9893
rect 13329 9853 13341 9887
rect 13375 9884 13387 9887
rect 13881 9887 13939 9893
rect 13881 9884 13893 9887
rect 13375 9856 13893 9884
rect 13375 9853 13387 9856
rect 13329 9847 13387 9853
rect 13881 9853 13893 9856
rect 13927 9853 13939 9887
rect 13881 9847 13939 9853
rect 14525 9887 14583 9893
rect 14525 9853 14537 9887
rect 14571 9884 14583 9887
rect 15077 9887 15135 9893
rect 15077 9884 15089 9887
rect 14571 9856 15089 9884
rect 14571 9853 14583 9856
rect 14525 9847 14583 9853
rect 15077 9853 15089 9856
rect 15123 9853 15135 9887
rect 15077 9847 15135 9853
rect 15721 9887 15779 9893
rect 15721 9853 15733 9887
rect 15767 9884 15779 9887
rect 16273 9887 16331 9893
rect 16273 9884 16285 9887
rect 15767 9856 16285 9884
rect 15767 9853 15779 9856
rect 15721 9847 15779 9853
rect 16273 9853 16285 9856
rect 16319 9853 16331 9887
rect 16273 9847 16331 9853
rect 16917 9887 16975 9893
rect 16917 9853 16929 9887
rect 16963 9884 16975 9887
rect 17469 9887 17527 9893
rect 17469 9884 17481 9887
rect 16963 9856 17481 9884
rect 16963 9853 16975 9856
rect 16917 9847 16975 9853
rect 17469 9853 17481 9856
rect 17515 9853 17527 9887
rect 17469 9847 17527 9853
rect 18113 9887 18171 9893
rect 18113 9853 18125 9887
rect 18159 9884 18171 9887
rect 18665 9887 18723 9893
rect 18665 9884 18677 9887
rect 18159 9856 18677 9884
rect 18159 9853 18171 9856
rect 18113 9847 18171 9853
rect 18665 9853 18677 9856
rect 18711 9853 18723 9887
rect 18665 9847 18723 9853
rect 19309 9887 19367 9893
rect 19309 9853 19321 9887
rect 19355 9884 19367 9887
rect 19861 9887 19919 9893
rect 19861 9884 19873 9887
rect 19355 9856 19873 9884
rect 19355 9853 19367 9856
rect 19309 9847 19367 9853
rect 19861 9853 19873 9856
rect 19907 9853 19919 9887
rect 19861 9847 19919 9853
rect 20505 9887 20563 9893
rect 20505 9853 20517 9887
rect 20551 9884 20563 9887
rect 21057 9887 21115 9893
rect 21057 9884 21069 9887
rect 20551 9856 21069 9884
rect 20551 9853 20563 9856
rect 20505 9847 20563 9853
rect 21057 9853 21069 9856
rect 21103 9853 21115 9887
rect 21057 9847 21115 9853
rect 1904 9658 22236 9680
rect 1904 9606 7110 9658
rect 7162 9606 7174 9658
rect 7226 9606 7238 9658
rect 7290 9606 7302 9658
rect 7354 9606 12438 9658
rect 12490 9606 12502 9658
rect 12554 9606 12566 9658
rect 12618 9606 12630 9658
rect 12682 9606 17766 9658
rect 17818 9606 17830 9658
rect 17882 9606 17894 9658
rect 17946 9606 17958 9658
rect 18010 9606 22236 9658
rect 1904 9584 22236 9606
rect 2470 9408 2476 9420
rect 2431 9380 2476 9408
rect 2470 9368 2476 9380
rect 2528 9368 2534 9420
rect 3117 9411 3175 9417
rect 3117 9377 3129 9411
rect 3163 9408 3175 9411
rect 4957 9411 5015 9417
rect 4957 9408 4969 9411
rect 3163 9380 4969 9408
rect 3163 9377 3175 9380
rect 3117 9371 3175 9377
rect 4957 9377 4969 9380
rect 5003 9377 5015 9411
rect 4957 9371 5015 9377
rect 5509 9411 5567 9417
rect 5509 9377 5521 9411
rect 5555 9408 5567 9411
rect 7349 9411 7407 9417
rect 7349 9408 7361 9411
rect 5555 9380 7361 9408
rect 5555 9377 5567 9380
rect 5509 9371 5567 9377
rect 7349 9377 7361 9380
rect 7395 9377 7407 9411
rect 8545 9411 8603 9417
rect 8545 9408 8557 9411
rect 7349 9371 7407 9377
rect 7456 9380 8557 9408
rect 2286 9300 2292 9352
rect 2344 9300 2350 9352
rect 4313 9343 4371 9349
rect 4313 9309 4325 9343
rect 4359 9340 4371 9343
rect 6153 9343 6211 9349
rect 6153 9340 6165 9343
rect 4359 9312 6165 9340
rect 4359 9309 4371 9312
rect 4313 9303 4371 9309
rect 6153 9309 6165 9312
rect 6199 9309 6211 9343
rect 6153 9303 6211 9309
rect 6705 9343 6763 9349
rect 6705 9309 6717 9343
rect 6751 9340 6763 9343
rect 7456 9340 7484 9380
rect 8545 9377 8557 9380
rect 8591 9377 8603 9411
rect 8545 9371 8603 9377
rect 9097 9411 9155 9417
rect 9097 9377 9109 9411
rect 9143 9408 9155 9411
rect 10937 9411 10995 9417
rect 10937 9408 10949 9411
rect 9143 9380 10949 9408
rect 9143 9377 9155 9380
rect 9097 9371 9155 9377
rect 10937 9377 10949 9380
rect 10983 9377 10995 9411
rect 10937 9371 10995 9377
rect 11489 9411 11547 9417
rect 11489 9377 11501 9411
rect 11535 9408 11547 9411
rect 13329 9411 13387 9417
rect 13329 9408 13341 9411
rect 11535 9380 13341 9408
rect 11535 9377 11547 9380
rect 11489 9371 11547 9377
rect 13329 9377 13341 9380
rect 13375 9377 13387 9411
rect 13329 9371 13387 9377
rect 13881 9411 13939 9417
rect 13881 9377 13893 9411
rect 13927 9408 13939 9411
rect 15721 9411 15779 9417
rect 15721 9408 15733 9411
rect 13927 9380 15733 9408
rect 13927 9377 13939 9380
rect 13881 9371 13939 9377
rect 15721 9377 15733 9380
rect 15767 9377 15779 9411
rect 15721 9371 15779 9377
rect 16273 9411 16331 9417
rect 16273 9377 16285 9411
rect 16319 9408 16331 9411
rect 18113 9411 18171 9417
rect 18113 9408 18125 9411
rect 16319 9380 18125 9408
rect 16319 9377 16331 9380
rect 16273 9371 16331 9377
rect 18113 9377 18125 9380
rect 18159 9377 18171 9411
rect 18113 9371 18171 9377
rect 18665 9411 18723 9417
rect 18665 9377 18677 9411
rect 18711 9408 18723 9411
rect 20505 9411 20563 9417
rect 20505 9408 20517 9411
rect 18711 9380 20517 9408
rect 18711 9377 18723 9380
rect 18665 9371 18723 9377
rect 20505 9377 20517 9380
rect 20551 9377 20563 9411
rect 20505 9371 20563 9377
rect 6751 9312 7484 9340
rect 7901 9343 7959 9349
rect 6751 9309 6763 9312
rect 6705 9303 6763 9309
rect 7901 9309 7913 9343
rect 7947 9340 7959 9343
rect 9741 9343 9799 9349
rect 9741 9340 9753 9343
rect 7947 9312 9753 9340
rect 7947 9309 7959 9312
rect 7901 9303 7959 9309
rect 9741 9309 9753 9312
rect 9787 9309 9799 9343
rect 9741 9303 9799 9309
rect 10293 9343 10351 9349
rect 10293 9309 10305 9343
rect 10339 9340 10351 9343
rect 12133 9343 12191 9349
rect 12133 9340 12145 9343
rect 10339 9312 12145 9340
rect 10339 9309 10351 9312
rect 10293 9303 10351 9309
rect 12133 9309 12145 9312
rect 12179 9309 12191 9343
rect 12133 9303 12191 9309
rect 12685 9343 12743 9349
rect 12685 9309 12697 9343
rect 12731 9340 12743 9343
rect 14525 9343 14583 9349
rect 14525 9340 14537 9343
rect 12731 9312 14537 9340
rect 12731 9309 12743 9312
rect 12685 9303 12743 9309
rect 14525 9309 14537 9312
rect 14571 9309 14583 9343
rect 14525 9303 14583 9309
rect 15077 9343 15135 9349
rect 15077 9309 15089 9343
rect 15123 9340 15135 9343
rect 16917 9343 16975 9349
rect 16917 9340 16929 9343
rect 15123 9312 16929 9340
rect 15123 9309 15135 9312
rect 15077 9303 15135 9309
rect 16917 9309 16929 9312
rect 16963 9309 16975 9343
rect 16917 9303 16975 9309
rect 17469 9343 17527 9349
rect 17469 9309 17481 9343
rect 17515 9340 17527 9343
rect 19309 9343 19367 9349
rect 19309 9340 19321 9343
rect 17515 9312 19321 9340
rect 17515 9309 17527 9312
rect 17469 9303 17527 9309
rect 19309 9309 19321 9312
rect 19355 9309 19367 9343
rect 19309 9303 19367 9309
rect 19861 9343 19919 9349
rect 19861 9309 19873 9343
rect 19907 9309 19919 9343
rect 21054 9340 21060 9352
rect 21015 9312 21060 9340
rect 19861 9303 19919 9309
rect 2304 9272 2332 9300
rect 1936 9244 2332 9272
rect 2381 9275 2439 9281
rect 1936 9213 1964 9244
rect 2381 9241 2393 9275
rect 2427 9272 2439 9275
rect 3761 9275 3819 9281
rect 3761 9272 3773 9275
rect 2427 9244 3773 9272
rect 2427 9241 2439 9244
rect 2381 9235 2439 9241
rect 3761 9241 3773 9244
rect 3807 9241 3819 9275
rect 3761 9235 3819 9241
rect 1921 9207 1979 9213
rect 1921 9173 1933 9207
rect 1967 9173 1979 9207
rect 1921 9167 1979 9173
rect 2286 9164 2292 9216
rect 2344 9204 2350 9216
rect 19876 9204 19904 9303
rect 21054 9300 21060 9312
rect 21112 9300 21118 9352
rect 21701 9207 21759 9213
rect 21701 9204 21713 9207
rect 2344 9176 2389 9204
rect 19876 9176 21713 9204
rect 2344 9164 2350 9176
rect 21701 9173 21713 9176
rect 21747 9173 21759 9207
rect 21701 9167 21759 9173
rect 1904 9114 22236 9136
rect 1904 9062 4446 9114
rect 4498 9062 4510 9114
rect 4562 9062 4574 9114
rect 4626 9062 4638 9114
rect 4690 9062 9774 9114
rect 9826 9062 9838 9114
rect 9890 9062 9902 9114
rect 9954 9062 9966 9114
rect 10018 9062 15102 9114
rect 15154 9062 15166 9114
rect 15218 9062 15230 9114
rect 15282 9062 15294 9114
rect 15346 9062 20430 9114
rect 20482 9062 20494 9114
rect 20546 9062 20558 9114
rect 20610 9062 20622 9114
rect 20674 9062 22236 9114
rect 1904 9040 22236 9062
rect 21054 8960 21060 9012
rect 21112 9000 21118 9012
rect 21701 9003 21759 9009
rect 21701 9000 21713 9003
rect 21112 8972 21713 9000
rect 21112 8960 21118 8972
rect 21701 8969 21713 8972
rect 21747 8969 21759 9003
rect 21701 8963 21759 8969
rect 3117 8867 3175 8873
rect 3117 8833 3129 8867
rect 3163 8864 3175 8867
rect 3850 8864 3856 8876
rect 3163 8836 3856 8864
rect 3163 8833 3175 8836
rect 3117 8827 3175 8833
rect 3850 8824 3856 8836
rect 3908 8824 3914 8876
rect 3761 8799 3819 8805
rect 3761 8765 3773 8799
rect 3807 8796 3819 8799
rect 4313 8799 4371 8805
rect 4313 8796 4325 8799
rect 3807 8768 4325 8796
rect 3807 8765 3819 8768
rect 3761 8759 3819 8765
rect 4313 8765 4325 8768
rect 4359 8765 4371 8799
rect 4313 8759 4371 8765
rect 4957 8799 5015 8805
rect 4957 8765 4969 8799
rect 5003 8796 5015 8799
rect 5509 8799 5567 8805
rect 5509 8796 5521 8799
rect 5003 8768 5521 8796
rect 5003 8765 5015 8768
rect 4957 8759 5015 8765
rect 5509 8765 5521 8768
rect 5555 8765 5567 8799
rect 5509 8759 5567 8765
rect 6153 8799 6211 8805
rect 6153 8765 6165 8799
rect 6199 8796 6211 8799
rect 6705 8799 6763 8805
rect 6705 8796 6717 8799
rect 6199 8768 6717 8796
rect 6199 8765 6211 8768
rect 6153 8759 6211 8765
rect 6705 8765 6717 8768
rect 6751 8765 6763 8799
rect 6705 8759 6763 8765
rect 7349 8799 7407 8805
rect 7349 8765 7361 8799
rect 7395 8796 7407 8799
rect 7901 8799 7959 8805
rect 7901 8796 7913 8799
rect 7395 8768 7913 8796
rect 7395 8765 7407 8768
rect 7349 8759 7407 8765
rect 7901 8765 7913 8768
rect 7947 8765 7959 8799
rect 7901 8759 7959 8765
rect 8545 8799 8603 8805
rect 8545 8765 8557 8799
rect 8591 8796 8603 8799
rect 9097 8799 9155 8805
rect 9097 8796 9109 8799
rect 8591 8768 9109 8796
rect 8591 8765 8603 8768
rect 8545 8759 8603 8765
rect 9097 8765 9109 8768
rect 9143 8765 9155 8799
rect 9097 8759 9155 8765
rect 9741 8799 9799 8805
rect 9741 8765 9753 8799
rect 9787 8796 9799 8799
rect 10293 8799 10351 8805
rect 10293 8796 10305 8799
rect 9787 8768 10305 8796
rect 9787 8765 9799 8768
rect 9741 8759 9799 8765
rect 10293 8765 10305 8768
rect 10339 8765 10351 8799
rect 10293 8759 10351 8765
rect 10937 8799 10995 8805
rect 10937 8765 10949 8799
rect 10983 8796 10995 8799
rect 11489 8799 11547 8805
rect 11489 8796 11501 8799
rect 10983 8768 11501 8796
rect 10983 8765 10995 8768
rect 10937 8759 10995 8765
rect 11489 8765 11501 8768
rect 11535 8765 11547 8799
rect 11489 8759 11547 8765
rect 12133 8799 12191 8805
rect 12133 8765 12145 8799
rect 12179 8796 12191 8799
rect 12685 8799 12743 8805
rect 12685 8796 12697 8799
rect 12179 8768 12697 8796
rect 12179 8765 12191 8768
rect 12133 8759 12191 8765
rect 12685 8765 12697 8768
rect 12731 8765 12743 8799
rect 12685 8759 12743 8765
rect 13329 8799 13387 8805
rect 13329 8765 13341 8799
rect 13375 8796 13387 8799
rect 13881 8799 13939 8805
rect 13881 8796 13893 8799
rect 13375 8768 13893 8796
rect 13375 8765 13387 8768
rect 13329 8759 13387 8765
rect 13881 8765 13893 8768
rect 13927 8765 13939 8799
rect 13881 8759 13939 8765
rect 14525 8799 14583 8805
rect 14525 8765 14537 8799
rect 14571 8796 14583 8799
rect 15077 8799 15135 8805
rect 15077 8796 15089 8799
rect 14571 8768 15089 8796
rect 14571 8765 14583 8768
rect 14525 8759 14583 8765
rect 15077 8765 15089 8768
rect 15123 8765 15135 8799
rect 15077 8759 15135 8765
rect 15721 8799 15779 8805
rect 15721 8765 15733 8799
rect 15767 8796 15779 8799
rect 16273 8799 16331 8805
rect 16273 8796 16285 8799
rect 15767 8768 16285 8796
rect 15767 8765 15779 8768
rect 15721 8759 15779 8765
rect 16273 8765 16285 8768
rect 16319 8765 16331 8799
rect 16273 8759 16331 8765
rect 16917 8799 16975 8805
rect 16917 8765 16929 8799
rect 16963 8796 16975 8799
rect 17469 8799 17527 8805
rect 17469 8796 17481 8799
rect 16963 8768 17481 8796
rect 16963 8765 16975 8768
rect 16917 8759 16975 8765
rect 17469 8765 17481 8768
rect 17515 8765 17527 8799
rect 17469 8759 17527 8765
rect 18113 8799 18171 8805
rect 18113 8765 18125 8799
rect 18159 8796 18171 8799
rect 18665 8799 18723 8805
rect 18665 8796 18677 8799
rect 18159 8768 18677 8796
rect 18159 8765 18171 8768
rect 18113 8759 18171 8765
rect 18665 8765 18677 8768
rect 18711 8765 18723 8799
rect 18665 8759 18723 8765
rect 19309 8799 19367 8805
rect 19309 8765 19321 8799
rect 19355 8796 19367 8799
rect 19861 8799 19919 8805
rect 19861 8796 19873 8799
rect 19355 8768 19873 8796
rect 19355 8765 19367 8768
rect 19309 8759 19367 8765
rect 19861 8765 19873 8768
rect 19907 8765 19919 8799
rect 19861 8759 19919 8765
rect 20505 8799 20563 8805
rect 20505 8765 20517 8799
rect 20551 8796 20563 8799
rect 21057 8799 21115 8805
rect 21057 8796 21069 8799
rect 20551 8768 21069 8796
rect 20551 8765 20563 8768
rect 20505 8759 20563 8765
rect 21057 8765 21069 8768
rect 21103 8765 21115 8799
rect 21057 8759 21115 8765
rect 1904 8570 22236 8592
rect 1904 8518 7110 8570
rect 7162 8518 7174 8570
rect 7226 8518 7238 8570
rect 7290 8518 7302 8570
rect 7354 8518 12438 8570
rect 12490 8518 12502 8570
rect 12554 8518 12566 8570
rect 12618 8518 12630 8570
rect 12682 8518 17766 8570
rect 17818 8518 17830 8570
rect 17882 8518 17894 8570
rect 17946 8518 17958 8570
rect 18010 8518 22236 8570
rect 1904 8496 22236 8518
rect 3761 8459 3819 8465
rect 3761 8425 3773 8459
rect 3807 8456 3819 8459
rect 3850 8456 3856 8468
rect 3807 8428 3856 8456
rect 3807 8425 3819 8428
rect 3761 8419 3819 8425
rect 3850 8416 3856 8428
rect 3908 8416 3914 8468
rect 3117 8323 3175 8329
rect 3117 8289 3129 8323
rect 3163 8320 3175 8323
rect 4957 8323 5015 8329
rect 4957 8320 4969 8323
rect 3163 8292 4969 8320
rect 3163 8289 3175 8292
rect 3117 8283 3175 8289
rect 4957 8289 4969 8292
rect 5003 8289 5015 8323
rect 4957 8283 5015 8289
rect 5509 8323 5567 8329
rect 5509 8289 5521 8323
rect 5555 8320 5567 8323
rect 7349 8323 7407 8329
rect 7349 8320 7361 8323
rect 5555 8292 7361 8320
rect 5555 8289 5567 8292
rect 5509 8283 5567 8289
rect 7349 8289 7361 8292
rect 7395 8289 7407 8323
rect 8545 8323 8603 8329
rect 8545 8320 8557 8323
rect 7349 8283 7407 8289
rect 7824 8292 8557 8320
rect 4313 8255 4371 8261
rect 4313 8221 4325 8255
rect 4359 8252 4371 8255
rect 6153 8255 6211 8261
rect 6153 8252 6165 8255
rect 4359 8224 6165 8252
rect 4359 8221 4371 8224
rect 4313 8215 4371 8221
rect 6153 8221 6165 8224
rect 6199 8221 6211 8255
rect 6153 8215 6211 8221
rect 6705 8255 6763 8261
rect 6705 8221 6717 8255
rect 6751 8252 6763 8255
rect 7824 8252 7852 8292
rect 8545 8289 8557 8292
rect 8591 8289 8603 8323
rect 8545 8283 8603 8289
rect 9097 8323 9155 8329
rect 9097 8289 9109 8323
rect 9143 8320 9155 8323
rect 10937 8323 10995 8329
rect 10937 8320 10949 8323
rect 9143 8292 10949 8320
rect 9143 8289 9155 8292
rect 9097 8283 9155 8289
rect 10937 8289 10949 8292
rect 10983 8289 10995 8323
rect 10937 8283 10995 8289
rect 11489 8323 11547 8329
rect 11489 8289 11501 8323
rect 11535 8320 11547 8323
rect 13329 8323 13387 8329
rect 13329 8320 13341 8323
rect 11535 8292 13341 8320
rect 11535 8289 11547 8292
rect 11489 8283 11547 8289
rect 13329 8289 13341 8292
rect 13375 8289 13387 8323
rect 13329 8283 13387 8289
rect 13881 8323 13939 8329
rect 13881 8289 13893 8323
rect 13927 8320 13939 8323
rect 15721 8323 15779 8329
rect 15721 8320 15733 8323
rect 13927 8292 15733 8320
rect 13927 8289 13939 8292
rect 13881 8283 13939 8289
rect 15721 8289 15733 8292
rect 15767 8289 15779 8323
rect 15721 8283 15779 8289
rect 16273 8323 16331 8329
rect 16273 8289 16285 8323
rect 16319 8320 16331 8323
rect 18113 8323 18171 8329
rect 18113 8320 18125 8323
rect 16319 8292 18125 8320
rect 16319 8289 16331 8292
rect 16273 8283 16331 8289
rect 18113 8289 18125 8292
rect 18159 8289 18171 8323
rect 18113 8283 18171 8289
rect 18665 8323 18723 8329
rect 18665 8289 18677 8323
rect 18711 8320 18723 8323
rect 20505 8323 20563 8329
rect 20505 8320 20517 8323
rect 18711 8292 20517 8320
rect 18711 8289 18723 8292
rect 18665 8283 18723 8289
rect 20505 8289 20517 8292
rect 20551 8289 20563 8323
rect 20505 8283 20563 8289
rect 6751 8224 7852 8252
rect 7901 8255 7959 8261
rect 6751 8221 6763 8224
rect 6705 8215 6763 8221
rect 7901 8221 7913 8255
rect 7947 8252 7959 8255
rect 9741 8255 9799 8261
rect 9741 8252 9753 8255
rect 7947 8224 9753 8252
rect 7947 8221 7959 8224
rect 7901 8215 7959 8221
rect 9741 8221 9753 8224
rect 9787 8221 9799 8255
rect 9741 8215 9799 8221
rect 10293 8255 10351 8261
rect 10293 8221 10305 8255
rect 10339 8252 10351 8255
rect 12133 8255 12191 8261
rect 12133 8252 12145 8255
rect 10339 8224 12145 8252
rect 10339 8221 10351 8224
rect 10293 8215 10351 8221
rect 12133 8221 12145 8224
rect 12179 8221 12191 8255
rect 12133 8215 12191 8221
rect 12685 8255 12743 8261
rect 12685 8221 12697 8255
rect 12731 8252 12743 8255
rect 14525 8255 14583 8261
rect 14525 8252 14537 8255
rect 12731 8224 14537 8252
rect 12731 8221 12743 8224
rect 12685 8215 12743 8221
rect 14525 8221 14537 8224
rect 14571 8221 14583 8255
rect 14525 8215 14583 8221
rect 15077 8255 15135 8261
rect 15077 8221 15089 8255
rect 15123 8252 15135 8255
rect 16917 8255 16975 8261
rect 16917 8252 16929 8255
rect 15123 8224 16929 8252
rect 15123 8221 15135 8224
rect 15077 8215 15135 8221
rect 16917 8221 16929 8224
rect 16963 8221 16975 8255
rect 16917 8215 16975 8221
rect 17469 8255 17527 8261
rect 17469 8221 17481 8255
rect 17515 8252 17527 8255
rect 19309 8255 19367 8261
rect 19309 8252 19321 8255
rect 17515 8224 19321 8252
rect 17515 8221 17527 8224
rect 17469 8215 17527 8221
rect 19309 8221 19321 8224
rect 19355 8221 19367 8255
rect 19309 8215 19367 8221
rect 19861 8255 19919 8261
rect 19861 8221 19873 8255
rect 19907 8221 19919 8255
rect 19861 8215 19919 8221
rect 21057 8255 21115 8261
rect 21057 8221 21069 8255
rect 21103 8252 21115 8255
rect 21606 8252 21612 8264
rect 21103 8224 21612 8252
rect 21103 8221 21115 8224
rect 21057 8215 21115 8221
rect 19876 8116 19904 8215
rect 21606 8212 21612 8224
rect 21664 8212 21670 8264
rect 21701 8119 21759 8125
rect 21701 8116 21713 8119
rect 19876 8088 21713 8116
rect 21701 8085 21713 8088
rect 21747 8085 21759 8119
rect 21701 8079 21759 8085
rect 1904 8026 22236 8048
rect 1904 7974 4446 8026
rect 4498 7974 4510 8026
rect 4562 7974 4574 8026
rect 4626 7974 4638 8026
rect 4690 7974 9774 8026
rect 9826 7974 9838 8026
rect 9890 7974 9902 8026
rect 9954 7974 9966 8026
rect 10018 7974 15102 8026
rect 15154 7974 15166 8026
rect 15218 7974 15230 8026
rect 15282 7974 15294 8026
rect 15346 7974 20430 8026
rect 20482 7974 20494 8026
rect 20546 7974 20558 8026
rect 20610 7974 20622 8026
rect 20674 7974 22236 8026
rect 1904 7952 22236 7974
rect 21606 7872 21612 7924
rect 21664 7912 21670 7924
rect 21701 7915 21759 7921
rect 21701 7912 21713 7915
rect 21664 7884 21713 7912
rect 21664 7872 21670 7884
rect 21701 7881 21713 7884
rect 21747 7881 21759 7915
rect 21701 7875 21759 7881
rect 3117 7779 3175 7785
rect 3117 7745 3129 7779
rect 3163 7776 3175 7779
rect 3850 7776 3856 7788
rect 3163 7748 3856 7776
rect 3163 7745 3175 7748
rect 3117 7739 3175 7745
rect 3850 7736 3856 7748
rect 3908 7736 3914 7788
rect 3761 7711 3819 7717
rect 3761 7677 3773 7711
rect 3807 7708 3819 7711
rect 4313 7711 4371 7717
rect 4313 7708 4325 7711
rect 3807 7680 4325 7708
rect 3807 7677 3819 7680
rect 3761 7671 3819 7677
rect 4313 7677 4325 7680
rect 4359 7677 4371 7711
rect 4313 7671 4371 7677
rect 4957 7711 5015 7717
rect 4957 7677 4969 7711
rect 5003 7708 5015 7711
rect 5509 7711 5567 7717
rect 5509 7708 5521 7711
rect 5003 7680 5521 7708
rect 5003 7677 5015 7680
rect 4957 7671 5015 7677
rect 5509 7677 5521 7680
rect 5555 7677 5567 7711
rect 5509 7671 5567 7677
rect 6153 7711 6211 7717
rect 6153 7677 6165 7711
rect 6199 7708 6211 7711
rect 6705 7711 6763 7717
rect 6705 7708 6717 7711
rect 6199 7680 6717 7708
rect 6199 7677 6211 7680
rect 6153 7671 6211 7677
rect 6705 7677 6717 7680
rect 6751 7677 6763 7711
rect 6705 7671 6763 7677
rect 7349 7711 7407 7717
rect 7349 7677 7361 7711
rect 7395 7708 7407 7711
rect 7901 7711 7959 7717
rect 7901 7708 7913 7711
rect 7395 7680 7913 7708
rect 7395 7677 7407 7680
rect 7349 7671 7407 7677
rect 7901 7677 7913 7680
rect 7947 7677 7959 7711
rect 7901 7671 7959 7677
rect 8545 7711 8603 7717
rect 8545 7677 8557 7711
rect 8591 7708 8603 7711
rect 9097 7711 9155 7717
rect 9097 7708 9109 7711
rect 8591 7680 9109 7708
rect 8591 7677 8603 7680
rect 8545 7671 8603 7677
rect 9097 7677 9109 7680
rect 9143 7677 9155 7711
rect 9097 7671 9155 7677
rect 9741 7711 9799 7717
rect 9741 7677 9753 7711
rect 9787 7708 9799 7711
rect 10293 7711 10351 7717
rect 10293 7708 10305 7711
rect 9787 7680 10305 7708
rect 9787 7677 9799 7680
rect 9741 7671 9799 7677
rect 10293 7677 10305 7680
rect 10339 7677 10351 7711
rect 10293 7671 10351 7677
rect 10937 7711 10995 7717
rect 10937 7677 10949 7711
rect 10983 7708 10995 7711
rect 11489 7711 11547 7717
rect 11489 7708 11501 7711
rect 10983 7680 11501 7708
rect 10983 7677 10995 7680
rect 10937 7671 10995 7677
rect 11489 7677 11501 7680
rect 11535 7677 11547 7711
rect 11489 7671 11547 7677
rect 12133 7711 12191 7717
rect 12133 7677 12145 7711
rect 12179 7708 12191 7711
rect 12685 7711 12743 7717
rect 12685 7708 12697 7711
rect 12179 7680 12697 7708
rect 12179 7677 12191 7680
rect 12133 7671 12191 7677
rect 12685 7677 12697 7680
rect 12731 7677 12743 7711
rect 12685 7671 12743 7677
rect 13329 7711 13387 7717
rect 13329 7677 13341 7711
rect 13375 7708 13387 7711
rect 13881 7711 13939 7717
rect 13881 7708 13893 7711
rect 13375 7680 13893 7708
rect 13375 7677 13387 7680
rect 13329 7671 13387 7677
rect 13881 7677 13893 7680
rect 13927 7677 13939 7711
rect 13881 7671 13939 7677
rect 14525 7711 14583 7717
rect 14525 7677 14537 7711
rect 14571 7708 14583 7711
rect 15077 7711 15135 7717
rect 15077 7708 15089 7711
rect 14571 7680 15089 7708
rect 14571 7677 14583 7680
rect 14525 7671 14583 7677
rect 15077 7677 15089 7680
rect 15123 7677 15135 7711
rect 15077 7671 15135 7677
rect 15721 7711 15779 7717
rect 15721 7677 15733 7711
rect 15767 7708 15779 7711
rect 16273 7711 16331 7717
rect 16273 7708 16285 7711
rect 15767 7680 16285 7708
rect 15767 7677 15779 7680
rect 15721 7671 15779 7677
rect 16273 7677 16285 7680
rect 16319 7677 16331 7711
rect 16273 7671 16331 7677
rect 16917 7711 16975 7717
rect 16917 7677 16929 7711
rect 16963 7708 16975 7711
rect 17469 7711 17527 7717
rect 17469 7708 17481 7711
rect 16963 7680 17481 7708
rect 16963 7677 16975 7680
rect 16917 7671 16975 7677
rect 17469 7677 17481 7680
rect 17515 7677 17527 7711
rect 17469 7671 17527 7677
rect 18113 7711 18171 7717
rect 18113 7677 18125 7711
rect 18159 7708 18171 7711
rect 18665 7711 18723 7717
rect 18665 7708 18677 7711
rect 18159 7680 18677 7708
rect 18159 7677 18171 7680
rect 18113 7671 18171 7677
rect 18665 7677 18677 7680
rect 18711 7677 18723 7711
rect 18665 7671 18723 7677
rect 19309 7711 19367 7717
rect 19309 7677 19321 7711
rect 19355 7708 19367 7711
rect 19861 7711 19919 7717
rect 19861 7708 19873 7711
rect 19355 7680 19873 7708
rect 19355 7677 19367 7680
rect 19309 7671 19367 7677
rect 19861 7677 19873 7680
rect 19907 7677 19919 7711
rect 19861 7671 19919 7677
rect 20505 7711 20563 7717
rect 20505 7677 20517 7711
rect 20551 7708 20563 7711
rect 21057 7711 21115 7717
rect 21057 7708 21069 7711
rect 20551 7680 21069 7708
rect 20551 7677 20563 7680
rect 20505 7671 20563 7677
rect 21057 7677 21069 7680
rect 21103 7677 21115 7711
rect 21057 7671 21115 7677
rect 1904 7482 22236 7504
rect 1904 7430 7110 7482
rect 7162 7430 7174 7482
rect 7226 7430 7238 7482
rect 7290 7430 7302 7482
rect 7354 7430 12438 7482
rect 12490 7430 12502 7482
rect 12554 7430 12566 7482
rect 12618 7430 12630 7482
rect 12682 7430 17766 7482
rect 17818 7430 17830 7482
rect 17882 7430 17894 7482
rect 17946 7430 17958 7482
rect 18010 7430 22236 7482
rect 1904 7408 22236 7430
rect 11320 7272 11624 7300
rect 3117 7167 3175 7173
rect 3117 7133 3129 7167
rect 3163 7133 3175 7167
rect 3117 7127 3175 7133
rect 3761 7167 3819 7173
rect 3761 7133 3773 7167
rect 3807 7164 3819 7167
rect 3850 7164 3856 7176
rect 3807 7136 3856 7164
rect 3807 7133 3819 7136
rect 3761 7127 3819 7133
rect 3132 7096 3160 7127
rect 3850 7124 3856 7136
rect 3908 7124 3914 7176
rect 4313 7167 4371 7173
rect 4313 7133 4325 7167
rect 4359 7164 4371 7167
rect 5509 7167 5567 7173
rect 4359 7136 5276 7164
rect 4359 7133 4371 7136
rect 4313 7127 4371 7133
rect 4957 7099 5015 7105
rect 4957 7096 4969 7099
rect 3132 7068 4969 7096
rect 4957 7065 4969 7068
rect 5003 7065 5015 7099
rect 4957 7059 5015 7065
rect 5248 7028 5276 7136
rect 5509 7133 5521 7167
rect 5555 7133 5567 7167
rect 5509 7127 5567 7133
rect 6705 7167 6763 7173
rect 6705 7133 6717 7167
rect 6751 7164 6763 7167
rect 7901 7167 7959 7173
rect 6751 7136 7852 7164
rect 6751 7133 6763 7136
rect 6705 7127 6763 7133
rect 5524 7096 5552 7127
rect 7349 7099 7407 7105
rect 7349 7096 7361 7099
rect 5524 7068 7361 7096
rect 7349 7065 7361 7068
rect 7395 7065 7407 7099
rect 7824 7096 7852 7136
rect 7901 7133 7913 7167
rect 7947 7164 7959 7167
rect 9097 7167 9155 7173
rect 7947 7136 8864 7164
rect 7947 7133 7959 7136
rect 7901 7127 7959 7133
rect 8545 7099 8603 7105
rect 8545 7096 8557 7099
rect 7824 7068 8557 7096
rect 7349 7059 7407 7065
rect 8545 7065 8557 7068
rect 8591 7065 8603 7099
rect 8836 7096 8864 7136
rect 9097 7133 9109 7167
rect 9143 7164 9155 7167
rect 10293 7167 10351 7173
rect 9143 7136 10060 7164
rect 9143 7133 9155 7136
rect 9097 7127 9155 7133
rect 9741 7099 9799 7105
rect 9741 7096 9753 7099
rect 8836 7068 9753 7096
rect 8545 7059 8603 7065
rect 9741 7065 9753 7068
rect 9787 7065 9799 7099
rect 9741 7059 9799 7065
rect 6153 7031 6211 7037
rect 6153 7028 6165 7031
rect 5248 7000 6165 7028
rect 6153 6997 6165 7000
rect 6199 6997 6211 7031
rect 10032 7028 10060 7136
rect 10293 7133 10305 7167
rect 10339 7164 10351 7167
rect 11320 7164 11348 7272
rect 11489 7235 11547 7241
rect 11489 7232 11501 7235
rect 10339 7136 11348 7164
rect 11412 7204 11501 7232
rect 10339 7133 10351 7136
rect 10293 7127 10351 7133
rect 10937 7031 10995 7037
rect 10937 7028 10949 7031
rect 10032 7000 10949 7028
rect 6153 6991 6211 6997
rect 10937 6997 10949 7000
rect 10983 6997 10995 7031
rect 11412 7028 11440 7204
rect 11489 7201 11501 7204
rect 11535 7201 11547 7235
rect 11489 7195 11547 7201
rect 11596 7164 11624 7272
rect 13712 7272 14016 7300
rect 12133 7167 12191 7173
rect 12133 7164 12145 7167
rect 11596 7136 12145 7164
rect 12133 7133 12145 7136
rect 12179 7133 12191 7167
rect 12133 7127 12191 7133
rect 12685 7167 12743 7173
rect 12685 7133 12697 7167
rect 12731 7164 12743 7167
rect 13712 7164 13740 7272
rect 13881 7235 13939 7241
rect 13881 7232 13893 7235
rect 12731 7136 13740 7164
rect 13804 7204 13893 7232
rect 12731 7133 12743 7136
rect 12685 7127 12743 7133
rect 13329 7031 13387 7037
rect 13329 7028 13341 7031
rect 11412 7000 13341 7028
rect 10937 6991 10995 6997
rect 13329 6997 13341 7000
rect 13375 6997 13387 7031
rect 13804 7028 13832 7204
rect 13881 7201 13893 7204
rect 13927 7201 13939 7235
rect 13881 7195 13939 7201
rect 13988 7164 14016 7272
rect 14525 7167 14583 7173
rect 14525 7164 14537 7167
rect 13988 7136 14537 7164
rect 14525 7133 14537 7136
rect 14571 7133 14583 7167
rect 14525 7127 14583 7133
rect 15077 7167 15135 7173
rect 15077 7133 15089 7167
rect 15123 7164 15135 7167
rect 16273 7167 16331 7173
rect 15123 7136 16040 7164
rect 15123 7133 15135 7136
rect 15077 7127 15135 7133
rect 15721 7099 15779 7105
rect 15721 7096 15733 7099
rect 14724 7068 15733 7096
rect 14724 7028 14752 7068
rect 15721 7065 15733 7068
rect 15767 7065 15779 7099
rect 15721 7059 15779 7065
rect 13804 7000 14752 7028
rect 16012 7028 16040 7136
rect 16273 7133 16285 7167
rect 16319 7133 16331 7167
rect 16273 7127 16331 7133
rect 17469 7167 17527 7173
rect 17469 7133 17481 7167
rect 17515 7164 17527 7167
rect 18665 7167 18723 7173
rect 17515 7136 18432 7164
rect 17515 7133 17527 7136
rect 17469 7127 17527 7133
rect 16288 7096 16316 7127
rect 18113 7099 18171 7105
rect 18113 7096 18125 7099
rect 16288 7068 18125 7096
rect 18113 7065 18125 7068
rect 18159 7065 18171 7099
rect 18113 7059 18171 7065
rect 16917 7031 16975 7037
rect 16917 7028 16929 7031
rect 16012 7000 16929 7028
rect 13329 6991 13387 6997
rect 16917 6997 16929 7000
rect 16963 6997 16975 7031
rect 18404 7028 18432 7136
rect 18665 7133 18677 7167
rect 18711 7133 18723 7167
rect 18665 7127 18723 7133
rect 19861 7167 19919 7173
rect 19861 7133 19873 7167
rect 19907 7164 19919 7167
rect 21057 7167 21115 7173
rect 19907 7136 20640 7164
rect 19907 7133 19919 7136
rect 19861 7127 19919 7133
rect 18680 7096 18708 7127
rect 20505 7099 20563 7105
rect 20505 7096 20517 7099
rect 18680 7068 20517 7096
rect 20505 7065 20517 7068
rect 20551 7065 20563 7099
rect 20505 7059 20563 7065
rect 19309 7031 19367 7037
rect 19309 7028 19321 7031
rect 18404 7000 19321 7028
rect 16917 6991 16975 6997
rect 19309 6997 19321 7000
rect 19355 6997 19367 7031
rect 20612 7028 20640 7136
rect 21057 7133 21069 7167
rect 21103 7164 21115 7167
rect 21698 7164 21704 7176
rect 21103 7136 21704 7164
rect 21103 7133 21115 7136
rect 21057 7127 21115 7133
rect 21698 7124 21704 7136
rect 21756 7124 21762 7176
rect 21701 7031 21759 7037
rect 21701 7028 21713 7031
rect 20612 7000 21713 7028
rect 19309 6991 19367 6997
rect 21701 6997 21713 7000
rect 21747 6997 21759 7031
rect 21701 6991 21759 6997
rect 1904 6938 22236 6960
rect 1904 6886 4446 6938
rect 4498 6886 4510 6938
rect 4562 6886 4574 6938
rect 4626 6886 4638 6938
rect 4690 6886 9774 6938
rect 9826 6886 9838 6938
rect 9890 6886 9902 6938
rect 9954 6886 9966 6938
rect 10018 6886 15102 6938
rect 15154 6886 15166 6938
rect 15218 6886 15230 6938
rect 15282 6886 15294 6938
rect 15346 6886 20430 6938
rect 20482 6886 20494 6938
rect 20546 6886 20558 6938
rect 20610 6886 20622 6938
rect 20674 6886 22236 6938
rect 1904 6864 22236 6886
rect 21698 6824 21704 6836
rect 21659 6796 21704 6824
rect 21698 6784 21704 6796
rect 21756 6784 21762 6836
rect 3117 6691 3175 6697
rect 3117 6657 3129 6691
rect 3163 6688 3175 6691
rect 3850 6688 3856 6700
rect 3163 6660 3856 6688
rect 3163 6657 3175 6660
rect 3117 6651 3175 6657
rect 3850 6648 3856 6660
rect 3908 6648 3914 6700
rect 3761 6623 3819 6629
rect 3761 6589 3773 6623
rect 3807 6620 3819 6623
rect 4313 6623 4371 6629
rect 4313 6620 4325 6623
rect 3807 6592 4325 6620
rect 3807 6589 3819 6592
rect 3761 6583 3819 6589
rect 4313 6589 4325 6592
rect 4359 6589 4371 6623
rect 4313 6583 4371 6589
rect 4957 6623 5015 6629
rect 4957 6589 4969 6623
rect 5003 6620 5015 6623
rect 5509 6623 5567 6629
rect 5509 6620 5521 6623
rect 5003 6592 5521 6620
rect 5003 6589 5015 6592
rect 4957 6583 5015 6589
rect 5509 6589 5521 6592
rect 5555 6589 5567 6623
rect 5509 6583 5567 6589
rect 6153 6623 6211 6629
rect 6153 6589 6165 6623
rect 6199 6620 6211 6623
rect 6705 6623 6763 6629
rect 6705 6620 6717 6623
rect 6199 6592 6717 6620
rect 6199 6589 6211 6592
rect 6153 6583 6211 6589
rect 6705 6589 6717 6592
rect 6751 6589 6763 6623
rect 6705 6583 6763 6589
rect 7349 6623 7407 6629
rect 7349 6589 7361 6623
rect 7395 6620 7407 6623
rect 7901 6623 7959 6629
rect 7901 6620 7913 6623
rect 7395 6592 7913 6620
rect 7395 6589 7407 6592
rect 7349 6583 7407 6589
rect 7901 6589 7913 6592
rect 7947 6589 7959 6623
rect 7901 6583 7959 6589
rect 8545 6623 8603 6629
rect 8545 6589 8557 6623
rect 8591 6620 8603 6623
rect 9097 6623 9155 6629
rect 9097 6620 9109 6623
rect 8591 6592 9109 6620
rect 8591 6589 8603 6592
rect 8545 6583 8603 6589
rect 9097 6589 9109 6592
rect 9143 6589 9155 6623
rect 9097 6583 9155 6589
rect 9741 6623 9799 6629
rect 9741 6589 9753 6623
rect 9787 6620 9799 6623
rect 10293 6623 10351 6629
rect 10293 6620 10305 6623
rect 9787 6592 10305 6620
rect 9787 6589 9799 6592
rect 9741 6583 9799 6589
rect 10293 6589 10305 6592
rect 10339 6589 10351 6623
rect 10293 6583 10351 6589
rect 10937 6623 10995 6629
rect 10937 6589 10949 6623
rect 10983 6620 10995 6623
rect 11489 6623 11547 6629
rect 11489 6620 11501 6623
rect 10983 6592 11501 6620
rect 10983 6589 10995 6592
rect 10937 6583 10995 6589
rect 11489 6589 11501 6592
rect 11535 6589 11547 6623
rect 11489 6583 11547 6589
rect 12133 6623 12191 6629
rect 12133 6589 12145 6623
rect 12179 6620 12191 6623
rect 12685 6623 12743 6629
rect 12685 6620 12697 6623
rect 12179 6592 12697 6620
rect 12179 6589 12191 6592
rect 12133 6583 12191 6589
rect 12685 6589 12697 6592
rect 12731 6589 12743 6623
rect 12685 6583 12743 6589
rect 13329 6623 13387 6629
rect 13329 6589 13341 6623
rect 13375 6620 13387 6623
rect 13881 6623 13939 6629
rect 13881 6620 13893 6623
rect 13375 6592 13893 6620
rect 13375 6589 13387 6592
rect 13329 6583 13387 6589
rect 13881 6589 13893 6592
rect 13927 6589 13939 6623
rect 13881 6583 13939 6589
rect 14525 6623 14583 6629
rect 14525 6589 14537 6623
rect 14571 6620 14583 6623
rect 15077 6623 15135 6629
rect 15077 6620 15089 6623
rect 14571 6592 15089 6620
rect 14571 6589 14583 6592
rect 14525 6583 14583 6589
rect 15077 6589 15089 6592
rect 15123 6589 15135 6623
rect 15077 6583 15135 6589
rect 15721 6623 15779 6629
rect 15721 6589 15733 6623
rect 15767 6620 15779 6623
rect 16273 6623 16331 6629
rect 16273 6620 16285 6623
rect 15767 6592 16285 6620
rect 15767 6589 15779 6592
rect 15721 6583 15779 6589
rect 16273 6589 16285 6592
rect 16319 6589 16331 6623
rect 16273 6583 16331 6589
rect 16917 6623 16975 6629
rect 16917 6589 16929 6623
rect 16963 6620 16975 6623
rect 17469 6623 17527 6629
rect 17469 6620 17481 6623
rect 16963 6592 17481 6620
rect 16963 6589 16975 6592
rect 16917 6583 16975 6589
rect 17469 6589 17481 6592
rect 17515 6589 17527 6623
rect 17469 6583 17527 6589
rect 18113 6623 18171 6629
rect 18113 6589 18125 6623
rect 18159 6620 18171 6623
rect 18665 6623 18723 6629
rect 18665 6620 18677 6623
rect 18159 6592 18677 6620
rect 18159 6589 18171 6592
rect 18113 6583 18171 6589
rect 18665 6589 18677 6592
rect 18711 6589 18723 6623
rect 18665 6583 18723 6589
rect 19309 6623 19367 6629
rect 19309 6589 19321 6623
rect 19355 6620 19367 6623
rect 19861 6623 19919 6629
rect 19861 6620 19873 6623
rect 19355 6592 19873 6620
rect 19355 6589 19367 6592
rect 19309 6583 19367 6589
rect 19861 6589 19873 6592
rect 19907 6589 19919 6623
rect 19861 6583 19919 6589
rect 20505 6623 20563 6629
rect 20505 6589 20517 6623
rect 20551 6620 20563 6623
rect 21057 6623 21115 6629
rect 21057 6620 21069 6623
rect 20551 6592 21069 6620
rect 20551 6589 20563 6592
rect 20505 6583 20563 6589
rect 21057 6589 21069 6592
rect 21103 6589 21115 6623
rect 21057 6583 21115 6589
rect 1904 6394 22236 6416
rect 1904 6342 7110 6394
rect 7162 6342 7174 6394
rect 7226 6342 7238 6394
rect 7290 6342 7302 6394
rect 7354 6342 12438 6394
rect 12490 6342 12502 6394
rect 12554 6342 12566 6394
rect 12618 6342 12630 6394
rect 12682 6342 17766 6394
rect 17818 6342 17830 6394
rect 17882 6342 17894 6394
rect 17946 6342 17958 6394
rect 18010 6342 22236 6394
rect 1904 6320 22236 6342
rect 3761 6283 3819 6289
rect 3761 6249 3773 6283
rect 3807 6280 3819 6283
rect 3850 6280 3856 6292
rect 3807 6252 3856 6280
rect 3807 6249 3819 6252
rect 3761 6243 3819 6249
rect 3850 6240 3856 6252
rect 3908 6240 3914 6292
rect 3117 6147 3175 6153
rect 3117 6113 3129 6147
rect 3163 6144 3175 6147
rect 4957 6147 5015 6153
rect 4957 6144 4969 6147
rect 3163 6116 4969 6144
rect 3163 6113 3175 6116
rect 3117 6107 3175 6113
rect 4957 6113 4969 6116
rect 5003 6113 5015 6147
rect 4957 6107 5015 6113
rect 5509 6147 5567 6153
rect 5509 6113 5521 6147
rect 5555 6144 5567 6147
rect 7349 6147 7407 6153
rect 7349 6144 7361 6147
rect 5555 6116 7361 6144
rect 5555 6113 5567 6116
rect 5509 6107 5567 6113
rect 7349 6113 7361 6116
rect 7395 6113 7407 6147
rect 7349 6107 7407 6113
rect 7901 6147 7959 6153
rect 7901 6113 7913 6147
rect 7947 6144 7959 6147
rect 9097 6147 9155 6153
rect 7947 6116 8772 6144
rect 7947 6113 7959 6116
rect 7901 6107 7959 6113
rect 4313 6079 4371 6085
rect 4313 6045 4325 6079
rect 4359 6076 4371 6079
rect 6153 6079 6211 6085
rect 6153 6076 6165 6079
rect 4359 6048 6165 6076
rect 4359 6045 4371 6048
rect 4313 6039 4371 6045
rect 6153 6045 6165 6048
rect 6199 6045 6211 6079
rect 6153 6039 6211 6045
rect 6705 6079 6763 6085
rect 6705 6045 6717 6079
rect 6751 6076 6763 6079
rect 8545 6079 8603 6085
rect 8545 6076 8557 6079
rect 6751 6048 8557 6076
rect 6751 6045 6763 6048
rect 6705 6039 6763 6045
rect 8545 6045 8557 6048
rect 8591 6045 8603 6079
rect 8744 6076 8772 6116
rect 9097 6113 9109 6147
rect 9143 6144 9155 6147
rect 10937 6147 10995 6153
rect 10937 6144 10949 6147
rect 9143 6116 10949 6144
rect 9143 6113 9155 6116
rect 9097 6107 9155 6113
rect 10937 6113 10949 6116
rect 10983 6113 10995 6147
rect 10937 6107 10995 6113
rect 11489 6147 11547 6153
rect 11489 6113 11501 6147
rect 11535 6144 11547 6147
rect 13329 6147 13387 6153
rect 13329 6144 13341 6147
rect 11535 6116 13341 6144
rect 11535 6113 11547 6116
rect 11489 6107 11547 6113
rect 13329 6113 13341 6116
rect 13375 6113 13387 6147
rect 13329 6107 13387 6113
rect 13881 6147 13939 6153
rect 13881 6113 13893 6147
rect 13927 6144 13939 6147
rect 15721 6147 15779 6153
rect 15721 6144 15733 6147
rect 13927 6116 15733 6144
rect 13927 6113 13939 6116
rect 13881 6107 13939 6113
rect 15721 6113 15733 6116
rect 15767 6113 15779 6147
rect 15721 6107 15779 6113
rect 16273 6147 16331 6153
rect 16273 6113 16285 6147
rect 16319 6144 16331 6147
rect 18113 6147 18171 6153
rect 18113 6144 18125 6147
rect 16319 6116 18125 6144
rect 16319 6113 16331 6116
rect 16273 6107 16331 6113
rect 18113 6113 18125 6116
rect 18159 6113 18171 6147
rect 19309 6147 19367 6153
rect 19309 6144 19321 6147
rect 18113 6107 18171 6113
rect 18496 6116 19321 6144
rect 9741 6079 9799 6085
rect 9741 6076 9753 6079
rect 8744 6048 9753 6076
rect 8545 6039 8603 6045
rect 9741 6045 9753 6048
rect 9787 6045 9799 6079
rect 9741 6039 9799 6045
rect 10293 6079 10351 6085
rect 10293 6045 10305 6079
rect 10339 6076 10351 6079
rect 12133 6079 12191 6085
rect 12133 6076 12145 6079
rect 10339 6048 12145 6076
rect 10339 6045 10351 6048
rect 10293 6039 10351 6045
rect 12133 6045 12145 6048
rect 12179 6045 12191 6079
rect 12133 6039 12191 6045
rect 12685 6079 12743 6085
rect 12685 6045 12697 6079
rect 12731 6076 12743 6079
rect 14525 6079 14583 6085
rect 14525 6076 14537 6079
rect 12731 6048 14537 6076
rect 12731 6045 12743 6048
rect 12685 6039 12743 6045
rect 14525 6045 14537 6048
rect 14571 6045 14583 6079
rect 14525 6039 14583 6045
rect 15077 6079 15135 6085
rect 15077 6045 15089 6079
rect 15123 6076 15135 6079
rect 16917 6079 16975 6085
rect 16917 6076 16929 6079
rect 15123 6048 16929 6076
rect 15123 6045 15135 6048
rect 15077 6039 15135 6045
rect 16917 6045 16929 6048
rect 16963 6045 16975 6079
rect 16917 6039 16975 6045
rect 17469 6079 17527 6085
rect 17469 6045 17481 6079
rect 17515 6076 17527 6079
rect 18496 6076 18524 6116
rect 19309 6113 19321 6116
rect 19355 6113 19367 6147
rect 19309 6107 19367 6113
rect 19861 6147 19919 6153
rect 19861 6113 19873 6147
rect 19907 6144 19919 6147
rect 21701 6147 21759 6153
rect 21701 6144 21713 6147
rect 19907 6116 21713 6144
rect 19907 6113 19919 6116
rect 19861 6107 19919 6113
rect 21701 6113 21713 6116
rect 21747 6113 21759 6147
rect 21701 6107 21759 6113
rect 17515 6048 18524 6076
rect 18665 6079 18723 6085
rect 17515 6045 17527 6048
rect 17469 6039 17527 6045
rect 18665 6045 18677 6079
rect 18711 6076 18723 6079
rect 20505 6079 20563 6085
rect 20505 6076 20517 6079
rect 18711 6048 20517 6076
rect 18711 6045 18723 6048
rect 18665 6039 18723 6045
rect 20505 6045 20517 6048
rect 20551 6045 20563 6079
rect 20505 6039 20563 6045
rect 21057 6079 21115 6085
rect 21057 6045 21069 6079
rect 21103 6076 21115 6079
rect 21606 6076 21612 6088
rect 21103 6048 21612 6076
rect 21103 6045 21115 6048
rect 21057 6039 21115 6045
rect 21606 6036 21612 6048
rect 21664 6036 21670 6088
rect 1904 5850 22236 5872
rect 1904 5798 4446 5850
rect 4498 5798 4510 5850
rect 4562 5798 4574 5850
rect 4626 5798 4638 5850
rect 4690 5798 9774 5850
rect 9826 5798 9838 5850
rect 9890 5798 9902 5850
rect 9954 5798 9966 5850
rect 10018 5798 15102 5850
rect 15154 5798 15166 5850
rect 15218 5798 15230 5850
rect 15282 5798 15294 5850
rect 15346 5798 20430 5850
rect 20482 5798 20494 5850
rect 20546 5798 20558 5850
rect 20610 5798 20622 5850
rect 20674 5798 22236 5850
rect 1904 5776 22236 5798
rect 21606 5696 21612 5748
rect 21664 5736 21670 5748
rect 21701 5739 21759 5745
rect 21701 5736 21713 5739
rect 21664 5708 21713 5736
rect 21664 5696 21670 5708
rect 21701 5705 21713 5708
rect 21747 5705 21759 5739
rect 21701 5699 21759 5705
rect 3117 5603 3175 5609
rect 3117 5569 3129 5603
rect 3163 5600 3175 5603
rect 3850 5600 3856 5612
rect 3163 5572 3856 5600
rect 3163 5569 3175 5572
rect 3117 5563 3175 5569
rect 3850 5560 3856 5572
rect 3908 5560 3914 5612
rect 3761 5535 3819 5541
rect 3761 5501 3773 5535
rect 3807 5532 3819 5535
rect 4313 5535 4371 5541
rect 4313 5532 4325 5535
rect 3807 5504 4325 5532
rect 3807 5501 3819 5504
rect 3761 5495 3819 5501
rect 4313 5501 4325 5504
rect 4359 5501 4371 5535
rect 4313 5495 4371 5501
rect 4957 5535 5015 5541
rect 4957 5501 4969 5535
rect 5003 5532 5015 5535
rect 5509 5535 5567 5541
rect 5509 5532 5521 5535
rect 5003 5504 5521 5532
rect 5003 5501 5015 5504
rect 4957 5495 5015 5501
rect 5509 5501 5521 5504
rect 5555 5501 5567 5535
rect 5509 5495 5567 5501
rect 6153 5535 6211 5541
rect 6153 5501 6165 5535
rect 6199 5532 6211 5535
rect 6705 5535 6763 5541
rect 6705 5532 6717 5535
rect 6199 5504 6717 5532
rect 6199 5501 6211 5504
rect 6153 5495 6211 5501
rect 6705 5501 6717 5504
rect 6751 5501 6763 5535
rect 6705 5495 6763 5501
rect 7349 5535 7407 5541
rect 7349 5501 7361 5535
rect 7395 5532 7407 5535
rect 7901 5535 7959 5541
rect 7901 5532 7913 5535
rect 7395 5504 7913 5532
rect 7395 5501 7407 5504
rect 7349 5495 7407 5501
rect 7901 5501 7913 5504
rect 7947 5501 7959 5535
rect 7901 5495 7959 5501
rect 8545 5535 8603 5541
rect 8545 5501 8557 5535
rect 8591 5532 8603 5535
rect 9097 5535 9155 5541
rect 9097 5532 9109 5535
rect 8591 5504 9109 5532
rect 8591 5501 8603 5504
rect 8545 5495 8603 5501
rect 9097 5501 9109 5504
rect 9143 5501 9155 5535
rect 9097 5495 9155 5501
rect 9741 5535 9799 5541
rect 9741 5501 9753 5535
rect 9787 5532 9799 5535
rect 10293 5535 10351 5541
rect 10293 5532 10305 5535
rect 9787 5504 10305 5532
rect 9787 5501 9799 5504
rect 9741 5495 9799 5501
rect 10293 5501 10305 5504
rect 10339 5501 10351 5535
rect 10293 5495 10351 5501
rect 10937 5535 10995 5541
rect 10937 5501 10949 5535
rect 10983 5532 10995 5535
rect 11489 5535 11547 5541
rect 11489 5532 11501 5535
rect 10983 5504 11501 5532
rect 10983 5501 10995 5504
rect 10937 5495 10995 5501
rect 11489 5501 11501 5504
rect 11535 5501 11547 5535
rect 11489 5495 11547 5501
rect 12133 5535 12191 5541
rect 12133 5501 12145 5535
rect 12179 5532 12191 5535
rect 12685 5535 12743 5541
rect 12685 5532 12697 5535
rect 12179 5504 12697 5532
rect 12179 5501 12191 5504
rect 12133 5495 12191 5501
rect 12685 5501 12697 5504
rect 12731 5501 12743 5535
rect 12685 5495 12743 5501
rect 13329 5535 13387 5541
rect 13329 5501 13341 5535
rect 13375 5532 13387 5535
rect 13881 5535 13939 5541
rect 13881 5532 13893 5535
rect 13375 5504 13893 5532
rect 13375 5501 13387 5504
rect 13329 5495 13387 5501
rect 13881 5501 13893 5504
rect 13927 5501 13939 5535
rect 13881 5495 13939 5501
rect 14525 5535 14583 5541
rect 14525 5501 14537 5535
rect 14571 5532 14583 5535
rect 15077 5535 15135 5541
rect 15077 5532 15089 5535
rect 14571 5504 15089 5532
rect 14571 5501 14583 5504
rect 14525 5495 14583 5501
rect 15077 5501 15089 5504
rect 15123 5501 15135 5535
rect 15077 5495 15135 5501
rect 15721 5535 15779 5541
rect 15721 5501 15733 5535
rect 15767 5532 15779 5535
rect 16273 5535 16331 5541
rect 16273 5532 16285 5535
rect 15767 5504 16285 5532
rect 15767 5501 15779 5504
rect 15721 5495 15779 5501
rect 16273 5501 16285 5504
rect 16319 5501 16331 5535
rect 16273 5495 16331 5501
rect 16917 5535 16975 5541
rect 16917 5501 16929 5535
rect 16963 5532 16975 5535
rect 17469 5535 17527 5541
rect 17469 5532 17481 5535
rect 16963 5504 17481 5532
rect 16963 5501 16975 5504
rect 16917 5495 16975 5501
rect 17469 5501 17481 5504
rect 17515 5501 17527 5535
rect 17469 5495 17527 5501
rect 18113 5535 18171 5541
rect 18113 5501 18125 5535
rect 18159 5532 18171 5535
rect 18665 5535 18723 5541
rect 18665 5532 18677 5535
rect 18159 5504 18677 5532
rect 18159 5501 18171 5504
rect 18113 5495 18171 5501
rect 18665 5501 18677 5504
rect 18711 5501 18723 5535
rect 18665 5495 18723 5501
rect 19309 5535 19367 5541
rect 19309 5501 19321 5535
rect 19355 5532 19367 5535
rect 19861 5535 19919 5541
rect 19861 5532 19873 5535
rect 19355 5504 19873 5532
rect 19355 5501 19367 5504
rect 19309 5495 19367 5501
rect 19861 5501 19873 5504
rect 19907 5501 19919 5535
rect 19861 5495 19919 5501
rect 20505 5535 20563 5541
rect 20505 5501 20517 5535
rect 20551 5532 20563 5535
rect 21057 5535 21115 5541
rect 21057 5532 21069 5535
rect 20551 5504 21069 5532
rect 20551 5501 20563 5504
rect 20505 5495 20563 5501
rect 21057 5501 21069 5504
rect 21103 5501 21115 5535
rect 21057 5495 21115 5501
rect 1904 5306 22236 5328
rect 1904 5254 7110 5306
rect 7162 5254 7174 5306
rect 7226 5254 7238 5306
rect 7290 5254 7302 5306
rect 7354 5254 12438 5306
rect 12490 5254 12502 5306
rect 12554 5254 12566 5306
rect 12618 5254 12630 5306
rect 12682 5254 17766 5306
rect 17818 5254 17830 5306
rect 17882 5254 17894 5306
rect 17946 5254 17958 5306
rect 18010 5254 22236 5306
rect 1904 5232 22236 5254
rect 12133 5195 12191 5201
rect 12133 5192 12145 5195
rect 10308 5164 12145 5192
rect 6153 5127 6211 5133
rect 6153 5124 6165 5127
rect 4328 5096 6165 5124
rect 4328 5065 4356 5096
rect 6153 5093 6165 5096
rect 6199 5093 6211 5127
rect 9741 5127 9799 5133
rect 9741 5124 9753 5127
rect 6153 5087 6211 5093
rect 7916 5096 9753 5124
rect 7916 5065 7944 5096
rect 9741 5093 9753 5096
rect 9787 5093 9799 5127
rect 9741 5087 9799 5093
rect 10308 5065 10336 5164
rect 12133 5161 12145 5164
rect 12179 5161 12191 5195
rect 12133 5155 12191 5161
rect 13329 5127 13387 5133
rect 13329 5124 13341 5127
rect 11504 5096 13341 5124
rect 11504 5065 11532 5096
rect 13329 5093 13341 5096
rect 13375 5093 13387 5127
rect 15721 5127 15779 5133
rect 15721 5124 15733 5127
rect 13329 5087 13387 5093
rect 13896 5096 15733 5124
rect 13896 5065 13924 5096
rect 15721 5093 15733 5096
rect 15767 5093 15779 5127
rect 19309 5127 19367 5133
rect 19309 5124 19321 5127
rect 15721 5087 15779 5093
rect 17484 5096 19321 5124
rect 3117 5059 3175 5065
rect 3117 5025 3129 5059
rect 3163 5056 3175 5059
rect 4313 5059 4371 5065
rect 3163 5028 4080 5056
rect 3163 5025 3175 5028
rect 3117 5019 3175 5025
rect 3761 4991 3819 4997
rect 3761 4957 3773 4991
rect 3807 4988 3819 4991
rect 3850 4988 3856 5000
rect 3807 4960 3856 4988
rect 3807 4957 3819 4960
rect 3761 4951 3819 4957
rect 3850 4948 3856 4960
rect 3908 4948 3914 5000
rect 4052 4988 4080 5028
rect 4313 5025 4325 5059
rect 4359 5025 4371 5059
rect 4313 5019 4371 5025
rect 5509 5059 5567 5065
rect 5509 5025 5521 5059
rect 5555 5056 5567 5059
rect 6705 5059 6763 5065
rect 5555 5028 6472 5056
rect 5555 5025 5567 5028
rect 5509 5019 5567 5025
rect 4957 4991 5015 4997
rect 4957 4988 4969 4991
rect 4052 4960 4969 4988
rect 4957 4957 4969 4960
rect 5003 4957 5015 4991
rect 6444 4988 6472 5028
rect 6705 5025 6717 5059
rect 6751 5056 6763 5059
rect 7901 5059 7959 5065
rect 6751 5028 7668 5056
rect 6751 5025 6763 5028
rect 6705 5019 6763 5025
rect 7349 4991 7407 4997
rect 7349 4988 7361 4991
rect 6444 4960 7361 4988
rect 4957 4951 5015 4957
rect 7349 4957 7361 4960
rect 7395 4957 7407 4991
rect 7640 4988 7668 5028
rect 7901 5025 7913 5059
rect 7947 5025 7959 5059
rect 7901 5019 7959 5025
rect 9097 5059 9155 5065
rect 9097 5025 9109 5059
rect 9143 5056 9155 5059
rect 10293 5059 10351 5065
rect 9143 5028 10244 5056
rect 9143 5025 9155 5028
rect 9097 5019 9155 5025
rect 8545 4991 8603 4997
rect 8545 4988 8557 4991
rect 7640 4960 8557 4988
rect 7349 4951 7407 4957
rect 8545 4957 8557 4960
rect 8591 4957 8603 4991
rect 8545 4951 8603 4957
rect 10216 4920 10244 5028
rect 10293 5025 10305 5059
rect 10339 5025 10351 5059
rect 10293 5019 10351 5025
rect 11489 5059 11547 5065
rect 11489 5025 11501 5059
rect 11535 5025 11547 5059
rect 11489 5019 11547 5025
rect 12685 5059 12743 5065
rect 12685 5025 12697 5059
rect 12731 5056 12743 5059
rect 13881 5059 13939 5065
rect 12731 5028 13648 5056
rect 12731 5025 12743 5028
rect 12685 5019 12743 5025
rect 13620 4988 13648 5028
rect 13881 5025 13893 5059
rect 13927 5025 13939 5059
rect 13881 5019 13939 5025
rect 15077 5059 15135 5065
rect 15077 5025 15089 5059
rect 15123 5056 15135 5059
rect 16273 5059 16331 5065
rect 15123 5028 16040 5056
rect 15123 5025 15135 5028
rect 15077 5019 15135 5025
rect 14525 4991 14583 4997
rect 14525 4988 14537 4991
rect 13620 4960 14537 4988
rect 14525 4957 14537 4960
rect 14571 4957 14583 4991
rect 16012 4988 16040 5028
rect 16273 5025 16285 5059
rect 16319 5056 16331 5059
rect 17374 5056 17380 5068
rect 16319 5028 17380 5056
rect 16319 5025 16331 5028
rect 16273 5019 16331 5025
rect 17374 5016 17380 5028
rect 17432 5016 17438 5068
rect 17484 4997 17512 5096
rect 19309 5093 19321 5096
rect 19355 5093 19367 5127
rect 19309 5087 19367 5093
rect 18665 5059 18723 5065
rect 18665 5025 18677 5059
rect 18711 5056 18723 5059
rect 19861 5059 19919 5065
rect 18711 5028 19444 5056
rect 18711 5025 18723 5028
rect 18665 5019 18723 5025
rect 16917 4991 16975 4997
rect 16917 4988 16929 4991
rect 16012 4960 16929 4988
rect 14525 4951 14583 4957
rect 16917 4957 16929 4960
rect 16963 4957 16975 4991
rect 16917 4951 16975 4957
rect 17469 4991 17527 4997
rect 17469 4957 17481 4991
rect 17515 4957 17527 4991
rect 17469 4951 17527 4957
rect 17558 4948 17564 5000
rect 17616 4988 17622 5000
rect 18113 4991 18171 4997
rect 18113 4988 18125 4991
rect 17616 4960 18125 4988
rect 17616 4948 17622 4960
rect 18113 4957 18125 4960
rect 18159 4957 18171 4991
rect 19416 4988 19444 5028
rect 19861 5025 19873 5059
rect 19907 5056 19919 5059
rect 21701 5059 21759 5065
rect 21701 5056 21713 5059
rect 19907 5028 21713 5056
rect 19907 5025 19919 5028
rect 19861 5019 19919 5025
rect 21701 5025 21713 5028
rect 21747 5025 21759 5059
rect 21701 5019 21759 5025
rect 20505 4991 20563 4997
rect 20505 4988 20517 4991
rect 19416 4960 20517 4988
rect 18113 4951 18171 4957
rect 20505 4957 20517 4960
rect 20551 4957 20563 4991
rect 20505 4951 20563 4957
rect 21057 4991 21115 4997
rect 21057 4957 21069 4991
rect 21103 4988 21115 4991
rect 21606 4988 21612 5000
rect 21103 4960 21612 4988
rect 21103 4957 21115 4960
rect 21057 4951 21115 4957
rect 21606 4948 21612 4960
rect 21664 4948 21670 5000
rect 10937 4923 10995 4929
rect 10937 4920 10949 4923
rect 10216 4892 10949 4920
rect 10937 4889 10949 4892
rect 10983 4889 10995 4923
rect 10937 4883 10995 4889
rect 1904 4762 22236 4784
rect 1904 4710 4446 4762
rect 4498 4710 4510 4762
rect 4562 4710 4574 4762
rect 4626 4710 4638 4762
rect 4690 4710 9774 4762
rect 9826 4710 9838 4762
rect 9890 4710 9902 4762
rect 9954 4710 9966 4762
rect 10018 4710 15102 4762
rect 15154 4710 15166 4762
rect 15218 4710 15230 4762
rect 15282 4710 15294 4762
rect 15346 4710 20430 4762
rect 20482 4710 20494 4762
rect 20546 4710 20558 4762
rect 20610 4710 20622 4762
rect 20674 4710 22236 4762
rect 1904 4688 22236 4710
rect 21606 4608 21612 4660
rect 21664 4648 21670 4660
rect 21701 4651 21759 4657
rect 21701 4648 21713 4651
rect 21664 4620 21713 4648
rect 21664 4608 21670 4620
rect 21701 4617 21713 4620
rect 21747 4617 21759 4651
rect 21701 4611 21759 4617
rect 3117 4515 3175 4521
rect 3117 4481 3129 4515
rect 3163 4512 3175 4515
rect 3850 4512 3856 4524
rect 3163 4484 3856 4512
rect 3163 4481 3175 4484
rect 3117 4475 3175 4481
rect 3850 4472 3856 4484
rect 3908 4472 3914 4524
rect 3761 4447 3819 4453
rect 3761 4413 3773 4447
rect 3807 4444 3819 4447
rect 4313 4447 4371 4453
rect 4313 4444 4325 4447
rect 3807 4416 4325 4444
rect 3807 4413 3819 4416
rect 3761 4407 3819 4413
rect 4313 4413 4325 4416
rect 4359 4413 4371 4447
rect 4313 4407 4371 4413
rect 4957 4447 5015 4453
rect 4957 4413 4969 4447
rect 5003 4444 5015 4447
rect 5509 4447 5567 4453
rect 5509 4444 5521 4447
rect 5003 4416 5521 4444
rect 5003 4413 5015 4416
rect 4957 4407 5015 4413
rect 5509 4413 5521 4416
rect 5555 4413 5567 4447
rect 5509 4407 5567 4413
rect 6153 4447 6211 4453
rect 6153 4413 6165 4447
rect 6199 4444 6211 4447
rect 6705 4447 6763 4453
rect 6705 4444 6717 4447
rect 6199 4416 6717 4444
rect 6199 4413 6211 4416
rect 6153 4407 6211 4413
rect 6705 4413 6717 4416
rect 6751 4413 6763 4447
rect 6705 4407 6763 4413
rect 7349 4447 7407 4453
rect 7349 4413 7361 4447
rect 7395 4444 7407 4447
rect 7901 4447 7959 4453
rect 7901 4444 7913 4447
rect 7395 4416 7913 4444
rect 7395 4413 7407 4416
rect 7349 4407 7407 4413
rect 7901 4413 7913 4416
rect 7947 4413 7959 4447
rect 7901 4407 7959 4413
rect 8545 4447 8603 4453
rect 8545 4413 8557 4447
rect 8591 4444 8603 4447
rect 9097 4447 9155 4453
rect 9097 4444 9109 4447
rect 8591 4416 9109 4444
rect 8591 4413 8603 4416
rect 8545 4407 8603 4413
rect 9097 4413 9109 4416
rect 9143 4413 9155 4447
rect 9097 4407 9155 4413
rect 9741 4447 9799 4453
rect 9741 4413 9753 4447
rect 9787 4444 9799 4447
rect 10293 4447 10351 4453
rect 10293 4444 10305 4447
rect 9787 4416 10305 4444
rect 9787 4413 9799 4416
rect 9741 4407 9799 4413
rect 10293 4413 10305 4416
rect 10339 4413 10351 4447
rect 10293 4407 10351 4413
rect 10937 4447 10995 4453
rect 10937 4413 10949 4447
rect 10983 4444 10995 4447
rect 11489 4447 11547 4453
rect 11489 4444 11501 4447
rect 10983 4416 11501 4444
rect 10983 4413 10995 4416
rect 10937 4407 10995 4413
rect 11489 4413 11501 4416
rect 11535 4413 11547 4447
rect 11489 4407 11547 4413
rect 12133 4447 12191 4453
rect 12133 4413 12145 4447
rect 12179 4444 12191 4447
rect 12685 4447 12743 4453
rect 12685 4444 12697 4447
rect 12179 4416 12697 4444
rect 12179 4413 12191 4416
rect 12133 4407 12191 4413
rect 12685 4413 12697 4416
rect 12731 4413 12743 4447
rect 12685 4407 12743 4413
rect 13329 4447 13387 4453
rect 13329 4413 13341 4447
rect 13375 4444 13387 4447
rect 13881 4447 13939 4453
rect 13881 4444 13893 4447
rect 13375 4416 13893 4444
rect 13375 4413 13387 4416
rect 13329 4407 13387 4413
rect 13881 4413 13893 4416
rect 13927 4413 13939 4447
rect 13881 4407 13939 4413
rect 14525 4447 14583 4453
rect 14525 4413 14537 4447
rect 14571 4444 14583 4447
rect 15077 4447 15135 4453
rect 15077 4444 15089 4447
rect 14571 4416 15089 4444
rect 14571 4413 14583 4416
rect 14525 4407 14583 4413
rect 15077 4413 15089 4416
rect 15123 4413 15135 4447
rect 15077 4407 15135 4413
rect 15721 4447 15779 4453
rect 15721 4413 15733 4447
rect 15767 4444 15779 4447
rect 16273 4447 16331 4453
rect 16273 4444 16285 4447
rect 15767 4416 16285 4444
rect 15767 4413 15779 4416
rect 15721 4407 15779 4413
rect 16273 4413 16285 4416
rect 16319 4413 16331 4447
rect 16273 4407 16331 4413
rect 16917 4447 16975 4453
rect 16917 4413 16929 4447
rect 16963 4444 16975 4447
rect 17469 4447 17527 4453
rect 17469 4444 17481 4447
rect 16963 4416 17481 4444
rect 16963 4413 16975 4416
rect 16917 4407 16975 4413
rect 17469 4413 17481 4416
rect 17515 4413 17527 4447
rect 17469 4407 17527 4413
rect 18113 4447 18171 4453
rect 18113 4413 18125 4447
rect 18159 4444 18171 4447
rect 18665 4447 18723 4453
rect 18665 4444 18677 4447
rect 18159 4416 18677 4444
rect 18159 4413 18171 4416
rect 18113 4407 18171 4413
rect 18665 4413 18677 4416
rect 18711 4413 18723 4447
rect 18665 4407 18723 4413
rect 19309 4447 19367 4453
rect 19309 4413 19321 4447
rect 19355 4444 19367 4447
rect 19861 4447 19919 4453
rect 19861 4444 19873 4447
rect 19355 4416 19873 4444
rect 19355 4413 19367 4416
rect 19309 4407 19367 4413
rect 19861 4413 19873 4416
rect 19907 4413 19919 4447
rect 19861 4407 19919 4413
rect 20505 4447 20563 4453
rect 20505 4413 20517 4447
rect 20551 4444 20563 4447
rect 21057 4447 21115 4453
rect 21057 4444 21069 4447
rect 20551 4416 21069 4444
rect 20551 4413 20563 4416
rect 20505 4407 20563 4413
rect 21057 4413 21069 4416
rect 21103 4413 21115 4447
rect 21057 4407 21115 4413
rect 1904 4218 22236 4240
rect 1904 4166 7110 4218
rect 7162 4166 7174 4218
rect 7226 4166 7238 4218
rect 7290 4166 7302 4218
rect 7354 4166 12438 4218
rect 12490 4166 12502 4218
rect 12554 4166 12566 4218
rect 12618 4166 12630 4218
rect 12682 4166 17766 4218
rect 17818 4166 17830 4218
rect 17882 4166 17894 4218
rect 17946 4166 17958 4218
rect 18010 4166 22236 4218
rect 1904 4144 22236 4166
rect 3761 4107 3819 4113
rect 3761 4073 3773 4107
rect 3807 4104 3819 4107
rect 3850 4104 3856 4116
rect 3807 4076 3856 4104
rect 3807 4073 3819 4076
rect 3761 4067 3819 4073
rect 3850 4064 3856 4076
rect 3908 4064 3914 4116
rect 3117 3971 3175 3977
rect 3117 3937 3129 3971
rect 3163 3968 3175 3971
rect 4957 3971 5015 3977
rect 4957 3968 4969 3971
rect 3163 3940 4969 3968
rect 3163 3937 3175 3940
rect 3117 3931 3175 3937
rect 4957 3937 4969 3940
rect 5003 3937 5015 3971
rect 4957 3931 5015 3937
rect 5509 3971 5567 3977
rect 5509 3937 5521 3971
rect 5555 3968 5567 3971
rect 7349 3971 7407 3977
rect 7349 3968 7361 3971
rect 5555 3940 7361 3968
rect 5555 3937 5567 3940
rect 5509 3931 5567 3937
rect 7349 3937 7361 3940
rect 7395 3937 7407 3971
rect 7349 3931 7407 3937
rect 7901 3971 7959 3977
rect 7901 3937 7913 3971
rect 7947 3968 7959 3971
rect 9097 3971 9155 3977
rect 7947 3940 8772 3968
rect 7947 3937 7959 3940
rect 7901 3931 7959 3937
rect 4313 3903 4371 3909
rect 4313 3869 4325 3903
rect 4359 3900 4371 3903
rect 6153 3903 6211 3909
rect 6153 3900 6165 3903
rect 4359 3872 6165 3900
rect 4359 3869 4371 3872
rect 4313 3863 4371 3869
rect 6153 3869 6165 3872
rect 6199 3869 6211 3903
rect 6153 3863 6211 3869
rect 6705 3903 6763 3909
rect 6705 3869 6717 3903
rect 6751 3900 6763 3903
rect 8545 3903 8603 3909
rect 8545 3900 8557 3903
rect 6751 3872 8557 3900
rect 6751 3869 6763 3872
rect 6705 3863 6763 3869
rect 8545 3869 8557 3872
rect 8591 3869 8603 3903
rect 8744 3900 8772 3940
rect 9097 3937 9109 3971
rect 9143 3968 9155 3971
rect 10937 3971 10995 3977
rect 10937 3968 10949 3971
rect 9143 3940 10949 3968
rect 9143 3937 9155 3940
rect 9097 3931 9155 3937
rect 10937 3937 10949 3940
rect 10983 3937 10995 3971
rect 10937 3931 10995 3937
rect 11489 3971 11547 3977
rect 11489 3937 11501 3971
rect 11535 3968 11547 3971
rect 13329 3971 13387 3977
rect 13329 3968 13341 3971
rect 11535 3940 13341 3968
rect 11535 3937 11547 3940
rect 11489 3931 11547 3937
rect 13329 3937 13341 3940
rect 13375 3937 13387 3971
rect 13329 3931 13387 3937
rect 13881 3971 13939 3977
rect 13881 3937 13893 3971
rect 13927 3968 13939 3971
rect 15721 3971 15779 3977
rect 15721 3968 15733 3971
rect 13927 3940 15733 3968
rect 13927 3937 13939 3940
rect 13881 3931 13939 3937
rect 15721 3937 15733 3940
rect 15767 3937 15779 3971
rect 15721 3931 15779 3937
rect 16273 3971 16331 3977
rect 16273 3937 16285 3971
rect 16319 3968 16331 3971
rect 18113 3971 18171 3977
rect 18113 3968 18125 3971
rect 16319 3940 18125 3968
rect 16319 3937 16331 3940
rect 16273 3931 16331 3937
rect 18113 3937 18125 3940
rect 18159 3937 18171 3971
rect 19309 3971 19367 3977
rect 19309 3968 19321 3971
rect 18113 3931 18171 3937
rect 18496 3940 19321 3968
rect 9741 3903 9799 3909
rect 9741 3900 9753 3903
rect 8744 3872 9753 3900
rect 8545 3863 8603 3869
rect 9741 3869 9753 3872
rect 9787 3869 9799 3903
rect 9741 3863 9799 3869
rect 10293 3903 10351 3909
rect 10293 3869 10305 3903
rect 10339 3900 10351 3903
rect 12133 3903 12191 3909
rect 12133 3900 12145 3903
rect 10339 3872 12145 3900
rect 10339 3869 10351 3872
rect 10293 3863 10351 3869
rect 12133 3869 12145 3872
rect 12179 3869 12191 3903
rect 12133 3863 12191 3869
rect 12685 3903 12743 3909
rect 12685 3869 12697 3903
rect 12731 3900 12743 3903
rect 14525 3903 14583 3909
rect 14525 3900 14537 3903
rect 12731 3872 14537 3900
rect 12731 3869 12743 3872
rect 12685 3863 12743 3869
rect 14525 3869 14537 3872
rect 14571 3869 14583 3903
rect 14525 3863 14583 3869
rect 15077 3903 15135 3909
rect 15077 3869 15089 3903
rect 15123 3900 15135 3903
rect 16917 3903 16975 3909
rect 16917 3900 16929 3903
rect 15123 3872 16929 3900
rect 15123 3869 15135 3872
rect 15077 3863 15135 3869
rect 16917 3869 16929 3872
rect 16963 3869 16975 3903
rect 16917 3863 16975 3869
rect 17469 3903 17527 3909
rect 17469 3869 17481 3903
rect 17515 3900 17527 3903
rect 18496 3900 18524 3940
rect 19309 3937 19321 3940
rect 19355 3937 19367 3971
rect 19309 3931 19367 3937
rect 19861 3971 19919 3977
rect 19861 3937 19873 3971
rect 19907 3968 19919 3971
rect 21701 3971 21759 3977
rect 21701 3968 21713 3971
rect 19907 3940 21713 3968
rect 19907 3937 19919 3940
rect 19861 3931 19919 3937
rect 21701 3937 21713 3940
rect 21747 3937 21759 3971
rect 21701 3931 21759 3937
rect 17515 3872 18524 3900
rect 18665 3903 18723 3909
rect 17515 3869 17527 3872
rect 17469 3863 17527 3869
rect 18665 3869 18677 3903
rect 18711 3900 18723 3903
rect 20505 3903 20563 3909
rect 20505 3900 20517 3903
rect 18711 3872 20517 3900
rect 18711 3869 18723 3872
rect 18665 3863 18723 3869
rect 20505 3869 20517 3872
rect 20551 3869 20563 3903
rect 20505 3863 20563 3869
rect 21057 3903 21115 3909
rect 21057 3869 21069 3903
rect 21103 3900 21115 3903
rect 21606 3900 21612 3912
rect 21103 3872 21612 3900
rect 21103 3869 21115 3872
rect 21057 3863 21115 3869
rect 21606 3860 21612 3872
rect 21664 3860 21670 3912
rect 1904 3674 22236 3696
rect 1904 3622 4446 3674
rect 4498 3622 4510 3674
rect 4562 3622 4574 3674
rect 4626 3622 4638 3674
rect 4690 3622 9774 3674
rect 9826 3622 9838 3674
rect 9890 3622 9902 3674
rect 9954 3622 9966 3674
rect 10018 3622 15102 3674
rect 15154 3622 15166 3674
rect 15218 3622 15230 3674
rect 15282 3622 15294 3674
rect 15346 3622 20430 3674
rect 20482 3622 20494 3674
rect 20546 3622 20558 3674
rect 20610 3622 20622 3674
rect 20674 3622 22236 3674
rect 1904 3600 22236 3622
rect 21606 3452 21612 3504
rect 21664 3492 21670 3504
rect 21701 3495 21759 3501
rect 21701 3492 21713 3495
rect 21664 3464 21713 3492
rect 21664 3452 21670 3464
rect 21701 3461 21713 3464
rect 21747 3461 21759 3495
rect 21701 3455 21759 3461
rect 3117 3427 3175 3433
rect 3117 3393 3129 3427
rect 3163 3424 3175 3427
rect 3850 3424 3856 3436
rect 3163 3396 3856 3424
rect 3163 3393 3175 3396
rect 3117 3387 3175 3393
rect 3850 3384 3856 3396
rect 3908 3384 3914 3436
rect 3761 3359 3819 3365
rect 3761 3325 3773 3359
rect 3807 3356 3819 3359
rect 4313 3359 4371 3365
rect 4313 3356 4325 3359
rect 3807 3328 4325 3356
rect 3807 3325 3819 3328
rect 3761 3319 3819 3325
rect 4313 3325 4325 3328
rect 4359 3325 4371 3359
rect 4313 3319 4371 3325
rect 4957 3359 5015 3365
rect 4957 3325 4969 3359
rect 5003 3356 5015 3359
rect 5509 3359 5567 3365
rect 5509 3356 5521 3359
rect 5003 3328 5521 3356
rect 5003 3325 5015 3328
rect 4957 3319 5015 3325
rect 5509 3325 5521 3328
rect 5555 3325 5567 3359
rect 5509 3319 5567 3325
rect 6153 3359 6211 3365
rect 6153 3325 6165 3359
rect 6199 3356 6211 3359
rect 6705 3359 6763 3365
rect 6705 3356 6717 3359
rect 6199 3328 6717 3356
rect 6199 3325 6211 3328
rect 6153 3319 6211 3325
rect 6705 3325 6717 3328
rect 6751 3325 6763 3359
rect 6705 3319 6763 3325
rect 7349 3359 7407 3365
rect 7349 3325 7361 3359
rect 7395 3356 7407 3359
rect 7901 3359 7959 3365
rect 7901 3356 7913 3359
rect 7395 3328 7913 3356
rect 7395 3325 7407 3328
rect 7349 3319 7407 3325
rect 7901 3325 7913 3328
rect 7947 3325 7959 3359
rect 7901 3319 7959 3325
rect 8545 3359 8603 3365
rect 8545 3325 8557 3359
rect 8591 3356 8603 3359
rect 9097 3359 9155 3365
rect 9097 3356 9109 3359
rect 8591 3328 9109 3356
rect 8591 3325 8603 3328
rect 8545 3319 8603 3325
rect 9097 3325 9109 3328
rect 9143 3325 9155 3359
rect 9097 3319 9155 3325
rect 9741 3359 9799 3365
rect 9741 3325 9753 3359
rect 9787 3356 9799 3359
rect 10293 3359 10351 3365
rect 10293 3356 10305 3359
rect 9787 3328 10305 3356
rect 9787 3325 9799 3328
rect 9741 3319 9799 3325
rect 10293 3325 10305 3328
rect 10339 3325 10351 3359
rect 10293 3319 10351 3325
rect 10937 3359 10995 3365
rect 10937 3325 10949 3359
rect 10983 3356 10995 3359
rect 11489 3359 11547 3365
rect 11489 3356 11501 3359
rect 10983 3328 11501 3356
rect 10983 3325 10995 3328
rect 10937 3319 10995 3325
rect 11489 3325 11501 3328
rect 11535 3325 11547 3359
rect 11489 3319 11547 3325
rect 12133 3359 12191 3365
rect 12133 3325 12145 3359
rect 12179 3356 12191 3359
rect 12685 3359 12743 3365
rect 12685 3356 12697 3359
rect 12179 3328 12697 3356
rect 12179 3325 12191 3328
rect 12133 3319 12191 3325
rect 12685 3325 12697 3328
rect 12731 3325 12743 3359
rect 12685 3319 12743 3325
rect 13329 3359 13387 3365
rect 13329 3325 13341 3359
rect 13375 3356 13387 3359
rect 13881 3359 13939 3365
rect 13881 3356 13893 3359
rect 13375 3328 13893 3356
rect 13375 3325 13387 3328
rect 13329 3319 13387 3325
rect 13881 3325 13893 3328
rect 13927 3325 13939 3359
rect 13881 3319 13939 3325
rect 14525 3359 14583 3365
rect 14525 3325 14537 3359
rect 14571 3356 14583 3359
rect 15077 3359 15135 3365
rect 15077 3356 15089 3359
rect 14571 3328 15089 3356
rect 14571 3325 14583 3328
rect 14525 3319 14583 3325
rect 15077 3325 15089 3328
rect 15123 3325 15135 3359
rect 15077 3319 15135 3325
rect 15721 3359 15779 3365
rect 15721 3325 15733 3359
rect 15767 3356 15779 3359
rect 16273 3359 16331 3365
rect 16273 3356 16285 3359
rect 15767 3328 16285 3356
rect 15767 3325 15779 3328
rect 15721 3319 15779 3325
rect 16273 3325 16285 3328
rect 16319 3325 16331 3359
rect 16273 3319 16331 3325
rect 16917 3359 16975 3365
rect 16917 3325 16929 3359
rect 16963 3356 16975 3359
rect 17469 3359 17527 3365
rect 17469 3356 17481 3359
rect 16963 3328 17481 3356
rect 16963 3325 16975 3328
rect 16917 3319 16975 3325
rect 17469 3325 17481 3328
rect 17515 3325 17527 3359
rect 17469 3319 17527 3325
rect 18113 3359 18171 3365
rect 18113 3325 18125 3359
rect 18159 3356 18171 3359
rect 18665 3359 18723 3365
rect 18665 3356 18677 3359
rect 18159 3328 18677 3356
rect 18159 3325 18171 3328
rect 18113 3319 18171 3325
rect 18665 3325 18677 3328
rect 18711 3325 18723 3359
rect 18665 3319 18723 3325
rect 19309 3359 19367 3365
rect 19309 3325 19321 3359
rect 19355 3356 19367 3359
rect 19861 3359 19919 3365
rect 19861 3356 19873 3359
rect 19355 3328 19873 3356
rect 19355 3325 19367 3328
rect 19309 3319 19367 3325
rect 19861 3325 19873 3328
rect 19907 3325 19919 3359
rect 19861 3319 19919 3325
rect 20505 3359 20563 3365
rect 20505 3325 20517 3359
rect 20551 3356 20563 3359
rect 21057 3359 21115 3365
rect 21057 3356 21069 3359
rect 20551 3328 21069 3356
rect 20551 3325 20563 3328
rect 20505 3319 20563 3325
rect 21057 3325 21069 3328
rect 21103 3325 21115 3359
rect 21057 3319 21115 3325
rect 1904 3130 22236 3152
rect 1904 3078 7110 3130
rect 7162 3078 7174 3130
rect 7226 3078 7238 3130
rect 7290 3078 7302 3130
rect 7354 3078 12438 3130
rect 12490 3078 12502 3130
rect 12554 3078 12566 3130
rect 12618 3078 12630 3130
rect 12682 3078 17766 3130
rect 17818 3078 17830 3130
rect 17882 3078 17894 3130
rect 17946 3078 17958 3130
rect 18010 3078 22236 3130
rect 1904 3056 22236 3078
rect 3761 3019 3819 3025
rect 3761 2985 3773 3019
rect 3807 3016 3819 3019
rect 3850 3016 3856 3028
rect 3807 2988 3856 3016
rect 3807 2985 3819 2988
rect 3761 2979 3819 2985
rect 3850 2976 3856 2988
rect 3908 2976 3914 3028
rect 4313 2883 4371 2889
rect 4313 2849 4325 2883
rect 4359 2880 4371 2883
rect 6153 2883 6211 2889
rect 6153 2880 6165 2883
rect 4359 2852 6165 2880
rect 4359 2849 4371 2852
rect 4313 2843 4371 2849
rect 6153 2849 6165 2852
rect 6199 2849 6211 2883
rect 6153 2843 6211 2849
rect 7901 2883 7959 2889
rect 7901 2849 7913 2883
rect 7947 2880 7959 2883
rect 9741 2883 9799 2889
rect 9741 2880 9753 2883
rect 7947 2852 9753 2880
rect 7947 2849 7959 2852
rect 7901 2843 7959 2849
rect 9741 2849 9753 2852
rect 9787 2849 9799 2883
rect 9741 2843 9799 2849
rect 11489 2883 11547 2889
rect 11489 2849 11501 2883
rect 11535 2880 11547 2883
rect 13329 2883 13387 2889
rect 13329 2880 13341 2883
rect 11535 2852 13341 2880
rect 11535 2849 11547 2852
rect 11489 2843 11547 2849
rect 13329 2849 13341 2852
rect 13375 2849 13387 2883
rect 13329 2843 13387 2849
rect 13881 2883 13939 2889
rect 13881 2849 13893 2883
rect 13927 2880 13939 2883
rect 15721 2883 15779 2889
rect 15721 2880 15733 2883
rect 13927 2852 15733 2880
rect 13927 2849 13939 2852
rect 13881 2843 13939 2849
rect 15721 2849 15733 2852
rect 15767 2849 15779 2883
rect 15721 2843 15779 2849
rect 16273 2883 16331 2889
rect 16273 2849 16285 2883
rect 16319 2880 16331 2883
rect 17006 2880 17012 2892
rect 16319 2852 17012 2880
rect 16319 2849 16331 2852
rect 16273 2843 16331 2849
rect 17006 2840 17012 2852
rect 17064 2840 17070 2892
rect 17469 2883 17527 2889
rect 17469 2849 17481 2883
rect 17515 2880 17527 2883
rect 19309 2883 19367 2889
rect 19309 2880 19321 2883
rect 17515 2852 19321 2880
rect 17515 2849 17527 2852
rect 17469 2843 17527 2849
rect 19309 2849 19321 2852
rect 19355 2849 19367 2883
rect 19309 2843 19367 2849
rect 19861 2883 19919 2889
rect 19861 2849 19873 2883
rect 19907 2880 19919 2883
rect 21701 2883 21759 2889
rect 21701 2880 21713 2883
rect 19907 2852 21713 2880
rect 19907 2849 19919 2852
rect 19861 2843 19919 2849
rect 21701 2849 21713 2852
rect 21747 2849 21759 2883
rect 21701 2843 21759 2849
rect 3117 2815 3175 2821
rect 3117 2781 3129 2815
rect 3163 2812 3175 2815
rect 5509 2815 5567 2821
rect 3163 2784 4080 2812
rect 3163 2781 3175 2784
rect 3117 2775 3175 2781
rect 4052 2744 4080 2784
rect 5509 2781 5521 2815
rect 5555 2812 5567 2815
rect 6705 2815 6763 2821
rect 5555 2784 6472 2812
rect 5555 2781 5567 2784
rect 5509 2775 5567 2781
rect 4957 2747 5015 2753
rect 4957 2744 4969 2747
rect 4052 2716 4969 2744
rect 4957 2713 4969 2716
rect 5003 2713 5015 2747
rect 6444 2744 6472 2784
rect 6705 2781 6717 2815
rect 6751 2812 6763 2815
rect 9097 2815 9155 2821
rect 6751 2784 7668 2812
rect 6751 2781 6763 2784
rect 6705 2775 6763 2781
rect 7349 2747 7407 2753
rect 7349 2744 7361 2747
rect 6444 2716 7361 2744
rect 4957 2707 5015 2713
rect 7349 2713 7361 2716
rect 7395 2713 7407 2747
rect 7640 2744 7668 2784
rect 9097 2781 9109 2815
rect 9143 2812 9155 2815
rect 9646 2812 9652 2824
rect 9143 2784 9652 2812
rect 9143 2781 9155 2784
rect 9097 2775 9155 2781
rect 9646 2772 9652 2784
rect 9704 2772 9710 2824
rect 10293 2815 10351 2821
rect 10293 2781 10305 2815
rect 10339 2812 10351 2815
rect 12133 2815 12191 2821
rect 12133 2812 12145 2815
rect 10339 2784 12145 2812
rect 10339 2781 10351 2784
rect 10293 2775 10351 2781
rect 12133 2781 12145 2784
rect 12179 2781 12191 2815
rect 12133 2775 12191 2781
rect 12685 2815 12743 2821
rect 12685 2781 12697 2815
rect 12731 2812 12743 2815
rect 15077 2815 15135 2821
rect 12731 2784 13648 2812
rect 12731 2781 12743 2784
rect 12685 2775 12743 2781
rect 8545 2747 8603 2753
rect 8545 2744 8557 2747
rect 7640 2716 8557 2744
rect 7349 2707 7407 2713
rect 8545 2713 8557 2716
rect 8591 2713 8603 2747
rect 13620 2744 13648 2784
rect 15077 2781 15089 2815
rect 15123 2812 15135 2815
rect 18665 2815 18723 2821
rect 15123 2784 16040 2812
rect 15123 2781 15135 2784
rect 15077 2775 15135 2781
rect 14525 2747 14583 2753
rect 14525 2744 14537 2747
rect 13620 2716 14537 2744
rect 8545 2707 8603 2713
rect 14525 2713 14537 2716
rect 14571 2713 14583 2747
rect 16012 2744 16040 2784
rect 18665 2781 18677 2815
rect 18711 2812 18723 2815
rect 21057 2815 21115 2821
rect 18711 2784 19628 2812
rect 18711 2781 18723 2784
rect 18665 2775 18723 2781
rect 16917 2747 16975 2753
rect 16917 2744 16929 2747
rect 16012 2716 16929 2744
rect 14525 2707 14583 2713
rect 16917 2713 16929 2716
rect 16963 2713 16975 2747
rect 16917 2707 16975 2713
rect 17006 2704 17012 2756
rect 17064 2744 17070 2756
rect 18113 2747 18171 2753
rect 18113 2744 18125 2747
rect 17064 2716 18125 2744
rect 17064 2704 17070 2716
rect 18113 2713 18125 2716
rect 18159 2713 18171 2747
rect 19600 2744 19628 2784
rect 21057 2781 21069 2815
rect 21103 2812 21115 2815
rect 21606 2812 21612 2824
rect 21103 2784 21612 2812
rect 21103 2781 21115 2784
rect 21057 2775 21115 2781
rect 21606 2772 21612 2784
rect 21664 2772 21670 2824
rect 20505 2747 20563 2753
rect 20505 2744 20517 2747
rect 19600 2716 20517 2744
rect 18113 2707 18171 2713
rect 20505 2713 20517 2716
rect 20551 2713 20563 2747
rect 20505 2707 20563 2713
rect 9646 2636 9652 2688
rect 9704 2676 9710 2688
rect 10937 2679 10995 2685
rect 10937 2676 10949 2679
rect 9704 2648 10949 2676
rect 9704 2636 9710 2648
rect 10937 2645 10949 2648
rect 10983 2645 10995 2679
rect 10937 2639 10995 2645
rect 1904 2586 22236 2608
rect 1904 2534 4446 2586
rect 4498 2534 4510 2586
rect 4562 2534 4574 2586
rect 4626 2534 4638 2586
rect 4690 2534 9774 2586
rect 9826 2534 9838 2586
rect 9890 2534 9902 2586
rect 9954 2534 9966 2586
rect 10018 2534 15102 2586
rect 15154 2534 15166 2586
rect 15218 2534 15230 2586
rect 15282 2534 15294 2586
rect 15346 2534 20430 2586
rect 20482 2534 20494 2586
rect 20546 2534 20558 2586
rect 20610 2534 20622 2586
rect 20674 2534 22236 2586
rect 1904 2512 22236 2534
rect 21606 2432 21612 2484
rect 21664 2472 21670 2484
rect 21701 2475 21759 2481
rect 21701 2472 21713 2475
rect 21664 2444 21713 2472
rect 21664 2432 21670 2444
rect 21701 2441 21713 2444
rect 21747 2441 21759 2475
rect 21701 2435 21759 2441
rect 3117 2339 3175 2345
rect 3117 2305 3129 2339
rect 3163 2336 3175 2339
rect 3850 2336 3856 2348
rect 3163 2308 3856 2336
rect 3163 2305 3175 2308
rect 3117 2299 3175 2305
rect 3850 2296 3856 2308
rect 3908 2296 3914 2348
rect 3761 2271 3819 2277
rect 3761 2237 3773 2271
rect 3807 2268 3819 2271
rect 4313 2271 4371 2277
rect 4313 2268 4325 2271
rect 3807 2240 4325 2268
rect 3807 2237 3819 2240
rect 3761 2231 3819 2237
rect 4313 2237 4325 2240
rect 4359 2237 4371 2271
rect 4313 2231 4371 2237
rect 4957 2271 5015 2277
rect 4957 2237 4969 2271
rect 5003 2268 5015 2271
rect 5509 2271 5567 2277
rect 5509 2268 5521 2271
rect 5003 2240 5521 2268
rect 5003 2237 5015 2240
rect 4957 2231 5015 2237
rect 5509 2237 5521 2240
rect 5555 2237 5567 2271
rect 5509 2231 5567 2237
rect 6153 2271 6211 2277
rect 6153 2237 6165 2271
rect 6199 2268 6211 2271
rect 6705 2271 6763 2277
rect 6705 2268 6717 2271
rect 6199 2240 6717 2268
rect 6199 2237 6211 2240
rect 6153 2231 6211 2237
rect 6705 2237 6717 2240
rect 6751 2237 6763 2271
rect 6705 2231 6763 2237
rect 7349 2271 7407 2277
rect 7349 2237 7361 2271
rect 7395 2268 7407 2271
rect 7901 2271 7959 2277
rect 7901 2268 7913 2271
rect 7395 2240 7913 2268
rect 7395 2237 7407 2240
rect 7349 2231 7407 2237
rect 7901 2237 7913 2240
rect 7947 2237 7959 2271
rect 7901 2231 7959 2237
rect 8545 2271 8603 2277
rect 8545 2237 8557 2271
rect 8591 2268 8603 2271
rect 9097 2271 9155 2277
rect 9097 2268 9109 2271
rect 8591 2240 9109 2268
rect 8591 2237 8603 2240
rect 8545 2231 8603 2237
rect 9097 2237 9109 2240
rect 9143 2237 9155 2271
rect 9097 2231 9155 2237
rect 9741 2271 9799 2277
rect 9741 2237 9753 2271
rect 9787 2268 9799 2271
rect 10293 2271 10351 2277
rect 10293 2268 10305 2271
rect 9787 2240 10305 2268
rect 9787 2237 9799 2240
rect 9741 2231 9799 2237
rect 10293 2237 10305 2240
rect 10339 2237 10351 2271
rect 10293 2231 10351 2237
rect 10937 2271 10995 2277
rect 10937 2237 10949 2271
rect 10983 2268 10995 2271
rect 11489 2271 11547 2277
rect 11489 2268 11501 2271
rect 10983 2240 11501 2268
rect 10983 2237 10995 2240
rect 10937 2231 10995 2237
rect 11489 2237 11501 2240
rect 11535 2237 11547 2271
rect 11489 2231 11547 2237
rect 12133 2271 12191 2277
rect 12133 2237 12145 2271
rect 12179 2268 12191 2271
rect 12685 2271 12743 2277
rect 12685 2268 12697 2271
rect 12179 2240 12697 2268
rect 12179 2237 12191 2240
rect 12133 2231 12191 2237
rect 12685 2237 12697 2240
rect 12731 2237 12743 2271
rect 12685 2231 12743 2237
rect 13329 2271 13387 2277
rect 13329 2237 13341 2271
rect 13375 2268 13387 2271
rect 13881 2271 13939 2277
rect 13881 2268 13893 2271
rect 13375 2240 13893 2268
rect 13375 2237 13387 2240
rect 13329 2231 13387 2237
rect 13881 2237 13893 2240
rect 13927 2237 13939 2271
rect 13881 2231 13939 2237
rect 14525 2271 14583 2277
rect 14525 2237 14537 2271
rect 14571 2268 14583 2271
rect 15077 2271 15135 2277
rect 15077 2268 15089 2271
rect 14571 2240 15089 2268
rect 14571 2237 14583 2240
rect 14525 2231 14583 2237
rect 15077 2237 15089 2240
rect 15123 2237 15135 2271
rect 15077 2231 15135 2237
rect 15721 2271 15779 2277
rect 15721 2237 15733 2271
rect 15767 2268 15779 2271
rect 16273 2271 16331 2277
rect 16273 2268 16285 2271
rect 15767 2240 16285 2268
rect 15767 2237 15779 2240
rect 15721 2231 15779 2237
rect 16273 2237 16285 2240
rect 16319 2237 16331 2271
rect 16273 2231 16331 2237
rect 16917 2271 16975 2277
rect 16917 2237 16929 2271
rect 16963 2268 16975 2271
rect 17469 2271 17527 2277
rect 17469 2268 17481 2271
rect 16963 2240 17481 2268
rect 16963 2237 16975 2240
rect 16917 2231 16975 2237
rect 17469 2237 17481 2240
rect 17515 2237 17527 2271
rect 17469 2231 17527 2237
rect 18113 2271 18171 2277
rect 18113 2237 18125 2271
rect 18159 2268 18171 2271
rect 18665 2271 18723 2277
rect 18665 2268 18677 2271
rect 18159 2240 18677 2268
rect 18159 2237 18171 2240
rect 18113 2231 18171 2237
rect 18665 2237 18677 2240
rect 18711 2237 18723 2271
rect 18665 2231 18723 2237
rect 19309 2271 19367 2277
rect 19309 2237 19321 2271
rect 19355 2268 19367 2271
rect 19861 2271 19919 2277
rect 19861 2268 19873 2271
rect 19355 2240 19873 2268
rect 19355 2237 19367 2240
rect 19309 2231 19367 2237
rect 19861 2237 19873 2240
rect 19907 2237 19919 2271
rect 19861 2231 19919 2237
rect 20505 2271 20563 2277
rect 20505 2237 20517 2271
rect 20551 2268 20563 2271
rect 21057 2271 21115 2277
rect 21057 2268 21069 2271
rect 20551 2240 21069 2268
rect 20551 2237 20563 2240
rect 20505 2231 20563 2237
rect 21057 2237 21069 2240
rect 21103 2237 21115 2271
rect 21057 2231 21115 2237
rect 1904 2042 22236 2064
rect 1904 1990 7110 2042
rect 7162 1990 7174 2042
rect 7226 1990 7238 2042
rect 7290 1990 7302 2042
rect 7354 1990 12438 2042
rect 12490 1990 12502 2042
rect 12554 1990 12566 2042
rect 12618 1990 12630 2042
rect 12682 1990 17766 2042
rect 17818 1990 17830 2042
rect 17882 1990 17894 2042
rect 17946 1990 17958 2042
rect 18010 1990 22236 2042
rect 1904 1968 22236 1990
rect 3761 1931 3819 1937
rect 3761 1897 3773 1931
rect 3807 1928 3819 1931
rect 3850 1928 3856 1940
rect 3807 1900 3856 1928
rect 3807 1897 3819 1900
rect 3761 1891 3819 1897
rect 3850 1888 3856 1900
rect 3908 1888 3914 1940
rect 3117 1795 3175 1801
rect 3117 1761 3129 1795
rect 3163 1792 3175 1795
rect 4957 1795 5015 1801
rect 4957 1792 4969 1795
rect 3163 1764 4969 1792
rect 3163 1761 3175 1764
rect 3117 1755 3175 1761
rect 4957 1761 4969 1764
rect 5003 1761 5015 1795
rect 4957 1755 5015 1761
rect 5509 1795 5567 1801
rect 5509 1761 5521 1795
rect 5555 1792 5567 1795
rect 7349 1795 7407 1801
rect 7349 1792 7361 1795
rect 5555 1764 7361 1792
rect 5555 1761 5567 1764
rect 5509 1755 5567 1761
rect 7349 1761 7361 1764
rect 7395 1761 7407 1795
rect 7349 1755 7407 1761
rect 7901 1795 7959 1801
rect 7901 1761 7913 1795
rect 7947 1792 7959 1795
rect 9097 1795 9155 1801
rect 7947 1764 8772 1792
rect 7947 1761 7959 1764
rect 7901 1755 7959 1761
rect 4313 1727 4371 1733
rect 4313 1693 4325 1727
rect 4359 1724 4371 1727
rect 6153 1727 6211 1733
rect 6153 1724 6165 1727
rect 4359 1696 6165 1724
rect 4359 1693 4371 1696
rect 4313 1687 4371 1693
rect 6153 1693 6165 1696
rect 6199 1693 6211 1727
rect 6153 1687 6211 1693
rect 6705 1727 6763 1733
rect 6705 1693 6717 1727
rect 6751 1724 6763 1727
rect 8545 1727 8603 1733
rect 8545 1724 8557 1727
rect 6751 1696 8557 1724
rect 6751 1693 6763 1696
rect 6705 1687 6763 1693
rect 8545 1693 8557 1696
rect 8591 1693 8603 1727
rect 8744 1724 8772 1764
rect 9097 1761 9109 1795
rect 9143 1792 9155 1795
rect 10937 1795 10995 1801
rect 10937 1792 10949 1795
rect 9143 1764 10949 1792
rect 9143 1761 9155 1764
rect 9097 1755 9155 1761
rect 10937 1761 10949 1764
rect 10983 1761 10995 1795
rect 10937 1755 10995 1761
rect 11489 1795 11547 1801
rect 11489 1761 11501 1795
rect 11535 1792 11547 1795
rect 13329 1795 13387 1801
rect 13329 1792 13341 1795
rect 11535 1764 13341 1792
rect 11535 1761 11547 1764
rect 11489 1755 11547 1761
rect 13329 1761 13341 1764
rect 13375 1761 13387 1795
rect 13329 1755 13387 1761
rect 13881 1795 13939 1801
rect 13881 1761 13893 1795
rect 13927 1792 13939 1795
rect 15721 1795 15779 1801
rect 15721 1792 15733 1795
rect 13927 1764 15733 1792
rect 13927 1761 13939 1764
rect 13881 1755 13939 1761
rect 15721 1761 15733 1764
rect 15767 1761 15779 1795
rect 15721 1755 15779 1761
rect 16273 1795 16331 1801
rect 16273 1761 16285 1795
rect 16319 1792 16331 1795
rect 18113 1795 18171 1801
rect 18113 1792 18125 1795
rect 16319 1764 18125 1792
rect 16319 1761 16331 1764
rect 16273 1755 16331 1761
rect 18113 1761 18125 1764
rect 18159 1761 18171 1795
rect 19309 1795 19367 1801
rect 19309 1792 19321 1795
rect 18113 1755 18171 1761
rect 18496 1764 19321 1792
rect 9741 1727 9799 1733
rect 9741 1724 9753 1727
rect 8744 1696 9753 1724
rect 8545 1687 8603 1693
rect 9741 1693 9753 1696
rect 9787 1693 9799 1727
rect 9741 1687 9799 1693
rect 10293 1727 10351 1733
rect 10293 1693 10305 1727
rect 10339 1724 10351 1727
rect 12133 1727 12191 1733
rect 12133 1724 12145 1727
rect 10339 1696 12145 1724
rect 10339 1693 10351 1696
rect 10293 1687 10351 1693
rect 12133 1693 12145 1696
rect 12179 1693 12191 1727
rect 12133 1687 12191 1693
rect 12685 1727 12743 1733
rect 12685 1693 12697 1727
rect 12731 1724 12743 1727
rect 14525 1727 14583 1733
rect 14525 1724 14537 1727
rect 12731 1696 14537 1724
rect 12731 1693 12743 1696
rect 12685 1687 12743 1693
rect 14525 1693 14537 1696
rect 14571 1693 14583 1727
rect 14525 1687 14583 1693
rect 15077 1727 15135 1733
rect 15077 1693 15089 1727
rect 15123 1724 15135 1727
rect 16917 1727 16975 1733
rect 16917 1724 16929 1727
rect 15123 1696 16929 1724
rect 15123 1693 15135 1696
rect 15077 1687 15135 1693
rect 16917 1693 16929 1696
rect 16963 1693 16975 1727
rect 16917 1687 16975 1693
rect 17469 1727 17527 1733
rect 17469 1693 17481 1727
rect 17515 1724 17527 1727
rect 18496 1724 18524 1764
rect 19309 1761 19321 1764
rect 19355 1761 19367 1795
rect 19309 1755 19367 1761
rect 19861 1795 19919 1801
rect 19861 1761 19873 1795
rect 19907 1792 19919 1795
rect 21701 1795 21759 1801
rect 21701 1792 21713 1795
rect 19907 1764 21713 1792
rect 19907 1761 19919 1764
rect 19861 1755 19919 1761
rect 21701 1761 21713 1764
rect 21747 1761 21759 1795
rect 21701 1755 21759 1761
rect 17515 1696 18524 1724
rect 18665 1727 18723 1733
rect 17515 1693 17527 1696
rect 17469 1687 17527 1693
rect 18665 1693 18677 1727
rect 18711 1724 18723 1727
rect 20505 1727 20563 1733
rect 20505 1724 20517 1727
rect 18711 1696 20517 1724
rect 18711 1693 18723 1696
rect 18665 1687 18723 1693
rect 20505 1693 20517 1696
rect 20551 1693 20563 1727
rect 20505 1687 20563 1693
rect 21057 1727 21115 1733
rect 21057 1693 21069 1727
rect 21103 1724 21115 1727
rect 21606 1724 21612 1736
rect 21103 1696 21612 1724
rect 21103 1693 21115 1696
rect 21057 1687 21115 1693
rect 21606 1684 21612 1696
rect 21664 1684 21670 1736
rect 1904 1498 22236 1520
rect 1904 1446 4446 1498
rect 4498 1446 4510 1498
rect 4562 1446 4574 1498
rect 4626 1446 4638 1498
rect 4690 1446 9774 1498
rect 9826 1446 9838 1498
rect 9890 1446 9902 1498
rect 9954 1446 9966 1498
rect 10018 1446 15102 1498
rect 15154 1446 15166 1498
rect 15218 1446 15230 1498
rect 15282 1446 15294 1498
rect 15346 1446 20430 1498
rect 20482 1446 20494 1498
rect 20546 1446 20558 1498
rect 20610 1446 20622 1498
rect 20674 1446 22236 1498
rect 1904 1424 22236 1446
rect 21606 1276 21612 1328
rect 21664 1316 21670 1328
rect 21701 1319 21759 1325
rect 21701 1316 21713 1319
rect 21664 1288 21713 1316
rect 21664 1276 21670 1288
rect 21701 1285 21713 1288
rect 21747 1285 21759 1319
rect 21701 1279 21759 1285
rect 2930 1140 2936 1192
rect 2988 1180 2994 1192
rect 3117 1183 3175 1189
rect 3117 1180 3129 1183
rect 2988 1152 3129 1180
rect 2988 1140 2994 1152
rect 3117 1149 3129 1152
rect 3163 1149 3175 1183
rect 3117 1143 3175 1149
rect 3761 1183 3819 1189
rect 3761 1149 3773 1183
rect 3807 1180 3819 1183
rect 4313 1183 4371 1189
rect 4313 1180 4325 1183
rect 3807 1152 4325 1180
rect 3807 1149 3819 1152
rect 3761 1143 3819 1149
rect 4313 1149 4325 1152
rect 4359 1149 4371 1183
rect 4313 1143 4371 1149
rect 4957 1183 5015 1189
rect 4957 1149 4969 1183
rect 5003 1180 5015 1183
rect 5509 1183 5567 1189
rect 5509 1180 5521 1183
rect 5003 1152 5521 1180
rect 5003 1149 5015 1152
rect 4957 1143 5015 1149
rect 5509 1149 5521 1152
rect 5555 1149 5567 1183
rect 5509 1143 5567 1149
rect 6153 1183 6211 1189
rect 6153 1149 6165 1183
rect 6199 1180 6211 1183
rect 6705 1183 6763 1189
rect 6705 1180 6717 1183
rect 6199 1152 6717 1180
rect 6199 1149 6211 1152
rect 6153 1143 6211 1149
rect 6705 1149 6717 1152
rect 6751 1149 6763 1183
rect 6705 1143 6763 1149
rect 7349 1183 7407 1189
rect 7349 1149 7361 1183
rect 7395 1180 7407 1183
rect 7901 1183 7959 1189
rect 7901 1180 7913 1183
rect 7395 1152 7913 1180
rect 7395 1149 7407 1152
rect 7349 1143 7407 1149
rect 7901 1149 7913 1152
rect 7947 1149 7959 1183
rect 7901 1143 7959 1149
rect 8545 1183 8603 1189
rect 8545 1149 8557 1183
rect 8591 1180 8603 1183
rect 9097 1183 9155 1189
rect 9097 1180 9109 1183
rect 8591 1152 9109 1180
rect 8591 1149 8603 1152
rect 8545 1143 8603 1149
rect 9097 1149 9109 1152
rect 9143 1149 9155 1183
rect 9097 1143 9155 1149
rect 9741 1183 9799 1189
rect 9741 1149 9753 1183
rect 9787 1180 9799 1183
rect 10293 1183 10351 1189
rect 10293 1180 10305 1183
rect 9787 1152 10305 1180
rect 9787 1149 9799 1152
rect 9741 1143 9799 1149
rect 10293 1149 10305 1152
rect 10339 1149 10351 1183
rect 10293 1143 10351 1149
rect 10937 1183 10995 1189
rect 10937 1149 10949 1183
rect 10983 1180 10995 1183
rect 11489 1183 11547 1189
rect 11489 1180 11501 1183
rect 10983 1152 11501 1180
rect 10983 1149 10995 1152
rect 10937 1143 10995 1149
rect 11489 1149 11501 1152
rect 11535 1149 11547 1183
rect 11489 1143 11547 1149
rect 12133 1183 12191 1189
rect 12133 1149 12145 1183
rect 12179 1180 12191 1183
rect 12685 1183 12743 1189
rect 12685 1180 12697 1183
rect 12179 1152 12697 1180
rect 12179 1149 12191 1152
rect 12133 1143 12191 1149
rect 12685 1149 12697 1152
rect 12731 1149 12743 1183
rect 12685 1143 12743 1149
rect 13329 1183 13387 1189
rect 13329 1149 13341 1183
rect 13375 1180 13387 1183
rect 13881 1183 13939 1189
rect 13881 1180 13893 1183
rect 13375 1152 13893 1180
rect 13375 1149 13387 1152
rect 13329 1143 13387 1149
rect 13881 1149 13893 1152
rect 13927 1149 13939 1183
rect 13881 1143 13939 1149
rect 14525 1183 14583 1189
rect 14525 1149 14537 1183
rect 14571 1180 14583 1183
rect 15077 1183 15135 1189
rect 15077 1180 15089 1183
rect 14571 1152 15089 1180
rect 14571 1149 14583 1152
rect 14525 1143 14583 1149
rect 15077 1149 15089 1152
rect 15123 1149 15135 1183
rect 15077 1143 15135 1149
rect 15721 1183 15779 1189
rect 15721 1149 15733 1183
rect 15767 1180 15779 1183
rect 16273 1183 16331 1189
rect 16273 1180 16285 1183
rect 15767 1152 16285 1180
rect 15767 1149 15779 1152
rect 15721 1143 15779 1149
rect 16273 1149 16285 1152
rect 16319 1149 16331 1183
rect 16273 1143 16331 1149
rect 16917 1183 16975 1189
rect 16917 1149 16929 1183
rect 16963 1180 16975 1183
rect 17469 1183 17527 1189
rect 17469 1180 17481 1183
rect 16963 1152 17481 1180
rect 16963 1149 16975 1152
rect 16917 1143 16975 1149
rect 17469 1149 17481 1152
rect 17515 1149 17527 1183
rect 17469 1143 17527 1149
rect 18113 1183 18171 1189
rect 18113 1149 18125 1183
rect 18159 1180 18171 1183
rect 18665 1183 18723 1189
rect 18665 1180 18677 1183
rect 18159 1152 18677 1180
rect 18159 1149 18171 1152
rect 18113 1143 18171 1149
rect 18665 1149 18677 1152
rect 18711 1149 18723 1183
rect 18665 1143 18723 1149
rect 19309 1183 19367 1189
rect 19309 1149 19321 1183
rect 19355 1180 19367 1183
rect 19861 1183 19919 1189
rect 19861 1180 19873 1183
rect 19355 1152 19873 1180
rect 19355 1149 19367 1152
rect 19309 1143 19367 1149
rect 19861 1149 19873 1152
rect 19907 1149 19919 1183
rect 19861 1143 19919 1149
rect 20505 1183 20563 1189
rect 20505 1149 20517 1183
rect 20551 1180 20563 1183
rect 21057 1183 21115 1189
rect 21057 1180 21069 1183
rect 20551 1152 21069 1180
rect 20551 1149 20563 1152
rect 20505 1143 20563 1149
rect 21057 1149 21069 1152
rect 21103 1149 21115 1183
rect 21057 1143 21115 1149
rect 1904 954 22236 976
rect 1904 902 7110 954
rect 7162 902 7174 954
rect 7226 902 7238 954
rect 7290 902 7302 954
rect 7354 902 12438 954
rect 12490 902 12502 954
rect 12554 902 12566 954
rect 12618 902 12630 954
rect 12682 902 17766 954
rect 17818 902 17830 954
rect 17882 902 17894 954
rect 17946 902 17958 954
rect 18010 902 22236 954
rect 1904 880 22236 902
<< via1 >>
rect 4446 22118 4498 22170
rect 4510 22118 4562 22170
rect 4574 22118 4626 22170
rect 4638 22118 4690 22170
rect 9774 22118 9826 22170
rect 9838 22118 9890 22170
rect 9902 22118 9954 22170
rect 9966 22118 10018 22170
rect 15102 22118 15154 22170
rect 15166 22118 15218 22170
rect 15230 22118 15282 22170
rect 15294 22118 15346 22170
rect 20430 22118 20482 22170
rect 20494 22118 20546 22170
rect 20558 22118 20610 22170
rect 20622 22118 20674 22170
rect 1924 22059 1976 22068
rect 1924 22025 1933 22059
rect 1933 22025 1967 22059
rect 1967 22025 1976 22059
rect 1924 22016 1976 22025
rect 2292 21991 2344 22000
rect 2292 21957 2301 21991
rect 2301 21957 2335 21991
rect 2335 21957 2344 21991
rect 2292 21948 2344 21957
rect 2476 21855 2528 21864
rect 2476 21821 2485 21855
rect 2485 21821 2519 21855
rect 2519 21821 2528 21855
rect 2476 21812 2528 21821
rect 2292 21744 2344 21796
rect 7110 21574 7162 21626
rect 7174 21574 7226 21626
rect 7238 21574 7290 21626
rect 7302 21574 7354 21626
rect 12438 21574 12490 21626
rect 12502 21574 12554 21626
rect 12566 21574 12618 21626
rect 12630 21574 12682 21626
rect 17766 21574 17818 21626
rect 17830 21574 17882 21626
rect 17894 21574 17946 21626
rect 17958 21574 18010 21626
rect 2292 21472 2344 21524
rect 2476 21379 2528 21388
rect 2476 21345 2485 21379
rect 2485 21345 2519 21379
rect 2519 21345 2528 21379
rect 2476 21336 2528 21345
rect 3764 21336 3816 21388
rect 2292 21175 2344 21184
rect 2292 21141 2301 21175
rect 2301 21141 2335 21175
rect 2335 21141 2344 21175
rect 2292 21132 2344 21141
rect 4446 21030 4498 21082
rect 4510 21030 4562 21082
rect 4574 21030 4626 21082
rect 4638 21030 4690 21082
rect 9774 21030 9826 21082
rect 9838 21030 9890 21082
rect 9902 21030 9954 21082
rect 9966 21030 10018 21082
rect 15102 21030 15154 21082
rect 15166 21030 15218 21082
rect 15230 21030 15282 21082
rect 15294 21030 15346 21082
rect 20430 21030 20482 21082
rect 20494 21030 20546 21082
rect 20558 21030 20610 21082
rect 20622 21030 20674 21082
rect 3764 20971 3816 20980
rect 3764 20937 3773 20971
rect 3773 20937 3807 20971
rect 3807 20937 3816 20971
rect 3764 20928 3816 20937
rect 2292 20724 2344 20776
rect 7110 20486 7162 20538
rect 7174 20486 7226 20538
rect 7238 20486 7290 20538
rect 7302 20486 7354 20538
rect 12438 20486 12490 20538
rect 12502 20486 12554 20538
rect 12566 20486 12618 20538
rect 12630 20486 12682 20538
rect 17766 20486 17818 20538
rect 17830 20486 17882 20538
rect 17894 20486 17946 20538
rect 17958 20486 18010 20538
rect 2292 20384 2344 20436
rect 2476 20291 2528 20300
rect 2476 20257 2485 20291
rect 2485 20257 2519 20291
rect 2519 20257 2528 20291
rect 2476 20248 2528 20257
rect 4316 20223 4368 20232
rect 4316 20189 4325 20223
rect 4325 20189 4359 20223
rect 4359 20189 4368 20223
rect 4316 20180 4368 20189
rect 2292 20087 2344 20096
rect 2292 20053 2301 20087
rect 2301 20053 2335 20087
rect 2335 20053 2344 20087
rect 2292 20044 2344 20053
rect 4446 19942 4498 19994
rect 4510 19942 4562 19994
rect 4574 19942 4626 19994
rect 4638 19942 4690 19994
rect 9774 19942 9826 19994
rect 9838 19942 9890 19994
rect 9902 19942 9954 19994
rect 9966 19942 10018 19994
rect 15102 19942 15154 19994
rect 15166 19942 15218 19994
rect 15230 19942 15282 19994
rect 15294 19942 15346 19994
rect 20430 19942 20482 19994
rect 20494 19942 20546 19994
rect 20558 19942 20610 19994
rect 20622 19942 20674 19994
rect 4316 19840 4368 19892
rect 2292 19636 2344 19688
rect 7110 19398 7162 19450
rect 7174 19398 7226 19450
rect 7238 19398 7290 19450
rect 7302 19398 7354 19450
rect 12438 19398 12490 19450
rect 12502 19398 12554 19450
rect 12566 19398 12618 19450
rect 12630 19398 12682 19450
rect 17766 19398 17818 19450
rect 17830 19398 17882 19450
rect 17894 19398 17946 19450
rect 17958 19398 18010 19450
rect 2292 19296 2344 19348
rect 2476 19203 2528 19212
rect 2476 19169 2485 19203
rect 2485 19169 2519 19203
rect 2519 19169 2528 19203
rect 2476 19160 2528 19169
rect 6708 19135 6760 19144
rect 6708 19101 6717 19135
rect 6717 19101 6751 19135
rect 6751 19101 6760 19135
rect 6708 19092 6760 19101
rect 2292 18999 2344 19008
rect 2292 18965 2301 18999
rect 2301 18965 2335 18999
rect 2335 18965 2344 18999
rect 2292 18956 2344 18965
rect 4446 18854 4498 18906
rect 4510 18854 4562 18906
rect 4574 18854 4626 18906
rect 4638 18854 4690 18906
rect 9774 18854 9826 18906
rect 9838 18854 9890 18906
rect 9902 18854 9954 18906
rect 9966 18854 10018 18906
rect 15102 18854 15154 18906
rect 15166 18854 15218 18906
rect 15230 18854 15282 18906
rect 15294 18854 15346 18906
rect 20430 18854 20482 18906
rect 20494 18854 20546 18906
rect 20558 18854 20610 18906
rect 20622 18854 20674 18906
rect 6708 18752 6760 18804
rect 2292 18548 2344 18600
rect 7110 18310 7162 18362
rect 7174 18310 7226 18362
rect 7238 18310 7290 18362
rect 7302 18310 7354 18362
rect 12438 18310 12490 18362
rect 12502 18310 12554 18362
rect 12566 18310 12618 18362
rect 12630 18310 12682 18362
rect 17766 18310 17818 18362
rect 17830 18310 17882 18362
rect 17894 18310 17946 18362
rect 17958 18310 18010 18362
rect 2292 18208 2344 18260
rect 2476 18115 2528 18124
rect 2476 18081 2485 18115
rect 2485 18081 2519 18115
rect 2519 18081 2528 18115
rect 2476 18072 2528 18081
rect 11492 18047 11544 18056
rect 11492 18013 11501 18047
rect 11501 18013 11535 18047
rect 11535 18013 11544 18047
rect 11492 18004 11544 18013
rect 2292 17911 2344 17920
rect 2292 17877 2301 17911
rect 2301 17877 2335 17911
rect 2335 17877 2344 17911
rect 2292 17868 2344 17877
rect 4446 17766 4498 17818
rect 4510 17766 4562 17818
rect 4574 17766 4626 17818
rect 4638 17766 4690 17818
rect 9774 17766 9826 17818
rect 9838 17766 9890 17818
rect 9902 17766 9954 17818
rect 9966 17766 10018 17818
rect 15102 17766 15154 17818
rect 15166 17766 15218 17818
rect 15230 17766 15282 17818
rect 15294 17766 15346 17818
rect 20430 17766 20482 17818
rect 20494 17766 20546 17818
rect 20558 17766 20610 17818
rect 20622 17766 20674 17818
rect 11492 17664 11544 17716
rect 2292 17528 2344 17580
rect 7110 17222 7162 17274
rect 7174 17222 7226 17274
rect 7238 17222 7290 17274
rect 7302 17222 7354 17274
rect 12438 17222 12490 17274
rect 12502 17222 12554 17274
rect 12566 17222 12618 17274
rect 12630 17222 12682 17274
rect 17766 17222 17818 17274
rect 17830 17222 17882 17274
rect 17894 17222 17946 17274
rect 17958 17222 18010 17274
rect 2292 17120 2344 17172
rect 2476 17027 2528 17036
rect 2476 16993 2485 17027
rect 2485 16993 2519 17027
rect 2519 16993 2528 17027
rect 2476 16984 2528 16993
rect 2292 16823 2344 16832
rect 2292 16789 2301 16823
rect 2301 16789 2335 16823
rect 2335 16789 2344 16823
rect 21612 16916 21664 16968
rect 2292 16780 2344 16789
rect 4446 16678 4498 16730
rect 4510 16678 4562 16730
rect 4574 16678 4626 16730
rect 4638 16678 4690 16730
rect 9774 16678 9826 16730
rect 9838 16678 9890 16730
rect 9902 16678 9954 16730
rect 9966 16678 10018 16730
rect 15102 16678 15154 16730
rect 15166 16678 15218 16730
rect 15230 16678 15282 16730
rect 15294 16678 15346 16730
rect 20430 16678 20482 16730
rect 20494 16678 20546 16730
rect 20558 16678 20610 16730
rect 20622 16678 20674 16730
rect 21612 16576 21664 16628
rect 2384 16372 2436 16424
rect 7110 16134 7162 16186
rect 7174 16134 7226 16186
rect 7238 16134 7290 16186
rect 7302 16134 7354 16186
rect 12438 16134 12490 16186
rect 12502 16134 12554 16186
rect 12566 16134 12618 16186
rect 12630 16134 12682 16186
rect 17766 16134 17818 16186
rect 17830 16134 17882 16186
rect 17894 16134 17946 16186
rect 17958 16134 18010 16186
rect 2384 15964 2436 16016
rect 2476 15939 2528 15948
rect 2476 15905 2485 15939
rect 2485 15905 2519 15939
rect 2519 15905 2528 15939
rect 2476 15896 2528 15905
rect 21060 15871 21112 15880
rect 2292 15735 2344 15744
rect 2292 15701 2301 15735
rect 2301 15701 2335 15735
rect 2335 15701 2344 15735
rect 21060 15837 21069 15871
rect 21069 15837 21103 15871
rect 21103 15837 21112 15871
rect 21060 15828 21112 15837
rect 2292 15692 2344 15701
rect 4446 15590 4498 15642
rect 4510 15590 4562 15642
rect 4574 15590 4626 15642
rect 4638 15590 4690 15642
rect 9774 15590 9826 15642
rect 9838 15590 9890 15642
rect 9902 15590 9954 15642
rect 9966 15590 10018 15642
rect 15102 15590 15154 15642
rect 15166 15590 15218 15642
rect 15230 15590 15282 15642
rect 15294 15590 15346 15642
rect 20430 15590 20482 15642
rect 20494 15590 20546 15642
rect 20558 15590 20610 15642
rect 20622 15590 20674 15642
rect 21060 15488 21112 15540
rect 3856 15352 3908 15404
rect 7110 15046 7162 15098
rect 7174 15046 7226 15098
rect 7238 15046 7290 15098
rect 7302 15046 7354 15098
rect 12438 15046 12490 15098
rect 12502 15046 12554 15098
rect 12566 15046 12618 15098
rect 12630 15046 12682 15098
rect 17766 15046 17818 15098
rect 17830 15046 17882 15098
rect 17894 15046 17946 15098
rect 17958 15046 18010 15098
rect 3856 14944 3908 14996
rect 21612 14740 21664 14792
rect 4446 14502 4498 14554
rect 4510 14502 4562 14554
rect 4574 14502 4626 14554
rect 4638 14502 4690 14554
rect 9774 14502 9826 14554
rect 9838 14502 9890 14554
rect 9902 14502 9954 14554
rect 9966 14502 10018 14554
rect 15102 14502 15154 14554
rect 15166 14502 15218 14554
rect 15230 14502 15282 14554
rect 15294 14502 15346 14554
rect 20430 14502 20482 14554
rect 20494 14502 20546 14554
rect 20558 14502 20610 14554
rect 20622 14502 20674 14554
rect 21612 14400 21664 14452
rect 2292 14264 2344 14316
rect 7110 13958 7162 14010
rect 7174 13958 7226 14010
rect 7238 13958 7290 14010
rect 7302 13958 7354 14010
rect 12438 13958 12490 14010
rect 12502 13958 12554 14010
rect 12566 13958 12618 14010
rect 12630 13958 12682 14010
rect 17766 13958 17818 14010
rect 17830 13958 17882 14010
rect 17894 13958 17946 14010
rect 17958 13958 18010 14010
rect 2292 13788 2344 13840
rect 2476 13763 2528 13772
rect 2476 13729 2485 13763
rect 2485 13729 2519 13763
rect 2519 13729 2528 13763
rect 2476 13720 2528 13729
rect 21060 13695 21112 13704
rect 2292 13559 2344 13568
rect 2292 13525 2301 13559
rect 2301 13525 2335 13559
rect 2335 13525 2344 13559
rect 21060 13661 21069 13695
rect 21069 13661 21103 13695
rect 21103 13661 21112 13695
rect 21060 13652 21112 13661
rect 2292 13516 2344 13525
rect 4446 13414 4498 13466
rect 4510 13414 4562 13466
rect 4574 13414 4626 13466
rect 4638 13414 4690 13466
rect 9774 13414 9826 13466
rect 9838 13414 9890 13466
rect 9902 13414 9954 13466
rect 9966 13414 10018 13466
rect 15102 13414 15154 13466
rect 15166 13414 15218 13466
rect 15230 13414 15282 13466
rect 15294 13414 15346 13466
rect 20430 13414 20482 13466
rect 20494 13414 20546 13466
rect 20558 13414 20610 13466
rect 20622 13414 20674 13466
rect 21060 13312 21112 13364
rect 3856 13176 3908 13228
rect 7110 12870 7162 12922
rect 7174 12870 7226 12922
rect 7238 12870 7290 12922
rect 7302 12870 7354 12922
rect 12438 12870 12490 12922
rect 12502 12870 12554 12922
rect 12566 12870 12618 12922
rect 12630 12870 12682 12922
rect 17766 12870 17818 12922
rect 17830 12870 17882 12922
rect 17894 12870 17946 12922
rect 17958 12870 18010 12922
rect 3856 12768 3908 12820
rect 21612 12564 21664 12616
rect 4446 12326 4498 12378
rect 4510 12326 4562 12378
rect 4574 12326 4626 12378
rect 4638 12326 4690 12378
rect 9774 12326 9826 12378
rect 9838 12326 9890 12378
rect 9902 12326 9954 12378
rect 9966 12326 10018 12378
rect 15102 12326 15154 12378
rect 15166 12326 15218 12378
rect 15230 12326 15282 12378
rect 15294 12326 15346 12378
rect 20430 12326 20482 12378
rect 20494 12326 20546 12378
rect 20558 12326 20610 12378
rect 20622 12326 20674 12378
rect 21612 12224 21664 12276
rect 3856 12088 3908 12140
rect 7110 11782 7162 11834
rect 7174 11782 7226 11834
rect 7238 11782 7290 11834
rect 7302 11782 7354 11834
rect 12438 11782 12490 11834
rect 12502 11782 12554 11834
rect 12566 11782 12618 11834
rect 12630 11782 12682 11834
rect 17766 11782 17818 11834
rect 17830 11782 17882 11834
rect 17894 11782 17946 11834
rect 17958 11782 18010 11834
rect 3856 11544 3908 11596
rect 21060 11519 21112 11528
rect 21060 11485 21069 11519
rect 21069 11485 21103 11519
rect 21103 11485 21112 11519
rect 21060 11476 21112 11485
rect 4446 11238 4498 11290
rect 4510 11238 4562 11290
rect 4574 11238 4626 11290
rect 4638 11238 4690 11290
rect 9774 11238 9826 11290
rect 9838 11238 9890 11290
rect 9902 11238 9954 11290
rect 9966 11238 10018 11290
rect 15102 11238 15154 11290
rect 15166 11238 15218 11290
rect 15230 11238 15282 11290
rect 15294 11238 15346 11290
rect 20430 11238 20482 11290
rect 20494 11238 20546 11290
rect 20558 11238 20610 11290
rect 20622 11238 20674 11290
rect 21060 11136 21112 11188
rect 3856 11000 3908 11052
rect 7110 10694 7162 10746
rect 7174 10694 7226 10746
rect 7238 10694 7290 10746
rect 7302 10694 7354 10746
rect 12438 10694 12490 10746
rect 12502 10694 12554 10746
rect 12566 10694 12618 10746
rect 12630 10694 12682 10746
rect 17766 10694 17818 10746
rect 17830 10694 17882 10746
rect 17894 10694 17946 10746
rect 17958 10694 18010 10746
rect 3856 10592 3908 10644
rect 21612 10388 21664 10440
rect 4446 10150 4498 10202
rect 4510 10150 4562 10202
rect 4574 10150 4626 10202
rect 4638 10150 4690 10202
rect 9774 10150 9826 10202
rect 9838 10150 9890 10202
rect 9902 10150 9954 10202
rect 9966 10150 10018 10202
rect 15102 10150 15154 10202
rect 15166 10150 15218 10202
rect 15230 10150 15282 10202
rect 15294 10150 15346 10202
rect 20430 10150 20482 10202
rect 20494 10150 20546 10202
rect 20558 10150 20610 10202
rect 20622 10150 20674 10202
rect 21612 10048 21664 10100
rect 2292 9912 2344 9964
rect 7110 9606 7162 9658
rect 7174 9606 7226 9658
rect 7238 9606 7290 9658
rect 7302 9606 7354 9658
rect 12438 9606 12490 9658
rect 12502 9606 12554 9658
rect 12566 9606 12618 9658
rect 12630 9606 12682 9658
rect 17766 9606 17818 9658
rect 17830 9606 17882 9658
rect 17894 9606 17946 9658
rect 17958 9606 18010 9658
rect 2476 9411 2528 9420
rect 2476 9377 2485 9411
rect 2485 9377 2519 9411
rect 2519 9377 2528 9411
rect 2476 9368 2528 9377
rect 2292 9300 2344 9352
rect 21060 9343 21112 9352
rect 2292 9207 2344 9216
rect 2292 9173 2301 9207
rect 2301 9173 2335 9207
rect 2335 9173 2344 9207
rect 21060 9309 21069 9343
rect 21069 9309 21103 9343
rect 21103 9309 21112 9343
rect 21060 9300 21112 9309
rect 2292 9164 2344 9173
rect 4446 9062 4498 9114
rect 4510 9062 4562 9114
rect 4574 9062 4626 9114
rect 4638 9062 4690 9114
rect 9774 9062 9826 9114
rect 9838 9062 9890 9114
rect 9902 9062 9954 9114
rect 9966 9062 10018 9114
rect 15102 9062 15154 9114
rect 15166 9062 15218 9114
rect 15230 9062 15282 9114
rect 15294 9062 15346 9114
rect 20430 9062 20482 9114
rect 20494 9062 20546 9114
rect 20558 9062 20610 9114
rect 20622 9062 20674 9114
rect 21060 8960 21112 9012
rect 3856 8824 3908 8876
rect 7110 8518 7162 8570
rect 7174 8518 7226 8570
rect 7238 8518 7290 8570
rect 7302 8518 7354 8570
rect 12438 8518 12490 8570
rect 12502 8518 12554 8570
rect 12566 8518 12618 8570
rect 12630 8518 12682 8570
rect 17766 8518 17818 8570
rect 17830 8518 17882 8570
rect 17894 8518 17946 8570
rect 17958 8518 18010 8570
rect 3856 8416 3908 8468
rect 21612 8212 21664 8264
rect 4446 7974 4498 8026
rect 4510 7974 4562 8026
rect 4574 7974 4626 8026
rect 4638 7974 4690 8026
rect 9774 7974 9826 8026
rect 9838 7974 9890 8026
rect 9902 7974 9954 8026
rect 9966 7974 10018 8026
rect 15102 7974 15154 8026
rect 15166 7974 15218 8026
rect 15230 7974 15282 8026
rect 15294 7974 15346 8026
rect 20430 7974 20482 8026
rect 20494 7974 20546 8026
rect 20558 7974 20610 8026
rect 20622 7974 20674 8026
rect 21612 7872 21664 7924
rect 3856 7736 3908 7788
rect 7110 7430 7162 7482
rect 7174 7430 7226 7482
rect 7238 7430 7290 7482
rect 7302 7430 7354 7482
rect 12438 7430 12490 7482
rect 12502 7430 12554 7482
rect 12566 7430 12618 7482
rect 12630 7430 12682 7482
rect 17766 7430 17818 7482
rect 17830 7430 17882 7482
rect 17894 7430 17946 7482
rect 17958 7430 18010 7482
rect 3856 7124 3908 7176
rect 21704 7124 21756 7176
rect 4446 6886 4498 6938
rect 4510 6886 4562 6938
rect 4574 6886 4626 6938
rect 4638 6886 4690 6938
rect 9774 6886 9826 6938
rect 9838 6886 9890 6938
rect 9902 6886 9954 6938
rect 9966 6886 10018 6938
rect 15102 6886 15154 6938
rect 15166 6886 15218 6938
rect 15230 6886 15282 6938
rect 15294 6886 15346 6938
rect 20430 6886 20482 6938
rect 20494 6886 20546 6938
rect 20558 6886 20610 6938
rect 20622 6886 20674 6938
rect 21704 6827 21756 6836
rect 21704 6793 21713 6827
rect 21713 6793 21747 6827
rect 21747 6793 21756 6827
rect 21704 6784 21756 6793
rect 3856 6648 3908 6700
rect 7110 6342 7162 6394
rect 7174 6342 7226 6394
rect 7238 6342 7290 6394
rect 7302 6342 7354 6394
rect 12438 6342 12490 6394
rect 12502 6342 12554 6394
rect 12566 6342 12618 6394
rect 12630 6342 12682 6394
rect 17766 6342 17818 6394
rect 17830 6342 17882 6394
rect 17894 6342 17946 6394
rect 17958 6342 18010 6394
rect 3856 6240 3908 6292
rect 21612 6036 21664 6088
rect 4446 5798 4498 5850
rect 4510 5798 4562 5850
rect 4574 5798 4626 5850
rect 4638 5798 4690 5850
rect 9774 5798 9826 5850
rect 9838 5798 9890 5850
rect 9902 5798 9954 5850
rect 9966 5798 10018 5850
rect 15102 5798 15154 5850
rect 15166 5798 15218 5850
rect 15230 5798 15282 5850
rect 15294 5798 15346 5850
rect 20430 5798 20482 5850
rect 20494 5798 20546 5850
rect 20558 5798 20610 5850
rect 20622 5798 20674 5850
rect 21612 5696 21664 5748
rect 3856 5560 3908 5612
rect 7110 5254 7162 5306
rect 7174 5254 7226 5306
rect 7238 5254 7290 5306
rect 7302 5254 7354 5306
rect 12438 5254 12490 5306
rect 12502 5254 12554 5306
rect 12566 5254 12618 5306
rect 12630 5254 12682 5306
rect 17766 5254 17818 5306
rect 17830 5254 17882 5306
rect 17894 5254 17946 5306
rect 17958 5254 18010 5306
rect 3856 4948 3908 5000
rect 17380 5016 17432 5068
rect 17564 4948 17616 5000
rect 21612 4948 21664 5000
rect 4446 4710 4498 4762
rect 4510 4710 4562 4762
rect 4574 4710 4626 4762
rect 4638 4710 4690 4762
rect 9774 4710 9826 4762
rect 9838 4710 9890 4762
rect 9902 4710 9954 4762
rect 9966 4710 10018 4762
rect 15102 4710 15154 4762
rect 15166 4710 15218 4762
rect 15230 4710 15282 4762
rect 15294 4710 15346 4762
rect 20430 4710 20482 4762
rect 20494 4710 20546 4762
rect 20558 4710 20610 4762
rect 20622 4710 20674 4762
rect 21612 4608 21664 4660
rect 3856 4472 3908 4524
rect 7110 4166 7162 4218
rect 7174 4166 7226 4218
rect 7238 4166 7290 4218
rect 7302 4166 7354 4218
rect 12438 4166 12490 4218
rect 12502 4166 12554 4218
rect 12566 4166 12618 4218
rect 12630 4166 12682 4218
rect 17766 4166 17818 4218
rect 17830 4166 17882 4218
rect 17894 4166 17946 4218
rect 17958 4166 18010 4218
rect 3856 4064 3908 4116
rect 21612 3860 21664 3912
rect 4446 3622 4498 3674
rect 4510 3622 4562 3674
rect 4574 3622 4626 3674
rect 4638 3622 4690 3674
rect 9774 3622 9826 3674
rect 9838 3622 9890 3674
rect 9902 3622 9954 3674
rect 9966 3622 10018 3674
rect 15102 3622 15154 3674
rect 15166 3622 15218 3674
rect 15230 3622 15282 3674
rect 15294 3622 15346 3674
rect 20430 3622 20482 3674
rect 20494 3622 20546 3674
rect 20558 3622 20610 3674
rect 20622 3622 20674 3674
rect 21612 3452 21664 3504
rect 3856 3384 3908 3436
rect 7110 3078 7162 3130
rect 7174 3078 7226 3130
rect 7238 3078 7290 3130
rect 7302 3078 7354 3130
rect 12438 3078 12490 3130
rect 12502 3078 12554 3130
rect 12566 3078 12618 3130
rect 12630 3078 12682 3130
rect 17766 3078 17818 3130
rect 17830 3078 17882 3130
rect 17894 3078 17946 3130
rect 17958 3078 18010 3130
rect 3856 2976 3908 3028
rect 17012 2840 17064 2892
rect 9652 2772 9704 2824
rect 17012 2704 17064 2756
rect 21612 2772 21664 2824
rect 9652 2636 9704 2688
rect 4446 2534 4498 2586
rect 4510 2534 4562 2586
rect 4574 2534 4626 2586
rect 4638 2534 4690 2586
rect 9774 2534 9826 2586
rect 9838 2534 9890 2586
rect 9902 2534 9954 2586
rect 9966 2534 10018 2586
rect 15102 2534 15154 2586
rect 15166 2534 15218 2586
rect 15230 2534 15282 2586
rect 15294 2534 15346 2586
rect 20430 2534 20482 2586
rect 20494 2534 20546 2586
rect 20558 2534 20610 2586
rect 20622 2534 20674 2586
rect 21612 2432 21664 2484
rect 3856 2296 3908 2348
rect 7110 1990 7162 2042
rect 7174 1990 7226 2042
rect 7238 1990 7290 2042
rect 7302 1990 7354 2042
rect 12438 1990 12490 2042
rect 12502 1990 12554 2042
rect 12566 1990 12618 2042
rect 12630 1990 12682 2042
rect 17766 1990 17818 2042
rect 17830 1990 17882 2042
rect 17894 1990 17946 2042
rect 17958 1990 18010 2042
rect 3856 1888 3908 1940
rect 21612 1684 21664 1736
rect 4446 1446 4498 1498
rect 4510 1446 4562 1498
rect 4574 1446 4626 1498
rect 4638 1446 4690 1498
rect 9774 1446 9826 1498
rect 9838 1446 9890 1498
rect 9902 1446 9954 1498
rect 9966 1446 10018 1498
rect 15102 1446 15154 1498
rect 15166 1446 15218 1498
rect 15230 1446 15282 1498
rect 15294 1446 15346 1498
rect 20430 1446 20482 1498
rect 20494 1446 20546 1498
rect 20558 1446 20610 1498
rect 20622 1446 20674 1498
rect 21612 1276 21664 1328
rect 2936 1140 2988 1192
rect 7110 902 7162 954
rect 7174 902 7226 954
rect 7238 902 7290 954
rect 7302 902 7354 954
rect 12438 902 12490 954
rect 12502 902 12554 954
rect 12566 902 12618 954
rect 12630 902 12682 954
rect 17766 902 17818 954
rect 17830 902 17882 954
rect 17894 902 17946 954
rect 17958 902 18010 954
<< metal2 >>
rect 1922 22376 1978 22385
rect 1922 22311 1978 22320
rect 1936 22074 1964 22311
rect 4420 22172 4716 22192
rect 4476 22170 4500 22172
rect 4556 22170 4580 22172
rect 4636 22170 4660 22172
rect 4498 22118 4500 22170
rect 4562 22118 4574 22170
rect 4636 22118 4638 22170
rect 4476 22116 4500 22118
rect 4556 22116 4580 22118
rect 4636 22116 4660 22118
rect 4420 22096 4716 22116
rect 9748 22172 10044 22192
rect 9804 22170 9828 22172
rect 9884 22170 9908 22172
rect 9964 22170 9988 22172
rect 9826 22118 9828 22170
rect 9890 22118 9902 22170
rect 9964 22118 9966 22170
rect 9804 22116 9828 22118
rect 9884 22116 9908 22118
rect 9964 22116 9988 22118
rect 9748 22096 10044 22116
rect 15076 22172 15372 22192
rect 15132 22170 15156 22172
rect 15212 22170 15236 22172
rect 15292 22170 15316 22172
rect 15154 22118 15156 22170
rect 15218 22118 15230 22170
rect 15292 22118 15294 22170
rect 15132 22116 15156 22118
rect 15212 22116 15236 22118
rect 15292 22116 15316 22118
rect 15076 22096 15372 22116
rect 20404 22172 20700 22192
rect 20460 22170 20484 22172
rect 20540 22170 20564 22172
rect 20620 22170 20644 22172
rect 20482 22118 20484 22170
rect 20546 22118 20558 22170
rect 20620 22118 20622 22170
rect 20460 22116 20484 22118
rect 20540 22116 20564 22118
rect 20620 22116 20644 22118
rect 20404 22096 20700 22116
rect 1924 22068 1976 22074
rect 1924 22010 1976 22016
rect 2292 22000 2344 22006
rect 2292 21942 2344 21948
rect 2304 21802 2332 21942
rect 2476 21864 2528 21870
rect 2474 21832 2476 21841
rect 2528 21832 2530 21841
rect 2292 21796 2344 21802
rect 2474 21767 2530 21776
rect 2292 21738 2344 21744
rect 2304 21530 2332 21738
rect 7084 21628 7380 21648
rect 7140 21626 7164 21628
rect 7220 21626 7244 21628
rect 7300 21626 7324 21628
rect 7162 21574 7164 21626
rect 7226 21574 7238 21626
rect 7300 21574 7302 21626
rect 7140 21572 7164 21574
rect 7220 21572 7244 21574
rect 7300 21572 7324 21574
rect 7084 21552 7380 21572
rect 12412 21628 12708 21648
rect 12468 21626 12492 21628
rect 12548 21626 12572 21628
rect 12628 21626 12652 21628
rect 12490 21574 12492 21626
rect 12554 21574 12566 21626
rect 12628 21574 12630 21626
rect 12468 21572 12492 21574
rect 12548 21572 12572 21574
rect 12628 21572 12652 21574
rect 12412 21552 12708 21572
rect 17740 21628 18036 21648
rect 17796 21626 17820 21628
rect 17876 21626 17900 21628
rect 17956 21626 17980 21628
rect 17818 21574 17820 21626
rect 17882 21574 17894 21626
rect 17956 21574 17958 21626
rect 17796 21572 17820 21574
rect 17876 21572 17900 21574
rect 17956 21572 17980 21574
rect 17740 21552 18036 21572
rect 2292 21524 2344 21530
rect 2292 21466 2344 21472
rect 2476 21388 2528 21394
rect 2476 21330 2528 21336
rect 3764 21388 3816 21394
rect 3764 21330 3816 21336
rect 2488 21297 2516 21330
rect 2474 21288 2530 21297
rect 2474 21223 2530 21232
rect 2292 21184 2344 21190
rect 2292 21126 2344 21132
rect 2304 20782 2332 21126
rect 3776 20986 3804 21330
rect 4420 21084 4716 21104
rect 4476 21082 4500 21084
rect 4556 21082 4580 21084
rect 4636 21082 4660 21084
rect 4498 21030 4500 21082
rect 4562 21030 4574 21082
rect 4636 21030 4638 21082
rect 4476 21028 4500 21030
rect 4556 21028 4580 21030
rect 4636 21028 4660 21030
rect 4420 21008 4716 21028
rect 9748 21084 10044 21104
rect 9804 21082 9828 21084
rect 9884 21082 9908 21084
rect 9964 21082 9988 21084
rect 9826 21030 9828 21082
rect 9890 21030 9902 21082
rect 9964 21030 9966 21082
rect 9804 21028 9828 21030
rect 9884 21028 9908 21030
rect 9964 21028 9988 21030
rect 9748 21008 10044 21028
rect 15076 21084 15372 21104
rect 15132 21082 15156 21084
rect 15212 21082 15236 21084
rect 15292 21082 15316 21084
rect 15154 21030 15156 21082
rect 15218 21030 15230 21082
rect 15292 21030 15294 21082
rect 15132 21028 15156 21030
rect 15212 21028 15236 21030
rect 15292 21028 15316 21030
rect 15076 21008 15372 21028
rect 20404 21084 20700 21104
rect 20460 21082 20484 21084
rect 20540 21082 20564 21084
rect 20620 21082 20644 21084
rect 20482 21030 20484 21082
rect 20546 21030 20558 21082
rect 20620 21030 20622 21082
rect 20460 21028 20484 21030
rect 20540 21028 20564 21030
rect 20620 21028 20644 21030
rect 20404 21008 20700 21028
rect 3764 20980 3816 20986
rect 3764 20922 3816 20928
rect 2292 20776 2344 20782
rect 2292 20718 2344 20724
rect 2304 20442 2332 20718
rect 7084 20540 7380 20560
rect 7140 20538 7164 20540
rect 7220 20538 7244 20540
rect 7300 20538 7324 20540
rect 7162 20486 7164 20538
rect 7226 20486 7238 20538
rect 7300 20486 7302 20538
rect 7140 20484 7164 20486
rect 7220 20484 7244 20486
rect 7300 20484 7324 20486
rect 7084 20464 7380 20484
rect 12412 20540 12708 20560
rect 12468 20538 12492 20540
rect 12548 20538 12572 20540
rect 12628 20538 12652 20540
rect 12490 20486 12492 20538
rect 12554 20486 12566 20538
rect 12628 20486 12630 20538
rect 12468 20484 12492 20486
rect 12548 20484 12572 20486
rect 12628 20484 12652 20486
rect 12412 20464 12708 20484
rect 17740 20540 18036 20560
rect 17796 20538 17820 20540
rect 17876 20538 17900 20540
rect 17956 20538 17980 20540
rect 17818 20486 17820 20538
rect 17882 20486 17894 20538
rect 17956 20486 17958 20538
rect 17796 20484 17820 20486
rect 17876 20484 17900 20486
rect 17956 20484 17980 20486
rect 17740 20464 18036 20484
rect 2292 20436 2344 20442
rect 2292 20378 2344 20384
rect 2476 20300 2528 20306
rect 2476 20242 2528 20248
rect 2488 20209 2516 20242
rect 4316 20232 4368 20238
rect 2474 20200 2530 20209
rect 4316 20174 4368 20180
rect 2474 20135 2530 20144
rect 2292 20096 2344 20102
rect 2292 20038 2344 20044
rect 2304 19694 2332 20038
rect 4328 19898 4356 20174
rect 4420 19996 4716 20016
rect 4476 19994 4500 19996
rect 4556 19994 4580 19996
rect 4636 19994 4660 19996
rect 4498 19942 4500 19994
rect 4562 19942 4574 19994
rect 4636 19942 4638 19994
rect 4476 19940 4500 19942
rect 4556 19940 4580 19942
rect 4636 19940 4660 19942
rect 4420 19920 4716 19940
rect 9748 19996 10044 20016
rect 9804 19994 9828 19996
rect 9884 19994 9908 19996
rect 9964 19994 9988 19996
rect 9826 19942 9828 19994
rect 9890 19942 9902 19994
rect 9964 19942 9966 19994
rect 9804 19940 9828 19942
rect 9884 19940 9908 19942
rect 9964 19940 9988 19942
rect 9748 19920 10044 19940
rect 15076 19996 15372 20016
rect 15132 19994 15156 19996
rect 15212 19994 15236 19996
rect 15292 19994 15316 19996
rect 15154 19942 15156 19994
rect 15218 19942 15230 19994
rect 15292 19942 15294 19994
rect 15132 19940 15156 19942
rect 15212 19940 15236 19942
rect 15292 19940 15316 19942
rect 15076 19920 15372 19940
rect 20404 19996 20700 20016
rect 20460 19994 20484 19996
rect 20540 19994 20564 19996
rect 20620 19994 20644 19996
rect 20482 19942 20484 19994
rect 20546 19942 20558 19994
rect 20620 19942 20622 19994
rect 20460 19940 20484 19942
rect 20540 19940 20564 19942
rect 20620 19940 20644 19942
rect 20404 19920 20700 19940
rect 4316 19892 4368 19898
rect 4316 19834 4368 19840
rect 2292 19688 2344 19694
rect 2292 19630 2344 19636
rect 2304 19354 2332 19630
rect 7084 19452 7380 19472
rect 7140 19450 7164 19452
rect 7220 19450 7244 19452
rect 7300 19450 7324 19452
rect 7162 19398 7164 19450
rect 7226 19398 7238 19450
rect 7300 19398 7302 19450
rect 7140 19396 7164 19398
rect 7220 19396 7244 19398
rect 7300 19396 7324 19398
rect 7084 19376 7380 19396
rect 12412 19452 12708 19472
rect 12468 19450 12492 19452
rect 12548 19450 12572 19452
rect 12628 19450 12652 19452
rect 12490 19398 12492 19450
rect 12554 19398 12566 19450
rect 12628 19398 12630 19450
rect 12468 19396 12492 19398
rect 12548 19396 12572 19398
rect 12628 19396 12652 19398
rect 12412 19376 12708 19396
rect 17740 19452 18036 19472
rect 17796 19450 17820 19452
rect 17876 19450 17900 19452
rect 17956 19450 17980 19452
rect 17818 19398 17820 19450
rect 17882 19398 17894 19450
rect 17956 19398 17958 19450
rect 17796 19396 17820 19398
rect 17876 19396 17900 19398
rect 17956 19396 17980 19398
rect 17740 19376 18036 19396
rect 2292 19348 2344 19354
rect 2292 19290 2344 19296
rect 2476 19212 2528 19218
rect 2476 19154 2528 19160
rect 2488 19121 2516 19154
rect 6708 19144 6760 19150
rect 2474 19112 2530 19121
rect 6708 19086 6760 19092
rect 2474 19047 2530 19056
rect 2292 19008 2344 19014
rect 2292 18950 2344 18956
rect 2304 18606 2332 18950
rect 4420 18908 4716 18928
rect 4476 18906 4500 18908
rect 4556 18906 4580 18908
rect 4636 18906 4660 18908
rect 4498 18854 4500 18906
rect 4562 18854 4574 18906
rect 4636 18854 4638 18906
rect 4476 18852 4500 18854
rect 4556 18852 4580 18854
rect 4636 18852 4660 18854
rect 4420 18832 4716 18852
rect 6720 18810 6748 19086
rect 9748 18908 10044 18928
rect 9804 18906 9828 18908
rect 9884 18906 9908 18908
rect 9964 18906 9988 18908
rect 9826 18854 9828 18906
rect 9890 18854 9902 18906
rect 9964 18854 9966 18906
rect 9804 18852 9828 18854
rect 9884 18852 9908 18854
rect 9964 18852 9988 18854
rect 9748 18832 10044 18852
rect 15076 18908 15372 18928
rect 15132 18906 15156 18908
rect 15212 18906 15236 18908
rect 15292 18906 15316 18908
rect 15154 18854 15156 18906
rect 15218 18854 15230 18906
rect 15292 18854 15294 18906
rect 15132 18852 15156 18854
rect 15212 18852 15236 18854
rect 15292 18852 15316 18854
rect 15076 18832 15372 18852
rect 20404 18908 20700 18928
rect 20460 18906 20484 18908
rect 20540 18906 20564 18908
rect 20620 18906 20644 18908
rect 20482 18854 20484 18906
rect 20546 18854 20558 18906
rect 20620 18854 20622 18906
rect 20460 18852 20484 18854
rect 20540 18852 20564 18854
rect 20620 18852 20644 18854
rect 20404 18832 20700 18852
rect 6708 18804 6760 18810
rect 6708 18746 6760 18752
rect 2292 18600 2344 18606
rect 2292 18542 2344 18548
rect 2304 18266 2332 18542
rect 7084 18364 7380 18384
rect 7140 18362 7164 18364
rect 7220 18362 7244 18364
rect 7300 18362 7324 18364
rect 7162 18310 7164 18362
rect 7226 18310 7238 18362
rect 7300 18310 7302 18362
rect 7140 18308 7164 18310
rect 7220 18308 7244 18310
rect 7300 18308 7324 18310
rect 7084 18288 7380 18308
rect 12412 18364 12708 18384
rect 12468 18362 12492 18364
rect 12548 18362 12572 18364
rect 12628 18362 12652 18364
rect 12490 18310 12492 18362
rect 12554 18310 12566 18362
rect 12628 18310 12630 18362
rect 12468 18308 12492 18310
rect 12548 18308 12572 18310
rect 12628 18308 12652 18310
rect 12412 18288 12708 18308
rect 17740 18364 18036 18384
rect 17796 18362 17820 18364
rect 17876 18362 17900 18364
rect 17956 18362 17980 18364
rect 17818 18310 17820 18362
rect 17882 18310 17894 18362
rect 17956 18310 17958 18362
rect 17796 18308 17820 18310
rect 17876 18308 17900 18310
rect 17956 18308 17980 18310
rect 17740 18288 18036 18308
rect 2292 18260 2344 18266
rect 2292 18202 2344 18208
rect 2476 18124 2528 18130
rect 2476 18066 2528 18072
rect 2488 18033 2516 18066
rect 11492 18056 11544 18062
rect 2474 18024 2530 18033
rect 11492 17998 11544 18004
rect 2474 17959 2530 17968
rect 2292 17920 2344 17926
rect 2292 17862 2344 17868
rect 2304 17586 2332 17862
rect 4420 17820 4716 17840
rect 4476 17818 4500 17820
rect 4556 17818 4580 17820
rect 4636 17818 4660 17820
rect 4498 17766 4500 17818
rect 4562 17766 4574 17818
rect 4636 17766 4638 17818
rect 4476 17764 4500 17766
rect 4556 17764 4580 17766
rect 4636 17764 4660 17766
rect 4420 17744 4716 17764
rect 9748 17820 10044 17840
rect 9804 17818 9828 17820
rect 9884 17818 9908 17820
rect 9964 17818 9988 17820
rect 9826 17766 9828 17818
rect 9890 17766 9902 17818
rect 9964 17766 9966 17818
rect 9804 17764 9828 17766
rect 9884 17764 9908 17766
rect 9964 17764 9988 17766
rect 9748 17744 10044 17764
rect 11504 17722 11532 17998
rect 15076 17820 15372 17840
rect 15132 17818 15156 17820
rect 15212 17818 15236 17820
rect 15292 17818 15316 17820
rect 15154 17766 15156 17818
rect 15218 17766 15230 17818
rect 15292 17766 15294 17818
rect 15132 17764 15156 17766
rect 15212 17764 15236 17766
rect 15292 17764 15316 17766
rect 15076 17744 15372 17764
rect 20404 17820 20700 17840
rect 20460 17818 20484 17820
rect 20540 17818 20564 17820
rect 20620 17818 20644 17820
rect 20482 17766 20484 17818
rect 20546 17766 20558 17818
rect 20620 17766 20622 17818
rect 20460 17764 20484 17766
rect 20540 17764 20564 17766
rect 20620 17764 20644 17766
rect 20404 17744 20700 17764
rect 11492 17716 11544 17722
rect 11492 17658 11544 17664
rect 2292 17580 2344 17586
rect 2292 17522 2344 17528
rect 2304 17178 2332 17522
rect 7084 17276 7380 17296
rect 7140 17274 7164 17276
rect 7220 17274 7244 17276
rect 7300 17274 7324 17276
rect 7162 17222 7164 17274
rect 7226 17222 7238 17274
rect 7300 17222 7302 17274
rect 7140 17220 7164 17222
rect 7220 17220 7244 17222
rect 7300 17220 7324 17222
rect 7084 17200 7380 17220
rect 12412 17276 12708 17296
rect 12468 17274 12492 17276
rect 12548 17274 12572 17276
rect 12628 17274 12652 17276
rect 12490 17222 12492 17274
rect 12554 17222 12566 17274
rect 12628 17222 12630 17274
rect 12468 17220 12492 17222
rect 12548 17220 12572 17222
rect 12628 17220 12652 17222
rect 12412 17200 12708 17220
rect 17740 17276 18036 17296
rect 17796 17274 17820 17276
rect 17876 17274 17900 17276
rect 17956 17274 17980 17276
rect 17818 17222 17820 17274
rect 17882 17222 17894 17274
rect 17956 17222 17958 17274
rect 17796 17220 17820 17222
rect 17876 17220 17900 17222
rect 17956 17220 17980 17222
rect 17740 17200 18036 17220
rect 2292 17172 2344 17178
rect 2292 17114 2344 17120
rect 2476 17036 2528 17042
rect 2476 16978 2528 16984
rect 2292 16832 2344 16838
rect 2292 16774 2344 16780
rect 2304 16514 2332 16774
rect 2304 16486 2424 16514
rect 2396 16430 2424 16486
rect 2384 16424 2436 16430
rect 2488 16401 2516 16978
rect 21612 16968 21664 16974
rect 21612 16910 21664 16916
rect 4420 16732 4716 16752
rect 4476 16730 4500 16732
rect 4556 16730 4580 16732
rect 4636 16730 4660 16732
rect 4498 16678 4500 16730
rect 4562 16678 4574 16730
rect 4636 16678 4638 16730
rect 4476 16676 4500 16678
rect 4556 16676 4580 16678
rect 4636 16676 4660 16678
rect 4420 16656 4716 16676
rect 9748 16732 10044 16752
rect 9804 16730 9828 16732
rect 9884 16730 9908 16732
rect 9964 16730 9988 16732
rect 9826 16678 9828 16730
rect 9890 16678 9902 16730
rect 9964 16678 9966 16730
rect 9804 16676 9828 16678
rect 9884 16676 9908 16678
rect 9964 16676 9988 16678
rect 9748 16656 10044 16676
rect 15076 16732 15372 16752
rect 15132 16730 15156 16732
rect 15212 16730 15236 16732
rect 15292 16730 15316 16732
rect 15154 16678 15156 16730
rect 15218 16678 15230 16730
rect 15292 16678 15294 16730
rect 15132 16676 15156 16678
rect 15212 16676 15236 16678
rect 15292 16676 15316 16678
rect 15076 16656 15372 16676
rect 20404 16732 20700 16752
rect 20460 16730 20484 16732
rect 20540 16730 20564 16732
rect 20620 16730 20644 16732
rect 20482 16678 20484 16730
rect 20546 16678 20558 16730
rect 20620 16678 20622 16730
rect 20460 16676 20484 16678
rect 20540 16676 20564 16678
rect 20620 16676 20644 16678
rect 20404 16656 20700 16676
rect 21624 16634 21652 16910
rect 21612 16628 21664 16634
rect 21612 16570 21664 16576
rect 2384 16366 2436 16372
rect 2474 16392 2530 16401
rect 2396 16022 2424 16366
rect 2474 16327 2530 16336
rect 7084 16188 7380 16208
rect 7140 16186 7164 16188
rect 7220 16186 7244 16188
rect 7300 16186 7324 16188
rect 7162 16134 7164 16186
rect 7226 16134 7238 16186
rect 7300 16134 7302 16186
rect 7140 16132 7164 16134
rect 7220 16132 7244 16134
rect 7300 16132 7324 16134
rect 7084 16112 7380 16132
rect 12412 16188 12708 16208
rect 12468 16186 12492 16188
rect 12548 16186 12572 16188
rect 12628 16186 12652 16188
rect 12490 16134 12492 16186
rect 12554 16134 12566 16186
rect 12628 16134 12630 16186
rect 12468 16132 12492 16134
rect 12548 16132 12572 16134
rect 12628 16132 12652 16134
rect 12412 16112 12708 16132
rect 17740 16188 18036 16208
rect 17796 16186 17820 16188
rect 17876 16186 17900 16188
rect 17956 16186 17980 16188
rect 17818 16134 17820 16186
rect 17882 16134 17894 16186
rect 17956 16134 17958 16186
rect 17796 16132 17820 16134
rect 17876 16132 17900 16134
rect 17956 16132 17980 16134
rect 17740 16112 18036 16132
rect 2384 16016 2436 16022
rect 2384 15958 2436 15964
rect 2476 15948 2528 15954
rect 2476 15890 2528 15896
rect 2488 15857 2516 15890
rect 21060 15880 21112 15886
rect 2474 15848 2530 15857
rect 21060 15822 21112 15828
rect 2474 15783 2530 15792
rect 2292 15744 2344 15750
rect 2292 15686 2344 15692
rect 2304 14322 2332 15686
rect 4420 15644 4716 15664
rect 4476 15642 4500 15644
rect 4556 15642 4580 15644
rect 4636 15642 4660 15644
rect 4498 15590 4500 15642
rect 4562 15590 4574 15642
rect 4636 15590 4638 15642
rect 4476 15588 4500 15590
rect 4556 15588 4580 15590
rect 4636 15588 4660 15590
rect 4420 15568 4716 15588
rect 9748 15644 10044 15664
rect 9804 15642 9828 15644
rect 9884 15642 9908 15644
rect 9964 15642 9988 15644
rect 9826 15590 9828 15642
rect 9890 15590 9902 15642
rect 9964 15590 9966 15642
rect 9804 15588 9828 15590
rect 9884 15588 9908 15590
rect 9964 15588 9988 15590
rect 9748 15568 10044 15588
rect 15076 15644 15372 15664
rect 15132 15642 15156 15644
rect 15212 15642 15236 15644
rect 15292 15642 15316 15644
rect 15154 15590 15156 15642
rect 15218 15590 15230 15642
rect 15292 15590 15294 15642
rect 15132 15588 15156 15590
rect 15212 15588 15236 15590
rect 15292 15588 15316 15590
rect 15076 15568 15372 15588
rect 20404 15644 20700 15664
rect 20460 15642 20484 15644
rect 20540 15642 20564 15644
rect 20620 15642 20644 15644
rect 20482 15590 20484 15642
rect 20546 15590 20558 15642
rect 20620 15590 20622 15642
rect 20460 15588 20484 15590
rect 20540 15588 20564 15590
rect 20620 15588 20644 15590
rect 20404 15568 20700 15588
rect 21072 15546 21100 15822
rect 21060 15540 21112 15546
rect 21060 15482 21112 15488
rect 3856 15404 3908 15410
rect 3856 15346 3908 15352
rect 3868 15002 3896 15346
rect 7084 15100 7380 15120
rect 7140 15098 7164 15100
rect 7220 15098 7244 15100
rect 7300 15098 7324 15100
rect 7162 15046 7164 15098
rect 7226 15046 7238 15098
rect 7300 15046 7302 15098
rect 7140 15044 7164 15046
rect 7220 15044 7244 15046
rect 7300 15044 7324 15046
rect 7084 15024 7380 15044
rect 12412 15100 12708 15120
rect 12468 15098 12492 15100
rect 12548 15098 12572 15100
rect 12628 15098 12652 15100
rect 12490 15046 12492 15098
rect 12554 15046 12566 15098
rect 12628 15046 12630 15098
rect 12468 15044 12492 15046
rect 12548 15044 12572 15046
rect 12628 15044 12652 15046
rect 12412 15024 12708 15044
rect 17740 15100 18036 15120
rect 17796 15098 17820 15100
rect 17876 15098 17900 15100
rect 17956 15098 17980 15100
rect 17818 15046 17820 15098
rect 17882 15046 17894 15098
rect 17956 15046 17958 15098
rect 17796 15044 17820 15046
rect 17876 15044 17900 15046
rect 17956 15044 17980 15046
rect 17740 15024 18036 15044
rect 3856 14996 3908 15002
rect 3856 14938 3908 14944
rect 21612 14792 21664 14798
rect 21612 14734 21664 14740
rect 4420 14556 4716 14576
rect 4476 14554 4500 14556
rect 4556 14554 4580 14556
rect 4636 14554 4660 14556
rect 4498 14502 4500 14554
rect 4562 14502 4574 14554
rect 4636 14502 4638 14554
rect 4476 14500 4500 14502
rect 4556 14500 4580 14502
rect 4636 14500 4660 14502
rect 4420 14480 4716 14500
rect 9748 14556 10044 14576
rect 9804 14554 9828 14556
rect 9884 14554 9908 14556
rect 9964 14554 9988 14556
rect 9826 14502 9828 14554
rect 9890 14502 9902 14554
rect 9964 14502 9966 14554
rect 9804 14500 9828 14502
rect 9884 14500 9908 14502
rect 9964 14500 9988 14502
rect 9748 14480 10044 14500
rect 15076 14556 15372 14576
rect 15132 14554 15156 14556
rect 15212 14554 15236 14556
rect 15292 14554 15316 14556
rect 15154 14502 15156 14554
rect 15218 14502 15230 14554
rect 15292 14502 15294 14554
rect 15132 14500 15156 14502
rect 15212 14500 15236 14502
rect 15292 14500 15316 14502
rect 15076 14480 15372 14500
rect 20404 14556 20700 14576
rect 20460 14554 20484 14556
rect 20540 14554 20564 14556
rect 20620 14554 20644 14556
rect 20482 14502 20484 14554
rect 20546 14502 20558 14554
rect 20620 14502 20622 14554
rect 20460 14500 20484 14502
rect 20540 14500 20564 14502
rect 20620 14500 20644 14502
rect 20404 14480 20700 14500
rect 21624 14458 21652 14734
rect 21612 14452 21664 14458
rect 21612 14394 21664 14400
rect 2292 14316 2344 14322
rect 2292 14258 2344 14264
rect 2304 13846 2332 14258
rect 7084 14012 7380 14032
rect 7140 14010 7164 14012
rect 7220 14010 7244 14012
rect 7300 14010 7324 14012
rect 7162 13958 7164 14010
rect 7226 13958 7238 14010
rect 7300 13958 7302 14010
rect 7140 13956 7164 13958
rect 7220 13956 7244 13958
rect 7300 13956 7324 13958
rect 7084 13936 7380 13956
rect 12412 14012 12708 14032
rect 12468 14010 12492 14012
rect 12548 14010 12572 14012
rect 12628 14010 12652 14012
rect 12490 13958 12492 14010
rect 12554 13958 12566 14010
rect 12628 13958 12630 14010
rect 12468 13956 12492 13958
rect 12548 13956 12572 13958
rect 12628 13956 12652 13958
rect 12412 13936 12708 13956
rect 17740 14012 18036 14032
rect 17796 14010 17820 14012
rect 17876 14010 17900 14012
rect 17956 14010 17980 14012
rect 17818 13958 17820 14010
rect 17882 13958 17894 14010
rect 17956 13958 17958 14010
rect 17796 13956 17820 13958
rect 17876 13956 17900 13958
rect 17956 13956 17980 13958
rect 17740 13936 18036 13956
rect 2292 13840 2344 13846
rect 2292 13782 2344 13788
rect 2476 13772 2528 13778
rect 2476 13714 2528 13720
rect 2488 13681 2516 13714
rect 21060 13704 21112 13710
rect 2474 13672 2530 13681
rect 21060 13646 21112 13652
rect 2474 13607 2530 13616
rect 2292 13568 2344 13574
rect 2292 13510 2344 13516
rect 2304 9970 2332 13510
rect 4420 13468 4716 13488
rect 4476 13466 4500 13468
rect 4556 13466 4580 13468
rect 4636 13466 4660 13468
rect 4498 13414 4500 13466
rect 4562 13414 4574 13466
rect 4636 13414 4638 13466
rect 4476 13412 4500 13414
rect 4556 13412 4580 13414
rect 4636 13412 4660 13414
rect 4420 13392 4716 13412
rect 9748 13468 10044 13488
rect 9804 13466 9828 13468
rect 9884 13466 9908 13468
rect 9964 13466 9988 13468
rect 9826 13414 9828 13466
rect 9890 13414 9902 13466
rect 9964 13414 9966 13466
rect 9804 13412 9828 13414
rect 9884 13412 9908 13414
rect 9964 13412 9988 13414
rect 9748 13392 10044 13412
rect 15076 13468 15372 13488
rect 15132 13466 15156 13468
rect 15212 13466 15236 13468
rect 15292 13466 15316 13468
rect 15154 13414 15156 13466
rect 15218 13414 15230 13466
rect 15292 13414 15294 13466
rect 15132 13412 15156 13414
rect 15212 13412 15236 13414
rect 15292 13412 15316 13414
rect 15076 13392 15372 13412
rect 20404 13468 20700 13488
rect 20460 13466 20484 13468
rect 20540 13466 20564 13468
rect 20620 13466 20644 13468
rect 20482 13414 20484 13466
rect 20546 13414 20558 13466
rect 20620 13414 20622 13466
rect 20460 13412 20484 13414
rect 20540 13412 20564 13414
rect 20620 13412 20644 13414
rect 20404 13392 20700 13412
rect 21072 13370 21100 13646
rect 21060 13364 21112 13370
rect 21060 13306 21112 13312
rect 3856 13228 3908 13234
rect 3856 13170 3908 13176
rect 3868 12826 3896 13170
rect 7084 12924 7380 12944
rect 7140 12922 7164 12924
rect 7220 12922 7244 12924
rect 7300 12922 7324 12924
rect 7162 12870 7164 12922
rect 7226 12870 7238 12922
rect 7300 12870 7302 12922
rect 7140 12868 7164 12870
rect 7220 12868 7244 12870
rect 7300 12868 7324 12870
rect 7084 12848 7380 12868
rect 12412 12924 12708 12944
rect 12468 12922 12492 12924
rect 12548 12922 12572 12924
rect 12628 12922 12652 12924
rect 12490 12870 12492 12922
rect 12554 12870 12566 12922
rect 12628 12870 12630 12922
rect 12468 12868 12492 12870
rect 12548 12868 12572 12870
rect 12628 12868 12652 12870
rect 12412 12848 12708 12868
rect 17740 12924 18036 12944
rect 17796 12922 17820 12924
rect 17876 12922 17900 12924
rect 17956 12922 17980 12924
rect 17818 12870 17820 12922
rect 17882 12870 17894 12922
rect 17956 12870 17958 12922
rect 17796 12868 17820 12870
rect 17876 12868 17900 12870
rect 17956 12868 17980 12870
rect 17740 12848 18036 12868
rect 3856 12820 3908 12826
rect 3856 12762 3908 12768
rect 21612 12616 21664 12622
rect 21612 12558 21664 12564
rect 4420 12380 4716 12400
rect 4476 12378 4500 12380
rect 4556 12378 4580 12380
rect 4636 12378 4660 12380
rect 4498 12326 4500 12378
rect 4562 12326 4574 12378
rect 4636 12326 4638 12378
rect 4476 12324 4500 12326
rect 4556 12324 4580 12326
rect 4636 12324 4660 12326
rect 4420 12304 4716 12324
rect 9748 12380 10044 12400
rect 9804 12378 9828 12380
rect 9884 12378 9908 12380
rect 9964 12378 9988 12380
rect 9826 12326 9828 12378
rect 9890 12326 9902 12378
rect 9964 12326 9966 12378
rect 9804 12324 9828 12326
rect 9884 12324 9908 12326
rect 9964 12324 9988 12326
rect 9748 12304 10044 12324
rect 15076 12380 15372 12400
rect 15132 12378 15156 12380
rect 15212 12378 15236 12380
rect 15292 12378 15316 12380
rect 15154 12326 15156 12378
rect 15218 12326 15230 12378
rect 15292 12326 15294 12378
rect 15132 12324 15156 12326
rect 15212 12324 15236 12326
rect 15292 12324 15316 12326
rect 15076 12304 15372 12324
rect 20404 12380 20700 12400
rect 20460 12378 20484 12380
rect 20540 12378 20564 12380
rect 20620 12378 20644 12380
rect 20482 12326 20484 12378
rect 20546 12326 20558 12378
rect 20620 12326 20622 12378
rect 20460 12324 20484 12326
rect 20540 12324 20564 12326
rect 20620 12324 20644 12326
rect 20404 12304 20700 12324
rect 21624 12282 21652 12558
rect 21612 12276 21664 12282
rect 21612 12218 21664 12224
rect 3856 12140 3908 12146
rect 3856 12082 3908 12088
rect 3868 11602 3896 12082
rect 7084 11836 7380 11856
rect 7140 11834 7164 11836
rect 7220 11834 7244 11836
rect 7300 11834 7324 11836
rect 7162 11782 7164 11834
rect 7226 11782 7238 11834
rect 7300 11782 7302 11834
rect 7140 11780 7164 11782
rect 7220 11780 7244 11782
rect 7300 11780 7324 11782
rect 7084 11760 7380 11780
rect 12412 11836 12708 11856
rect 12468 11834 12492 11836
rect 12548 11834 12572 11836
rect 12628 11834 12652 11836
rect 12490 11782 12492 11834
rect 12554 11782 12566 11834
rect 12628 11782 12630 11834
rect 12468 11780 12492 11782
rect 12548 11780 12572 11782
rect 12628 11780 12652 11782
rect 12412 11760 12708 11780
rect 17740 11836 18036 11856
rect 17796 11834 17820 11836
rect 17876 11834 17900 11836
rect 17956 11834 17980 11836
rect 17818 11782 17820 11834
rect 17882 11782 17894 11834
rect 17956 11782 17958 11834
rect 17796 11780 17820 11782
rect 17876 11780 17900 11782
rect 17956 11780 17980 11782
rect 17740 11760 18036 11780
rect 3856 11596 3908 11602
rect 3856 11538 3908 11544
rect 21060 11528 21112 11534
rect 21060 11470 21112 11476
rect 4420 11292 4716 11312
rect 4476 11290 4500 11292
rect 4556 11290 4580 11292
rect 4636 11290 4660 11292
rect 4498 11238 4500 11290
rect 4562 11238 4574 11290
rect 4636 11238 4638 11290
rect 4476 11236 4500 11238
rect 4556 11236 4580 11238
rect 4636 11236 4660 11238
rect 4420 11216 4716 11236
rect 9748 11292 10044 11312
rect 9804 11290 9828 11292
rect 9884 11290 9908 11292
rect 9964 11290 9988 11292
rect 9826 11238 9828 11290
rect 9890 11238 9902 11290
rect 9964 11238 9966 11290
rect 9804 11236 9828 11238
rect 9884 11236 9908 11238
rect 9964 11236 9988 11238
rect 9748 11216 10044 11236
rect 15076 11292 15372 11312
rect 15132 11290 15156 11292
rect 15212 11290 15236 11292
rect 15292 11290 15316 11292
rect 15154 11238 15156 11290
rect 15218 11238 15230 11290
rect 15292 11238 15294 11290
rect 15132 11236 15156 11238
rect 15212 11236 15236 11238
rect 15292 11236 15316 11238
rect 15076 11216 15372 11236
rect 20404 11292 20700 11312
rect 20460 11290 20484 11292
rect 20540 11290 20564 11292
rect 20620 11290 20644 11292
rect 20482 11238 20484 11290
rect 20546 11238 20558 11290
rect 20620 11238 20622 11290
rect 20460 11236 20484 11238
rect 20540 11236 20564 11238
rect 20620 11236 20644 11238
rect 20404 11216 20700 11236
rect 21072 11194 21100 11470
rect 21060 11188 21112 11194
rect 21060 11130 21112 11136
rect 3856 11052 3908 11058
rect 3856 10994 3908 11000
rect 3868 10650 3896 10994
rect 7084 10748 7380 10768
rect 7140 10746 7164 10748
rect 7220 10746 7244 10748
rect 7300 10746 7324 10748
rect 7162 10694 7164 10746
rect 7226 10694 7238 10746
rect 7300 10694 7302 10746
rect 7140 10692 7164 10694
rect 7220 10692 7244 10694
rect 7300 10692 7324 10694
rect 7084 10672 7380 10692
rect 12412 10748 12708 10768
rect 12468 10746 12492 10748
rect 12548 10746 12572 10748
rect 12628 10746 12652 10748
rect 12490 10694 12492 10746
rect 12554 10694 12566 10746
rect 12628 10694 12630 10746
rect 12468 10692 12492 10694
rect 12548 10692 12572 10694
rect 12628 10692 12652 10694
rect 12412 10672 12708 10692
rect 17740 10748 18036 10768
rect 17796 10746 17820 10748
rect 17876 10746 17900 10748
rect 17956 10746 17980 10748
rect 17818 10694 17820 10746
rect 17882 10694 17894 10746
rect 17956 10694 17958 10746
rect 17796 10692 17820 10694
rect 17876 10692 17900 10694
rect 17956 10692 17980 10694
rect 17740 10672 18036 10692
rect 3856 10644 3908 10650
rect 3856 10586 3908 10592
rect 21612 10440 21664 10446
rect 21612 10382 21664 10388
rect 4420 10204 4716 10224
rect 4476 10202 4500 10204
rect 4556 10202 4580 10204
rect 4636 10202 4660 10204
rect 4498 10150 4500 10202
rect 4562 10150 4574 10202
rect 4636 10150 4638 10202
rect 4476 10148 4500 10150
rect 4556 10148 4580 10150
rect 4636 10148 4660 10150
rect 4420 10128 4716 10148
rect 9748 10204 10044 10224
rect 9804 10202 9828 10204
rect 9884 10202 9908 10204
rect 9964 10202 9988 10204
rect 9826 10150 9828 10202
rect 9890 10150 9902 10202
rect 9964 10150 9966 10202
rect 9804 10148 9828 10150
rect 9884 10148 9908 10150
rect 9964 10148 9988 10150
rect 9748 10128 10044 10148
rect 15076 10204 15372 10224
rect 15132 10202 15156 10204
rect 15212 10202 15236 10204
rect 15292 10202 15316 10204
rect 15154 10150 15156 10202
rect 15218 10150 15230 10202
rect 15292 10150 15294 10202
rect 15132 10148 15156 10150
rect 15212 10148 15236 10150
rect 15292 10148 15316 10150
rect 15076 10128 15372 10148
rect 20404 10204 20700 10224
rect 20460 10202 20484 10204
rect 20540 10202 20564 10204
rect 20620 10202 20644 10204
rect 20482 10150 20484 10202
rect 20546 10150 20558 10202
rect 20620 10150 20622 10202
rect 20460 10148 20484 10150
rect 20540 10148 20564 10150
rect 20620 10148 20644 10150
rect 20404 10128 20700 10148
rect 21624 10106 21652 10382
rect 21612 10100 21664 10106
rect 21612 10042 21664 10048
rect 2292 9964 2344 9970
rect 2292 9906 2344 9912
rect 2304 9358 2332 9906
rect 7084 9660 7380 9680
rect 7140 9658 7164 9660
rect 7220 9658 7244 9660
rect 7300 9658 7324 9660
rect 7162 9606 7164 9658
rect 7226 9606 7238 9658
rect 7300 9606 7302 9658
rect 7140 9604 7164 9606
rect 7220 9604 7244 9606
rect 7300 9604 7324 9606
rect 7084 9584 7380 9604
rect 12412 9660 12708 9680
rect 12468 9658 12492 9660
rect 12548 9658 12572 9660
rect 12628 9658 12652 9660
rect 12490 9606 12492 9658
rect 12554 9606 12566 9658
rect 12628 9606 12630 9658
rect 12468 9604 12492 9606
rect 12548 9604 12572 9606
rect 12628 9604 12652 9606
rect 12412 9584 12708 9604
rect 17740 9660 18036 9680
rect 17796 9658 17820 9660
rect 17876 9658 17900 9660
rect 17956 9658 17980 9660
rect 17818 9606 17820 9658
rect 17882 9606 17894 9658
rect 17956 9606 17958 9658
rect 17796 9604 17820 9606
rect 17876 9604 17900 9606
rect 17956 9604 17980 9606
rect 17740 9584 18036 9604
rect 2476 9420 2528 9426
rect 2476 9362 2528 9368
rect 2292 9352 2344 9358
rect 2292 9294 2344 9300
rect 2292 9216 2344 9222
rect 2292 9158 2344 9164
rect 2304 1169 2332 9158
rect 2488 8785 2516 9362
rect 21060 9352 21112 9358
rect 21060 9294 21112 9300
rect 4420 9116 4716 9136
rect 4476 9114 4500 9116
rect 4556 9114 4580 9116
rect 4636 9114 4660 9116
rect 4498 9062 4500 9114
rect 4562 9062 4574 9114
rect 4636 9062 4638 9114
rect 4476 9060 4500 9062
rect 4556 9060 4580 9062
rect 4636 9060 4660 9062
rect 4420 9040 4716 9060
rect 9748 9116 10044 9136
rect 9804 9114 9828 9116
rect 9884 9114 9908 9116
rect 9964 9114 9988 9116
rect 9826 9062 9828 9114
rect 9890 9062 9902 9114
rect 9964 9062 9966 9114
rect 9804 9060 9828 9062
rect 9884 9060 9908 9062
rect 9964 9060 9988 9062
rect 9748 9040 10044 9060
rect 15076 9116 15372 9136
rect 15132 9114 15156 9116
rect 15212 9114 15236 9116
rect 15292 9114 15316 9116
rect 15154 9062 15156 9114
rect 15218 9062 15230 9114
rect 15292 9062 15294 9114
rect 15132 9060 15156 9062
rect 15212 9060 15236 9062
rect 15292 9060 15316 9062
rect 15076 9040 15372 9060
rect 20404 9116 20700 9136
rect 20460 9114 20484 9116
rect 20540 9114 20564 9116
rect 20620 9114 20644 9116
rect 20482 9062 20484 9114
rect 20546 9062 20558 9114
rect 20620 9062 20622 9114
rect 20460 9060 20484 9062
rect 20540 9060 20564 9062
rect 20620 9060 20644 9062
rect 20404 9040 20700 9060
rect 21072 9018 21100 9294
rect 21060 9012 21112 9018
rect 21060 8954 21112 8960
rect 3856 8876 3908 8882
rect 3856 8818 3908 8824
rect 2474 8776 2530 8785
rect 2474 8711 2530 8720
rect 3868 8474 3896 8818
rect 7084 8572 7380 8592
rect 7140 8570 7164 8572
rect 7220 8570 7244 8572
rect 7300 8570 7324 8572
rect 7162 8518 7164 8570
rect 7226 8518 7238 8570
rect 7300 8518 7302 8570
rect 7140 8516 7164 8518
rect 7220 8516 7244 8518
rect 7300 8516 7324 8518
rect 7084 8496 7380 8516
rect 12412 8572 12708 8592
rect 12468 8570 12492 8572
rect 12548 8570 12572 8572
rect 12628 8570 12652 8572
rect 12490 8518 12492 8570
rect 12554 8518 12566 8570
rect 12628 8518 12630 8570
rect 12468 8516 12492 8518
rect 12548 8516 12572 8518
rect 12628 8516 12652 8518
rect 12412 8496 12708 8516
rect 17740 8572 18036 8592
rect 17796 8570 17820 8572
rect 17876 8570 17900 8572
rect 17956 8570 17980 8572
rect 17818 8518 17820 8570
rect 17882 8518 17894 8570
rect 17956 8518 17958 8570
rect 17796 8516 17820 8518
rect 17876 8516 17900 8518
rect 17956 8516 17980 8518
rect 17740 8496 18036 8516
rect 3856 8468 3908 8474
rect 3856 8410 3908 8416
rect 21612 8264 21664 8270
rect 21612 8206 21664 8212
rect 4420 8028 4716 8048
rect 4476 8026 4500 8028
rect 4556 8026 4580 8028
rect 4636 8026 4660 8028
rect 4498 7974 4500 8026
rect 4562 7974 4574 8026
rect 4636 7974 4638 8026
rect 4476 7972 4500 7974
rect 4556 7972 4580 7974
rect 4636 7972 4660 7974
rect 4420 7952 4716 7972
rect 9748 8028 10044 8048
rect 9804 8026 9828 8028
rect 9884 8026 9908 8028
rect 9964 8026 9988 8028
rect 9826 7974 9828 8026
rect 9890 7974 9902 8026
rect 9964 7974 9966 8026
rect 9804 7972 9828 7974
rect 9884 7972 9908 7974
rect 9964 7972 9988 7974
rect 9748 7952 10044 7972
rect 15076 8028 15372 8048
rect 15132 8026 15156 8028
rect 15212 8026 15236 8028
rect 15292 8026 15316 8028
rect 15154 7974 15156 8026
rect 15218 7974 15230 8026
rect 15292 7974 15294 8026
rect 15132 7972 15156 7974
rect 15212 7972 15236 7974
rect 15292 7972 15316 7974
rect 15076 7952 15372 7972
rect 20404 8028 20700 8048
rect 20460 8026 20484 8028
rect 20540 8026 20564 8028
rect 20620 8026 20644 8028
rect 20482 7974 20484 8026
rect 20546 7974 20558 8026
rect 20620 7974 20622 8026
rect 20460 7972 20484 7974
rect 20540 7972 20564 7974
rect 20620 7972 20644 7974
rect 20404 7952 20700 7972
rect 21624 7930 21652 8206
rect 21612 7924 21664 7930
rect 21612 7866 21664 7872
rect 3856 7788 3908 7794
rect 3856 7730 3908 7736
rect 3868 7182 3896 7730
rect 7084 7484 7380 7504
rect 7140 7482 7164 7484
rect 7220 7482 7244 7484
rect 7300 7482 7324 7484
rect 7162 7430 7164 7482
rect 7226 7430 7238 7482
rect 7300 7430 7302 7482
rect 7140 7428 7164 7430
rect 7220 7428 7244 7430
rect 7300 7428 7324 7430
rect 7084 7408 7380 7428
rect 12412 7484 12708 7504
rect 12468 7482 12492 7484
rect 12548 7482 12572 7484
rect 12628 7482 12652 7484
rect 12490 7430 12492 7482
rect 12554 7430 12566 7482
rect 12628 7430 12630 7482
rect 12468 7428 12492 7430
rect 12548 7428 12572 7430
rect 12628 7428 12652 7430
rect 12412 7408 12708 7428
rect 17740 7484 18036 7504
rect 17796 7482 17820 7484
rect 17876 7482 17900 7484
rect 17956 7482 17980 7484
rect 17818 7430 17820 7482
rect 17882 7430 17894 7482
rect 17956 7430 17958 7482
rect 17796 7428 17820 7430
rect 17876 7428 17900 7430
rect 17956 7428 17980 7430
rect 17740 7408 18036 7428
rect 3856 7176 3908 7182
rect 3856 7118 3908 7124
rect 21704 7176 21756 7182
rect 21704 7118 21756 7124
rect 4420 6940 4716 6960
rect 4476 6938 4500 6940
rect 4556 6938 4580 6940
rect 4636 6938 4660 6940
rect 4498 6886 4500 6938
rect 4562 6886 4574 6938
rect 4636 6886 4638 6938
rect 4476 6884 4500 6886
rect 4556 6884 4580 6886
rect 4636 6884 4660 6886
rect 4420 6864 4716 6884
rect 9748 6940 10044 6960
rect 9804 6938 9828 6940
rect 9884 6938 9908 6940
rect 9964 6938 9988 6940
rect 9826 6886 9828 6938
rect 9890 6886 9902 6938
rect 9964 6886 9966 6938
rect 9804 6884 9828 6886
rect 9884 6884 9908 6886
rect 9964 6884 9988 6886
rect 9748 6864 10044 6884
rect 15076 6940 15372 6960
rect 15132 6938 15156 6940
rect 15212 6938 15236 6940
rect 15292 6938 15316 6940
rect 15154 6886 15156 6938
rect 15218 6886 15230 6938
rect 15292 6886 15294 6938
rect 15132 6884 15156 6886
rect 15212 6884 15236 6886
rect 15292 6884 15316 6886
rect 15076 6864 15372 6884
rect 20404 6940 20700 6960
rect 20460 6938 20484 6940
rect 20540 6938 20564 6940
rect 20620 6938 20644 6940
rect 20482 6886 20484 6938
rect 20546 6886 20558 6938
rect 20620 6886 20622 6938
rect 20460 6884 20484 6886
rect 20540 6884 20564 6886
rect 20620 6884 20644 6886
rect 20404 6864 20700 6884
rect 21716 6842 21744 7118
rect 21704 6836 21756 6842
rect 21704 6778 21756 6784
rect 3856 6700 3908 6706
rect 3856 6642 3908 6648
rect 3868 6298 3896 6642
rect 7084 6396 7380 6416
rect 7140 6394 7164 6396
rect 7220 6394 7244 6396
rect 7300 6394 7324 6396
rect 7162 6342 7164 6394
rect 7226 6342 7238 6394
rect 7300 6342 7302 6394
rect 7140 6340 7164 6342
rect 7220 6340 7244 6342
rect 7300 6340 7324 6342
rect 7084 6320 7380 6340
rect 12412 6396 12708 6416
rect 12468 6394 12492 6396
rect 12548 6394 12572 6396
rect 12628 6394 12652 6396
rect 12490 6342 12492 6394
rect 12554 6342 12566 6394
rect 12628 6342 12630 6394
rect 12468 6340 12492 6342
rect 12548 6340 12572 6342
rect 12628 6340 12652 6342
rect 12412 6320 12708 6340
rect 17740 6396 18036 6416
rect 17796 6394 17820 6396
rect 17876 6394 17900 6396
rect 17956 6394 17980 6396
rect 17818 6342 17820 6394
rect 17882 6342 17894 6394
rect 17956 6342 17958 6394
rect 17796 6340 17820 6342
rect 17876 6340 17900 6342
rect 17956 6340 17980 6342
rect 17740 6320 18036 6340
rect 3856 6292 3908 6298
rect 3856 6234 3908 6240
rect 21612 6088 21664 6094
rect 21612 6030 21664 6036
rect 4420 5852 4716 5872
rect 4476 5850 4500 5852
rect 4556 5850 4580 5852
rect 4636 5850 4660 5852
rect 4498 5798 4500 5850
rect 4562 5798 4574 5850
rect 4636 5798 4638 5850
rect 4476 5796 4500 5798
rect 4556 5796 4580 5798
rect 4636 5796 4660 5798
rect 4420 5776 4716 5796
rect 9748 5852 10044 5872
rect 9804 5850 9828 5852
rect 9884 5850 9908 5852
rect 9964 5850 9988 5852
rect 9826 5798 9828 5850
rect 9890 5798 9902 5850
rect 9964 5798 9966 5850
rect 9804 5796 9828 5798
rect 9884 5796 9908 5798
rect 9964 5796 9988 5798
rect 9748 5776 10044 5796
rect 15076 5852 15372 5872
rect 15132 5850 15156 5852
rect 15212 5850 15236 5852
rect 15292 5850 15316 5852
rect 15154 5798 15156 5850
rect 15218 5798 15230 5850
rect 15292 5798 15294 5850
rect 15132 5796 15156 5798
rect 15212 5796 15236 5798
rect 15292 5796 15316 5798
rect 15076 5776 15372 5796
rect 20404 5852 20700 5872
rect 20460 5850 20484 5852
rect 20540 5850 20564 5852
rect 20620 5850 20644 5852
rect 20482 5798 20484 5850
rect 20546 5798 20558 5850
rect 20620 5798 20622 5850
rect 20460 5796 20484 5798
rect 20540 5796 20564 5798
rect 20620 5796 20644 5798
rect 20404 5776 20700 5796
rect 21624 5754 21652 6030
rect 21612 5748 21664 5754
rect 21612 5690 21664 5696
rect 3856 5612 3908 5618
rect 3856 5554 3908 5560
rect 3868 5006 3896 5554
rect 7084 5308 7380 5328
rect 7140 5306 7164 5308
rect 7220 5306 7244 5308
rect 7300 5306 7324 5308
rect 7162 5254 7164 5306
rect 7226 5254 7238 5306
rect 7300 5254 7302 5306
rect 7140 5252 7164 5254
rect 7220 5252 7244 5254
rect 7300 5252 7324 5254
rect 7084 5232 7380 5252
rect 12412 5308 12708 5328
rect 12468 5306 12492 5308
rect 12548 5306 12572 5308
rect 12628 5306 12652 5308
rect 12490 5254 12492 5306
rect 12554 5254 12566 5306
rect 12628 5254 12630 5306
rect 12468 5252 12492 5254
rect 12548 5252 12572 5254
rect 12628 5252 12652 5254
rect 12412 5232 12708 5252
rect 17740 5308 18036 5328
rect 17796 5306 17820 5308
rect 17876 5306 17900 5308
rect 17956 5306 17980 5308
rect 17818 5254 17820 5306
rect 17882 5254 17894 5306
rect 17956 5254 17958 5306
rect 17796 5252 17820 5254
rect 17876 5252 17900 5254
rect 17956 5252 17980 5254
rect 17740 5232 18036 5252
rect 17380 5068 17432 5074
rect 17380 5010 17432 5016
rect 3856 5000 3908 5006
rect 3856 4942 3908 4948
rect 17392 4954 17420 5010
rect 17564 5000 17616 5006
rect 17392 4948 17564 4954
rect 17392 4942 17616 4948
rect 21612 5000 21664 5006
rect 21612 4942 21664 4948
rect 17392 4926 17604 4942
rect 4420 4764 4716 4784
rect 4476 4762 4500 4764
rect 4556 4762 4580 4764
rect 4636 4762 4660 4764
rect 4498 4710 4500 4762
rect 4562 4710 4574 4762
rect 4636 4710 4638 4762
rect 4476 4708 4500 4710
rect 4556 4708 4580 4710
rect 4636 4708 4660 4710
rect 4420 4688 4716 4708
rect 9748 4764 10044 4784
rect 9804 4762 9828 4764
rect 9884 4762 9908 4764
rect 9964 4762 9988 4764
rect 9826 4710 9828 4762
rect 9890 4710 9902 4762
rect 9964 4710 9966 4762
rect 9804 4708 9828 4710
rect 9884 4708 9908 4710
rect 9964 4708 9988 4710
rect 9748 4688 10044 4708
rect 15076 4764 15372 4784
rect 15132 4762 15156 4764
rect 15212 4762 15236 4764
rect 15292 4762 15316 4764
rect 15154 4710 15156 4762
rect 15218 4710 15230 4762
rect 15292 4710 15294 4762
rect 15132 4708 15156 4710
rect 15212 4708 15236 4710
rect 15292 4708 15316 4710
rect 15076 4688 15372 4708
rect 20404 4764 20700 4784
rect 20460 4762 20484 4764
rect 20540 4762 20564 4764
rect 20620 4762 20644 4764
rect 20482 4710 20484 4762
rect 20546 4710 20558 4762
rect 20620 4710 20622 4762
rect 20460 4708 20484 4710
rect 20540 4708 20564 4710
rect 20620 4708 20644 4710
rect 20404 4688 20700 4708
rect 21624 4666 21652 4942
rect 21612 4660 21664 4666
rect 21612 4602 21664 4608
rect 3856 4524 3908 4530
rect 3856 4466 3908 4472
rect 3868 4122 3896 4466
rect 7084 4220 7380 4240
rect 7140 4218 7164 4220
rect 7220 4218 7244 4220
rect 7300 4218 7324 4220
rect 7162 4166 7164 4218
rect 7226 4166 7238 4218
rect 7300 4166 7302 4218
rect 7140 4164 7164 4166
rect 7220 4164 7244 4166
rect 7300 4164 7324 4166
rect 7084 4144 7380 4164
rect 12412 4220 12708 4240
rect 12468 4218 12492 4220
rect 12548 4218 12572 4220
rect 12628 4218 12652 4220
rect 12490 4166 12492 4218
rect 12554 4166 12566 4218
rect 12628 4166 12630 4218
rect 12468 4164 12492 4166
rect 12548 4164 12572 4166
rect 12628 4164 12652 4166
rect 12412 4144 12708 4164
rect 17740 4220 18036 4240
rect 17796 4218 17820 4220
rect 17876 4218 17900 4220
rect 17956 4218 17980 4220
rect 17818 4166 17820 4218
rect 17882 4166 17894 4218
rect 17956 4166 17958 4218
rect 17796 4164 17820 4166
rect 17876 4164 17900 4166
rect 17956 4164 17980 4166
rect 17740 4144 18036 4164
rect 3856 4116 3908 4122
rect 3856 4058 3908 4064
rect 21612 3912 21664 3918
rect 21612 3854 21664 3860
rect 4420 3676 4716 3696
rect 4476 3674 4500 3676
rect 4556 3674 4580 3676
rect 4636 3674 4660 3676
rect 4498 3622 4500 3674
rect 4562 3622 4574 3674
rect 4636 3622 4638 3674
rect 4476 3620 4500 3622
rect 4556 3620 4580 3622
rect 4636 3620 4660 3622
rect 4420 3600 4716 3620
rect 9748 3676 10044 3696
rect 9804 3674 9828 3676
rect 9884 3674 9908 3676
rect 9964 3674 9988 3676
rect 9826 3622 9828 3674
rect 9890 3622 9902 3674
rect 9964 3622 9966 3674
rect 9804 3620 9828 3622
rect 9884 3620 9908 3622
rect 9964 3620 9988 3622
rect 9748 3600 10044 3620
rect 15076 3676 15372 3696
rect 15132 3674 15156 3676
rect 15212 3674 15236 3676
rect 15292 3674 15316 3676
rect 15154 3622 15156 3674
rect 15218 3622 15230 3674
rect 15292 3622 15294 3674
rect 15132 3620 15156 3622
rect 15212 3620 15236 3622
rect 15292 3620 15316 3622
rect 15076 3600 15372 3620
rect 20404 3676 20700 3696
rect 20460 3674 20484 3676
rect 20540 3674 20564 3676
rect 20620 3674 20644 3676
rect 20482 3622 20484 3674
rect 20546 3622 20558 3674
rect 20620 3622 20622 3674
rect 20460 3620 20484 3622
rect 20540 3620 20564 3622
rect 20620 3620 20644 3622
rect 20404 3600 20700 3620
rect 21624 3510 21652 3854
rect 21612 3504 21664 3510
rect 21612 3446 21664 3452
rect 3856 3436 3908 3442
rect 3856 3378 3908 3384
rect 3868 3034 3896 3378
rect 7084 3132 7380 3152
rect 7140 3130 7164 3132
rect 7220 3130 7244 3132
rect 7300 3130 7324 3132
rect 7162 3078 7164 3130
rect 7226 3078 7238 3130
rect 7300 3078 7302 3130
rect 7140 3076 7164 3078
rect 7220 3076 7244 3078
rect 7300 3076 7324 3078
rect 7084 3056 7380 3076
rect 12412 3132 12708 3152
rect 12468 3130 12492 3132
rect 12548 3130 12572 3132
rect 12628 3130 12652 3132
rect 12490 3078 12492 3130
rect 12554 3078 12566 3130
rect 12628 3078 12630 3130
rect 12468 3076 12492 3078
rect 12548 3076 12572 3078
rect 12628 3076 12652 3078
rect 12412 3056 12708 3076
rect 17740 3132 18036 3152
rect 17796 3130 17820 3132
rect 17876 3130 17900 3132
rect 17956 3130 17980 3132
rect 17818 3078 17820 3130
rect 17882 3078 17894 3130
rect 17956 3078 17958 3130
rect 17796 3076 17820 3078
rect 17876 3076 17900 3078
rect 17956 3076 17980 3078
rect 17740 3056 18036 3076
rect 3856 3028 3908 3034
rect 3856 2970 3908 2976
rect 17012 2892 17064 2898
rect 17012 2834 17064 2840
rect 9652 2824 9704 2830
rect 9652 2766 9704 2772
rect 9664 2694 9692 2766
rect 17024 2762 17052 2834
rect 21612 2824 21664 2830
rect 21612 2766 21664 2772
rect 17012 2756 17064 2762
rect 17012 2698 17064 2704
rect 9652 2688 9704 2694
rect 9652 2630 9704 2636
rect 4420 2588 4716 2608
rect 4476 2586 4500 2588
rect 4556 2586 4580 2588
rect 4636 2586 4660 2588
rect 4498 2534 4500 2586
rect 4562 2534 4574 2586
rect 4636 2534 4638 2586
rect 4476 2532 4500 2534
rect 4556 2532 4580 2534
rect 4636 2532 4660 2534
rect 4420 2512 4716 2532
rect 9748 2588 10044 2608
rect 9804 2586 9828 2588
rect 9884 2586 9908 2588
rect 9964 2586 9988 2588
rect 9826 2534 9828 2586
rect 9890 2534 9902 2586
rect 9964 2534 9966 2586
rect 9804 2532 9828 2534
rect 9884 2532 9908 2534
rect 9964 2532 9988 2534
rect 9748 2512 10044 2532
rect 15076 2588 15372 2608
rect 15132 2586 15156 2588
rect 15212 2586 15236 2588
rect 15292 2586 15316 2588
rect 15154 2534 15156 2586
rect 15218 2534 15230 2586
rect 15292 2534 15294 2586
rect 15132 2532 15156 2534
rect 15212 2532 15236 2534
rect 15292 2532 15316 2534
rect 15076 2512 15372 2532
rect 20404 2588 20700 2608
rect 20460 2586 20484 2588
rect 20540 2586 20564 2588
rect 20620 2586 20644 2588
rect 20482 2534 20484 2586
rect 20546 2534 20558 2586
rect 20620 2534 20622 2586
rect 20460 2532 20484 2534
rect 20540 2532 20564 2534
rect 20620 2532 20644 2534
rect 20404 2512 20700 2532
rect 21624 2490 21652 2766
rect 21612 2484 21664 2490
rect 21612 2426 21664 2432
rect 3856 2348 3908 2354
rect 3856 2290 3908 2296
rect 3868 1946 3896 2290
rect 7084 2044 7380 2064
rect 7140 2042 7164 2044
rect 7220 2042 7244 2044
rect 7300 2042 7324 2044
rect 7162 1990 7164 2042
rect 7226 1990 7238 2042
rect 7300 1990 7302 2042
rect 7140 1988 7164 1990
rect 7220 1988 7244 1990
rect 7300 1988 7324 1990
rect 7084 1968 7380 1988
rect 12412 2044 12708 2064
rect 12468 2042 12492 2044
rect 12548 2042 12572 2044
rect 12628 2042 12652 2044
rect 12490 1990 12492 2042
rect 12554 1990 12566 2042
rect 12628 1990 12630 2042
rect 12468 1988 12492 1990
rect 12548 1988 12572 1990
rect 12628 1988 12652 1990
rect 12412 1968 12708 1988
rect 17740 2044 18036 2064
rect 17796 2042 17820 2044
rect 17876 2042 17900 2044
rect 17956 2042 17980 2044
rect 17818 1990 17820 2042
rect 17882 1990 17894 2042
rect 17956 1990 17958 2042
rect 17796 1988 17820 1990
rect 17876 1988 17900 1990
rect 17956 1988 17980 1990
rect 17740 1968 18036 1988
rect 3856 1940 3908 1946
rect 3856 1882 3908 1888
rect 21612 1736 21664 1742
rect 21612 1678 21664 1684
rect 4420 1500 4716 1520
rect 4476 1498 4500 1500
rect 4556 1498 4580 1500
rect 4636 1498 4660 1500
rect 4498 1446 4500 1498
rect 4562 1446 4574 1498
rect 4636 1446 4638 1498
rect 4476 1444 4500 1446
rect 4556 1444 4580 1446
rect 4636 1444 4660 1446
rect 4420 1424 4716 1444
rect 9748 1500 10044 1520
rect 9804 1498 9828 1500
rect 9884 1498 9908 1500
rect 9964 1498 9988 1500
rect 9826 1446 9828 1498
rect 9890 1446 9902 1498
rect 9964 1446 9966 1498
rect 9804 1444 9828 1446
rect 9884 1444 9908 1446
rect 9964 1444 9988 1446
rect 9748 1424 10044 1444
rect 15076 1500 15372 1520
rect 15132 1498 15156 1500
rect 15212 1498 15236 1500
rect 15292 1498 15316 1500
rect 15154 1446 15156 1498
rect 15218 1446 15230 1498
rect 15292 1446 15294 1498
rect 15132 1444 15156 1446
rect 15212 1444 15236 1446
rect 15292 1444 15316 1446
rect 15076 1424 15372 1444
rect 20404 1500 20700 1520
rect 20460 1498 20484 1500
rect 20540 1498 20564 1500
rect 20620 1498 20644 1500
rect 20482 1446 20484 1498
rect 20546 1446 20558 1498
rect 20620 1446 20622 1498
rect 20460 1444 20484 1446
rect 20540 1444 20564 1446
rect 20620 1444 20644 1446
rect 20404 1424 20700 1444
rect 21624 1334 21652 1678
rect 21612 1328 21664 1334
rect 21612 1270 21664 1276
rect 2936 1192 2988 1198
rect 2290 1160 2346 1169
rect 2290 1095 2346 1104
rect 2934 1160 2936 1169
rect 2988 1160 2990 1169
rect 2934 1095 2990 1104
rect 7084 956 7380 976
rect 7140 954 7164 956
rect 7220 954 7244 956
rect 7300 954 7324 956
rect 7162 902 7164 954
rect 7226 902 7238 954
rect 7300 902 7302 954
rect 7140 900 7164 902
rect 7220 900 7244 902
rect 7300 900 7324 902
rect 7084 880 7380 900
rect 12412 956 12708 976
rect 12468 954 12492 956
rect 12548 954 12572 956
rect 12628 954 12652 956
rect 12490 902 12492 954
rect 12554 902 12566 954
rect 12628 902 12630 954
rect 12468 900 12492 902
rect 12548 900 12572 902
rect 12628 900 12652 902
rect 12412 880 12708 900
rect 17740 956 18036 976
rect 17796 954 17820 956
rect 17876 954 17900 956
rect 17956 954 17980 956
rect 17818 902 17820 954
rect 17882 902 17894 954
rect 17956 902 17958 954
rect 17796 900 17820 902
rect 17876 900 17900 902
rect 17956 900 17980 902
rect 17740 880 18036 900
<< via2 >>
rect 1922 22320 1978 22376
rect 4420 22170 4476 22172
rect 4500 22170 4556 22172
rect 4580 22170 4636 22172
rect 4660 22170 4716 22172
rect 4420 22118 4446 22170
rect 4446 22118 4476 22170
rect 4500 22118 4510 22170
rect 4510 22118 4556 22170
rect 4580 22118 4626 22170
rect 4626 22118 4636 22170
rect 4660 22118 4690 22170
rect 4690 22118 4716 22170
rect 4420 22116 4476 22118
rect 4500 22116 4556 22118
rect 4580 22116 4636 22118
rect 4660 22116 4716 22118
rect 9748 22170 9804 22172
rect 9828 22170 9884 22172
rect 9908 22170 9964 22172
rect 9988 22170 10044 22172
rect 9748 22118 9774 22170
rect 9774 22118 9804 22170
rect 9828 22118 9838 22170
rect 9838 22118 9884 22170
rect 9908 22118 9954 22170
rect 9954 22118 9964 22170
rect 9988 22118 10018 22170
rect 10018 22118 10044 22170
rect 9748 22116 9804 22118
rect 9828 22116 9884 22118
rect 9908 22116 9964 22118
rect 9988 22116 10044 22118
rect 15076 22170 15132 22172
rect 15156 22170 15212 22172
rect 15236 22170 15292 22172
rect 15316 22170 15372 22172
rect 15076 22118 15102 22170
rect 15102 22118 15132 22170
rect 15156 22118 15166 22170
rect 15166 22118 15212 22170
rect 15236 22118 15282 22170
rect 15282 22118 15292 22170
rect 15316 22118 15346 22170
rect 15346 22118 15372 22170
rect 15076 22116 15132 22118
rect 15156 22116 15212 22118
rect 15236 22116 15292 22118
rect 15316 22116 15372 22118
rect 20404 22170 20460 22172
rect 20484 22170 20540 22172
rect 20564 22170 20620 22172
rect 20644 22170 20700 22172
rect 20404 22118 20430 22170
rect 20430 22118 20460 22170
rect 20484 22118 20494 22170
rect 20494 22118 20540 22170
rect 20564 22118 20610 22170
rect 20610 22118 20620 22170
rect 20644 22118 20674 22170
rect 20674 22118 20700 22170
rect 20404 22116 20460 22118
rect 20484 22116 20540 22118
rect 20564 22116 20620 22118
rect 20644 22116 20700 22118
rect 2474 21812 2476 21832
rect 2476 21812 2528 21832
rect 2528 21812 2530 21832
rect 2474 21776 2530 21812
rect 7084 21626 7140 21628
rect 7164 21626 7220 21628
rect 7244 21626 7300 21628
rect 7324 21626 7380 21628
rect 7084 21574 7110 21626
rect 7110 21574 7140 21626
rect 7164 21574 7174 21626
rect 7174 21574 7220 21626
rect 7244 21574 7290 21626
rect 7290 21574 7300 21626
rect 7324 21574 7354 21626
rect 7354 21574 7380 21626
rect 7084 21572 7140 21574
rect 7164 21572 7220 21574
rect 7244 21572 7300 21574
rect 7324 21572 7380 21574
rect 12412 21626 12468 21628
rect 12492 21626 12548 21628
rect 12572 21626 12628 21628
rect 12652 21626 12708 21628
rect 12412 21574 12438 21626
rect 12438 21574 12468 21626
rect 12492 21574 12502 21626
rect 12502 21574 12548 21626
rect 12572 21574 12618 21626
rect 12618 21574 12628 21626
rect 12652 21574 12682 21626
rect 12682 21574 12708 21626
rect 12412 21572 12468 21574
rect 12492 21572 12548 21574
rect 12572 21572 12628 21574
rect 12652 21572 12708 21574
rect 17740 21626 17796 21628
rect 17820 21626 17876 21628
rect 17900 21626 17956 21628
rect 17980 21626 18036 21628
rect 17740 21574 17766 21626
rect 17766 21574 17796 21626
rect 17820 21574 17830 21626
rect 17830 21574 17876 21626
rect 17900 21574 17946 21626
rect 17946 21574 17956 21626
rect 17980 21574 18010 21626
rect 18010 21574 18036 21626
rect 17740 21572 17796 21574
rect 17820 21572 17876 21574
rect 17900 21572 17956 21574
rect 17980 21572 18036 21574
rect 2474 21232 2530 21288
rect 4420 21082 4476 21084
rect 4500 21082 4556 21084
rect 4580 21082 4636 21084
rect 4660 21082 4716 21084
rect 4420 21030 4446 21082
rect 4446 21030 4476 21082
rect 4500 21030 4510 21082
rect 4510 21030 4556 21082
rect 4580 21030 4626 21082
rect 4626 21030 4636 21082
rect 4660 21030 4690 21082
rect 4690 21030 4716 21082
rect 4420 21028 4476 21030
rect 4500 21028 4556 21030
rect 4580 21028 4636 21030
rect 4660 21028 4716 21030
rect 9748 21082 9804 21084
rect 9828 21082 9884 21084
rect 9908 21082 9964 21084
rect 9988 21082 10044 21084
rect 9748 21030 9774 21082
rect 9774 21030 9804 21082
rect 9828 21030 9838 21082
rect 9838 21030 9884 21082
rect 9908 21030 9954 21082
rect 9954 21030 9964 21082
rect 9988 21030 10018 21082
rect 10018 21030 10044 21082
rect 9748 21028 9804 21030
rect 9828 21028 9884 21030
rect 9908 21028 9964 21030
rect 9988 21028 10044 21030
rect 15076 21082 15132 21084
rect 15156 21082 15212 21084
rect 15236 21082 15292 21084
rect 15316 21082 15372 21084
rect 15076 21030 15102 21082
rect 15102 21030 15132 21082
rect 15156 21030 15166 21082
rect 15166 21030 15212 21082
rect 15236 21030 15282 21082
rect 15282 21030 15292 21082
rect 15316 21030 15346 21082
rect 15346 21030 15372 21082
rect 15076 21028 15132 21030
rect 15156 21028 15212 21030
rect 15236 21028 15292 21030
rect 15316 21028 15372 21030
rect 20404 21082 20460 21084
rect 20484 21082 20540 21084
rect 20564 21082 20620 21084
rect 20644 21082 20700 21084
rect 20404 21030 20430 21082
rect 20430 21030 20460 21082
rect 20484 21030 20494 21082
rect 20494 21030 20540 21082
rect 20564 21030 20610 21082
rect 20610 21030 20620 21082
rect 20644 21030 20674 21082
rect 20674 21030 20700 21082
rect 20404 21028 20460 21030
rect 20484 21028 20540 21030
rect 20564 21028 20620 21030
rect 20644 21028 20700 21030
rect 7084 20538 7140 20540
rect 7164 20538 7220 20540
rect 7244 20538 7300 20540
rect 7324 20538 7380 20540
rect 7084 20486 7110 20538
rect 7110 20486 7140 20538
rect 7164 20486 7174 20538
rect 7174 20486 7220 20538
rect 7244 20486 7290 20538
rect 7290 20486 7300 20538
rect 7324 20486 7354 20538
rect 7354 20486 7380 20538
rect 7084 20484 7140 20486
rect 7164 20484 7220 20486
rect 7244 20484 7300 20486
rect 7324 20484 7380 20486
rect 12412 20538 12468 20540
rect 12492 20538 12548 20540
rect 12572 20538 12628 20540
rect 12652 20538 12708 20540
rect 12412 20486 12438 20538
rect 12438 20486 12468 20538
rect 12492 20486 12502 20538
rect 12502 20486 12548 20538
rect 12572 20486 12618 20538
rect 12618 20486 12628 20538
rect 12652 20486 12682 20538
rect 12682 20486 12708 20538
rect 12412 20484 12468 20486
rect 12492 20484 12548 20486
rect 12572 20484 12628 20486
rect 12652 20484 12708 20486
rect 17740 20538 17796 20540
rect 17820 20538 17876 20540
rect 17900 20538 17956 20540
rect 17980 20538 18036 20540
rect 17740 20486 17766 20538
rect 17766 20486 17796 20538
rect 17820 20486 17830 20538
rect 17830 20486 17876 20538
rect 17900 20486 17946 20538
rect 17946 20486 17956 20538
rect 17980 20486 18010 20538
rect 18010 20486 18036 20538
rect 17740 20484 17796 20486
rect 17820 20484 17876 20486
rect 17900 20484 17956 20486
rect 17980 20484 18036 20486
rect 2474 20144 2530 20200
rect 4420 19994 4476 19996
rect 4500 19994 4556 19996
rect 4580 19994 4636 19996
rect 4660 19994 4716 19996
rect 4420 19942 4446 19994
rect 4446 19942 4476 19994
rect 4500 19942 4510 19994
rect 4510 19942 4556 19994
rect 4580 19942 4626 19994
rect 4626 19942 4636 19994
rect 4660 19942 4690 19994
rect 4690 19942 4716 19994
rect 4420 19940 4476 19942
rect 4500 19940 4556 19942
rect 4580 19940 4636 19942
rect 4660 19940 4716 19942
rect 9748 19994 9804 19996
rect 9828 19994 9884 19996
rect 9908 19994 9964 19996
rect 9988 19994 10044 19996
rect 9748 19942 9774 19994
rect 9774 19942 9804 19994
rect 9828 19942 9838 19994
rect 9838 19942 9884 19994
rect 9908 19942 9954 19994
rect 9954 19942 9964 19994
rect 9988 19942 10018 19994
rect 10018 19942 10044 19994
rect 9748 19940 9804 19942
rect 9828 19940 9884 19942
rect 9908 19940 9964 19942
rect 9988 19940 10044 19942
rect 15076 19994 15132 19996
rect 15156 19994 15212 19996
rect 15236 19994 15292 19996
rect 15316 19994 15372 19996
rect 15076 19942 15102 19994
rect 15102 19942 15132 19994
rect 15156 19942 15166 19994
rect 15166 19942 15212 19994
rect 15236 19942 15282 19994
rect 15282 19942 15292 19994
rect 15316 19942 15346 19994
rect 15346 19942 15372 19994
rect 15076 19940 15132 19942
rect 15156 19940 15212 19942
rect 15236 19940 15292 19942
rect 15316 19940 15372 19942
rect 20404 19994 20460 19996
rect 20484 19994 20540 19996
rect 20564 19994 20620 19996
rect 20644 19994 20700 19996
rect 20404 19942 20430 19994
rect 20430 19942 20460 19994
rect 20484 19942 20494 19994
rect 20494 19942 20540 19994
rect 20564 19942 20610 19994
rect 20610 19942 20620 19994
rect 20644 19942 20674 19994
rect 20674 19942 20700 19994
rect 20404 19940 20460 19942
rect 20484 19940 20540 19942
rect 20564 19940 20620 19942
rect 20644 19940 20700 19942
rect 7084 19450 7140 19452
rect 7164 19450 7220 19452
rect 7244 19450 7300 19452
rect 7324 19450 7380 19452
rect 7084 19398 7110 19450
rect 7110 19398 7140 19450
rect 7164 19398 7174 19450
rect 7174 19398 7220 19450
rect 7244 19398 7290 19450
rect 7290 19398 7300 19450
rect 7324 19398 7354 19450
rect 7354 19398 7380 19450
rect 7084 19396 7140 19398
rect 7164 19396 7220 19398
rect 7244 19396 7300 19398
rect 7324 19396 7380 19398
rect 12412 19450 12468 19452
rect 12492 19450 12548 19452
rect 12572 19450 12628 19452
rect 12652 19450 12708 19452
rect 12412 19398 12438 19450
rect 12438 19398 12468 19450
rect 12492 19398 12502 19450
rect 12502 19398 12548 19450
rect 12572 19398 12618 19450
rect 12618 19398 12628 19450
rect 12652 19398 12682 19450
rect 12682 19398 12708 19450
rect 12412 19396 12468 19398
rect 12492 19396 12548 19398
rect 12572 19396 12628 19398
rect 12652 19396 12708 19398
rect 17740 19450 17796 19452
rect 17820 19450 17876 19452
rect 17900 19450 17956 19452
rect 17980 19450 18036 19452
rect 17740 19398 17766 19450
rect 17766 19398 17796 19450
rect 17820 19398 17830 19450
rect 17830 19398 17876 19450
rect 17900 19398 17946 19450
rect 17946 19398 17956 19450
rect 17980 19398 18010 19450
rect 18010 19398 18036 19450
rect 17740 19396 17796 19398
rect 17820 19396 17876 19398
rect 17900 19396 17956 19398
rect 17980 19396 18036 19398
rect 2474 19056 2530 19112
rect 4420 18906 4476 18908
rect 4500 18906 4556 18908
rect 4580 18906 4636 18908
rect 4660 18906 4716 18908
rect 4420 18854 4446 18906
rect 4446 18854 4476 18906
rect 4500 18854 4510 18906
rect 4510 18854 4556 18906
rect 4580 18854 4626 18906
rect 4626 18854 4636 18906
rect 4660 18854 4690 18906
rect 4690 18854 4716 18906
rect 4420 18852 4476 18854
rect 4500 18852 4556 18854
rect 4580 18852 4636 18854
rect 4660 18852 4716 18854
rect 9748 18906 9804 18908
rect 9828 18906 9884 18908
rect 9908 18906 9964 18908
rect 9988 18906 10044 18908
rect 9748 18854 9774 18906
rect 9774 18854 9804 18906
rect 9828 18854 9838 18906
rect 9838 18854 9884 18906
rect 9908 18854 9954 18906
rect 9954 18854 9964 18906
rect 9988 18854 10018 18906
rect 10018 18854 10044 18906
rect 9748 18852 9804 18854
rect 9828 18852 9884 18854
rect 9908 18852 9964 18854
rect 9988 18852 10044 18854
rect 15076 18906 15132 18908
rect 15156 18906 15212 18908
rect 15236 18906 15292 18908
rect 15316 18906 15372 18908
rect 15076 18854 15102 18906
rect 15102 18854 15132 18906
rect 15156 18854 15166 18906
rect 15166 18854 15212 18906
rect 15236 18854 15282 18906
rect 15282 18854 15292 18906
rect 15316 18854 15346 18906
rect 15346 18854 15372 18906
rect 15076 18852 15132 18854
rect 15156 18852 15212 18854
rect 15236 18852 15292 18854
rect 15316 18852 15372 18854
rect 20404 18906 20460 18908
rect 20484 18906 20540 18908
rect 20564 18906 20620 18908
rect 20644 18906 20700 18908
rect 20404 18854 20430 18906
rect 20430 18854 20460 18906
rect 20484 18854 20494 18906
rect 20494 18854 20540 18906
rect 20564 18854 20610 18906
rect 20610 18854 20620 18906
rect 20644 18854 20674 18906
rect 20674 18854 20700 18906
rect 20404 18852 20460 18854
rect 20484 18852 20540 18854
rect 20564 18852 20620 18854
rect 20644 18852 20700 18854
rect 7084 18362 7140 18364
rect 7164 18362 7220 18364
rect 7244 18362 7300 18364
rect 7324 18362 7380 18364
rect 7084 18310 7110 18362
rect 7110 18310 7140 18362
rect 7164 18310 7174 18362
rect 7174 18310 7220 18362
rect 7244 18310 7290 18362
rect 7290 18310 7300 18362
rect 7324 18310 7354 18362
rect 7354 18310 7380 18362
rect 7084 18308 7140 18310
rect 7164 18308 7220 18310
rect 7244 18308 7300 18310
rect 7324 18308 7380 18310
rect 12412 18362 12468 18364
rect 12492 18362 12548 18364
rect 12572 18362 12628 18364
rect 12652 18362 12708 18364
rect 12412 18310 12438 18362
rect 12438 18310 12468 18362
rect 12492 18310 12502 18362
rect 12502 18310 12548 18362
rect 12572 18310 12618 18362
rect 12618 18310 12628 18362
rect 12652 18310 12682 18362
rect 12682 18310 12708 18362
rect 12412 18308 12468 18310
rect 12492 18308 12548 18310
rect 12572 18308 12628 18310
rect 12652 18308 12708 18310
rect 17740 18362 17796 18364
rect 17820 18362 17876 18364
rect 17900 18362 17956 18364
rect 17980 18362 18036 18364
rect 17740 18310 17766 18362
rect 17766 18310 17796 18362
rect 17820 18310 17830 18362
rect 17830 18310 17876 18362
rect 17900 18310 17946 18362
rect 17946 18310 17956 18362
rect 17980 18310 18010 18362
rect 18010 18310 18036 18362
rect 17740 18308 17796 18310
rect 17820 18308 17876 18310
rect 17900 18308 17956 18310
rect 17980 18308 18036 18310
rect 2474 17968 2530 18024
rect 4420 17818 4476 17820
rect 4500 17818 4556 17820
rect 4580 17818 4636 17820
rect 4660 17818 4716 17820
rect 4420 17766 4446 17818
rect 4446 17766 4476 17818
rect 4500 17766 4510 17818
rect 4510 17766 4556 17818
rect 4580 17766 4626 17818
rect 4626 17766 4636 17818
rect 4660 17766 4690 17818
rect 4690 17766 4716 17818
rect 4420 17764 4476 17766
rect 4500 17764 4556 17766
rect 4580 17764 4636 17766
rect 4660 17764 4716 17766
rect 9748 17818 9804 17820
rect 9828 17818 9884 17820
rect 9908 17818 9964 17820
rect 9988 17818 10044 17820
rect 9748 17766 9774 17818
rect 9774 17766 9804 17818
rect 9828 17766 9838 17818
rect 9838 17766 9884 17818
rect 9908 17766 9954 17818
rect 9954 17766 9964 17818
rect 9988 17766 10018 17818
rect 10018 17766 10044 17818
rect 9748 17764 9804 17766
rect 9828 17764 9884 17766
rect 9908 17764 9964 17766
rect 9988 17764 10044 17766
rect 15076 17818 15132 17820
rect 15156 17818 15212 17820
rect 15236 17818 15292 17820
rect 15316 17818 15372 17820
rect 15076 17766 15102 17818
rect 15102 17766 15132 17818
rect 15156 17766 15166 17818
rect 15166 17766 15212 17818
rect 15236 17766 15282 17818
rect 15282 17766 15292 17818
rect 15316 17766 15346 17818
rect 15346 17766 15372 17818
rect 15076 17764 15132 17766
rect 15156 17764 15212 17766
rect 15236 17764 15292 17766
rect 15316 17764 15372 17766
rect 20404 17818 20460 17820
rect 20484 17818 20540 17820
rect 20564 17818 20620 17820
rect 20644 17818 20700 17820
rect 20404 17766 20430 17818
rect 20430 17766 20460 17818
rect 20484 17766 20494 17818
rect 20494 17766 20540 17818
rect 20564 17766 20610 17818
rect 20610 17766 20620 17818
rect 20644 17766 20674 17818
rect 20674 17766 20700 17818
rect 20404 17764 20460 17766
rect 20484 17764 20540 17766
rect 20564 17764 20620 17766
rect 20644 17764 20700 17766
rect 7084 17274 7140 17276
rect 7164 17274 7220 17276
rect 7244 17274 7300 17276
rect 7324 17274 7380 17276
rect 7084 17222 7110 17274
rect 7110 17222 7140 17274
rect 7164 17222 7174 17274
rect 7174 17222 7220 17274
rect 7244 17222 7290 17274
rect 7290 17222 7300 17274
rect 7324 17222 7354 17274
rect 7354 17222 7380 17274
rect 7084 17220 7140 17222
rect 7164 17220 7220 17222
rect 7244 17220 7300 17222
rect 7324 17220 7380 17222
rect 12412 17274 12468 17276
rect 12492 17274 12548 17276
rect 12572 17274 12628 17276
rect 12652 17274 12708 17276
rect 12412 17222 12438 17274
rect 12438 17222 12468 17274
rect 12492 17222 12502 17274
rect 12502 17222 12548 17274
rect 12572 17222 12618 17274
rect 12618 17222 12628 17274
rect 12652 17222 12682 17274
rect 12682 17222 12708 17274
rect 12412 17220 12468 17222
rect 12492 17220 12548 17222
rect 12572 17220 12628 17222
rect 12652 17220 12708 17222
rect 17740 17274 17796 17276
rect 17820 17274 17876 17276
rect 17900 17274 17956 17276
rect 17980 17274 18036 17276
rect 17740 17222 17766 17274
rect 17766 17222 17796 17274
rect 17820 17222 17830 17274
rect 17830 17222 17876 17274
rect 17900 17222 17946 17274
rect 17946 17222 17956 17274
rect 17980 17222 18010 17274
rect 18010 17222 18036 17274
rect 17740 17220 17796 17222
rect 17820 17220 17876 17222
rect 17900 17220 17956 17222
rect 17980 17220 18036 17222
rect 4420 16730 4476 16732
rect 4500 16730 4556 16732
rect 4580 16730 4636 16732
rect 4660 16730 4716 16732
rect 4420 16678 4446 16730
rect 4446 16678 4476 16730
rect 4500 16678 4510 16730
rect 4510 16678 4556 16730
rect 4580 16678 4626 16730
rect 4626 16678 4636 16730
rect 4660 16678 4690 16730
rect 4690 16678 4716 16730
rect 4420 16676 4476 16678
rect 4500 16676 4556 16678
rect 4580 16676 4636 16678
rect 4660 16676 4716 16678
rect 9748 16730 9804 16732
rect 9828 16730 9884 16732
rect 9908 16730 9964 16732
rect 9988 16730 10044 16732
rect 9748 16678 9774 16730
rect 9774 16678 9804 16730
rect 9828 16678 9838 16730
rect 9838 16678 9884 16730
rect 9908 16678 9954 16730
rect 9954 16678 9964 16730
rect 9988 16678 10018 16730
rect 10018 16678 10044 16730
rect 9748 16676 9804 16678
rect 9828 16676 9884 16678
rect 9908 16676 9964 16678
rect 9988 16676 10044 16678
rect 15076 16730 15132 16732
rect 15156 16730 15212 16732
rect 15236 16730 15292 16732
rect 15316 16730 15372 16732
rect 15076 16678 15102 16730
rect 15102 16678 15132 16730
rect 15156 16678 15166 16730
rect 15166 16678 15212 16730
rect 15236 16678 15282 16730
rect 15282 16678 15292 16730
rect 15316 16678 15346 16730
rect 15346 16678 15372 16730
rect 15076 16676 15132 16678
rect 15156 16676 15212 16678
rect 15236 16676 15292 16678
rect 15316 16676 15372 16678
rect 20404 16730 20460 16732
rect 20484 16730 20540 16732
rect 20564 16730 20620 16732
rect 20644 16730 20700 16732
rect 20404 16678 20430 16730
rect 20430 16678 20460 16730
rect 20484 16678 20494 16730
rect 20494 16678 20540 16730
rect 20564 16678 20610 16730
rect 20610 16678 20620 16730
rect 20644 16678 20674 16730
rect 20674 16678 20700 16730
rect 20404 16676 20460 16678
rect 20484 16676 20540 16678
rect 20564 16676 20620 16678
rect 20644 16676 20700 16678
rect 2474 16336 2530 16392
rect 7084 16186 7140 16188
rect 7164 16186 7220 16188
rect 7244 16186 7300 16188
rect 7324 16186 7380 16188
rect 7084 16134 7110 16186
rect 7110 16134 7140 16186
rect 7164 16134 7174 16186
rect 7174 16134 7220 16186
rect 7244 16134 7290 16186
rect 7290 16134 7300 16186
rect 7324 16134 7354 16186
rect 7354 16134 7380 16186
rect 7084 16132 7140 16134
rect 7164 16132 7220 16134
rect 7244 16132 7300 16134
rect 7324 16132 7380 16134
rect 12412 16186 12468 16188
rect 12492 16186 12548 16188
rect 12572 16186 12628 16188
rect 12652 16186 12708 16188
rect 12412 16134 12438 16186
rect 12438 16134 12468 16186
rect 12492 16134 12502 16186
rect 12502 16134 12548 16186
rect 12572 16134 12618 16186
rect 12618 16134 12628 16186
rect 12652 16134 12682 16186
rect 12682 16134 12708 16186
rect 12412 16132 12468 16134
rect 12492 16132 12548 16134
rect 12572 16132 12628 16134
rect 12652 16132 12708 16134
rect 17740 16186 17796 16188
rect 17820 16186 17876 16188
rect 17900 16186 17956 16188
rect 17980 16186 18036 16188
rect 17740 16134 17766 16186
rect 17766 16134 17796 16186
rect 17820 16134 17830 16186
rect 17830 16134 17876 16186
rect 17900 16134 17946 16186
rect 17946 16134 17956 16186
rect 17980 16134 18010 16186
rect 18010 16134 18036 16186
rect 17740 16132 17796 16134
rect 17820 16132 17876 16134
rect 17900 16132 17956 16134
rect 17980 16132 18036 16134
rect 2474 15792 2530 15848
rect 4420 15642 4476 15644
rect 4500 15642 4556 15644
rect 4580 15642 4636 15644
rect 4660 15642 4716 15644
rect 4420 15590 4446 15642
rect 4446 15590 4476 15642
rect 4500 15590 4510 15642
rect 4510 15590 4556 15642
rect 4580 15590 4626 15642
rect 4626 15590 4636 15642
rect 4660 15590 4690 15642
rect 4690 15590 4716 15642
rect 4420 15588 4476 15590
rect 4500 15588 4556 15590
rect 4580 15588 4636 15590
rect 4660 15588 4716 15590
rect 9748 15642 9804 15644
rect 9828 15642 9884 15644
rect 9908 15642 9964 15644
rect 9988 15642 10044 15644
rect 9748 15590 9774 15642
rect 9774 15590 9804 15642
rect 9828 15590 9838 15642
rect 9838 15590 9884 15642
rect 9908 15590 9954 15642
rect 9954 15590 9964 15642
rect 9988 15590 10018 15642
rect 10018 15590 10044 15642
rect 9748 15588 9804 15590
rect 9828 15588 9884 15590
rect 9908 15588 9964 15590
rect 9988 15588 10044 15590
rect 15076 15642 15132 15644
rect 15156 15642 15212 15644
rect 15236 15642 15292 15644
rect 15316 15642 15372 15644
rect 15076 15590 15102 15642
rect 15102 15590 15132 15642
rect 15156 15590 15166 15642
rect 15166 15590 15212 15642
rect 15236 15590 15282 15642
rect 15282 15590 15292 15642
rect 15316 15590 15346 15642
rect 15346 15590 15372 15642
rect 15076 15588 15132 15590
rect 15156 15588 15212 15590
rect 15236 15588 15292 15590
rect 15316 15588 15372 15590
rect 20404 15642 20460 15644
rect 20484 15642 20540 15644
rect 20564 15642 20620 15644
rect 20644 15642 20700 15644
rect 20404 15590 20430 15642
rect 20430 15590 20460 15642
rect 20484 15590 20494 15642
rect 20494 15590 20540 15642
rect 20564 15590 20610 15642
rect 20610 15590 20620 15642
rect 20644 15590 20674 15642
rect 20674 15590 20700 15642
rect 20404 15588 20460 15590
rect 20484 15588 20540 15590
rect 20564 15588 20620 15590
rect 20644 15588 20700 15590
rect 7084 15098 7140 15100
rect 7164 15098 7220 15100
rect 7244 15098 7300 15100
rect 7324 15098 7380 15100
rect 7084 15046 7110 15098
rect 7110 15046 7140 15098
rect 7164 15046 7174 15098
rect 7174 15046 7220 15098
rect 7244 15046 7290 15098
rect 7290 15046 7300 15098
rect 7324 15046 7354 15098
rect 7354 15046 7380 15098
rect 7084 15044 7140 15046
rect 7164 15044 7220 15046
rect 7244 15044 7300 15046
rect 7324 15044 7380 15046
rect 12412 15098 12468 15100
rect 12492 15098 12548 15100
rect 12572 15098 12628 15100
rect 12652 15098 12708 15100
rect 12412 15046 12438 15098
rect 12438 15046 12468 15098
rect 12492 15046 12502 15098
rect 12502 15046 12548 15098
rect 12572 15046 12618 15098
rect 12618 15046 12628 15098
rect 12652 15046 12682 15098
rect 12682 15046 12708 15098
rect 12412 15044 12468 15046
rect 12492 15044 12548 15046
rect 12572 15044 12628 15046
rect 12652 15044 12708 15046
rect 17740 15098 17796 15100
rect 17820 15098 17876 15100
rect 17900 15098 17956 15100
rect 17980 15098 18036 15100
rect 17740 15046 17766 15098
rect 17766 15046 17796 15098
rect 17820 15046 17830 15098
rect 17830 15046 17876 15098
rect 17900 15046 17946 15098
rect 17946 15046 17956 15098
rect 17980 15046 18010 15098
rect 18010 15046 18036 15098
rect 17740 15044 17796 15046
rect 17820 15044 17876 15046
rect 17900 15044 17956 15046
rect 17980 15044 18036 15046
rect 4420 14554 4476 14556
rect 4500 14554 4556 14556
rect 4580 14554 4636 14556
rect 4660 14554 4716 14556
rect 4420 14502 4446 14554
rect 4446 14502 4476 14554
rect 4500 14502 4510 14554
rect 4510 14502 4556 14554
rect 4580 14502 4626 14554
rect 4626 14502 4636 14554
rect 4660 14502 4690 14554
rect 4690 14502 4716 14554
rect 4420 14500 4476 14502
rect 4500 14500 4556 14502
rect 4580 14500 4636 14502
rect 4660 14500 4716 14502
rect 9748 14554 9804 14556
rect 9828 14554 9884 14556
rect 9908 14554 9964 14556
rect 9988 14554 10044 14556
rect 9748 14502 9774 14554
rect 9774 14502 9804 14554
rect 9828 14502 9838 14554
rect 9838 14502 9884 14554
rect 9908 14502 9954 14554
rect 9954 14502 9964 14554
rect 9988 14502 10018 14554
rect 10018 14502 10044 14554
rect 9748 14500 9804 14502
rect 9828 14500 9884 14502
rect 9908 14500 9964 14502
rect 9988 14500 10044 14502
rect 15076 14554 15132 14556
rect 15156 14554 15212 14556
rect 15236 14554 15292 14556
rect 15316 14554 15372 14556
rect 15076 14502 15102 14554
rect 15102 14502 15132 14554
rect 15156 14502 15166 14554
rect 15166 14502 15212 14554
rect 15236 14502 15282 14554
rect 15282 14502 15292 14554
rect 15316 14502 15346 14554
rect 15346 14502 15372 14554
rect 15076 14500 15132 14502
rect 15156 14500 15212 14502
rect 15236 14500 15292 14502
rect 15316 14500 15372 14502
rect 20404 14554 20460 14556
rect 20484 14554 20540 14556
rect 20564 14554 20620 14556
rect 20644 14554 20700 14556
rect 20404 14502 20430 14554
rect 20430 14502 20460 14554
rect 20484 14502 20494 14554
rect 20494 14502 20540 14554
rect 20564 14502 20610 14554
rect 20610 14502 20620 14554
rect 20644 14502 20674 14554
rect 20674 14502 20700 14554
rect 20404 14500 20460 14502
rect 20484 14500 20540 14502
rect 20564 14500 20620 14502
rect 20644 14500 20700 14502
rect 7084 14010 7140 14012
rect 7164 14010 7220 14012
rect 7244 14010 7300 14012
rect 7324 14010 7380 14012
rect 7084 13958 7110 14010
rect 7110 13958 7140 14010
rect 7164 13958 7174 14010
rect 7174 13958 7220 14010
rect 7244 13958 7290 14010
rect 7290 13958 7300 14010
rect 7324 13958 7354 14010
rect 7354 13958 7380 14010
rect 7084 13956 7140 13958
rect 7164 13956 7220 13958
rect 7244 13956 7300 13958
rect 7324 13956 7380 13958
rect 12412 14010 12468 14012
rect 12492 14010 12548 14012
rect 12572 14010 12628 14012
rect 12652 14010 12708 14012
rect 12412 13958 12438 14010
rect 12438 13958 12468 14010
rect 12492 13958 12502 14010
rect 12502 13958 12548 14010
rect 12572 13958 12618 14010
rect 12618 13958 12628 14010
rect 12652 13958 12682 14010
rect 12682 13958 12708 14010
rect 12412 13956 12468 13958
rect 12492 13956 12548 13958
rect 12572 13956 12628 13958
rect 12652 13956 12708 13958
rect 17740 14010 17796 14012
rect 17820 14010 17876 14012
rect 17900 14010 17956 14012
rect 17980 14010 18036 14012
rect 17740 13958 17766 14010
rect 17766 13958 17796 14010
rect 17820 13958 17830 14010
rect 17830 13958 17876 14010
rect 17900 13958 17946 14010
rect 17946 13958 17956 14010
rect 17980 13958 18010 14010
rect 18010 13958 18036 14010
rect 17740 13956 17796 13958
rect 17820 13956 17876 13958
rect 17900 13956 17956 13958
rect 17980 13956 18036 13958
rect 2474 13616 2530 13672
rect 4420 13466 4476 13468
rect 4500 13466 4556 13468
rect 4580 13466 4636 13468
rect 4660 13466 4716 13468
rect 4420 13414 4446 13466
rect 4446 13414 4476 13466
rect 4500 13414 4510 13466
rect 4510 13414 4556 13466
rect 4580 13414 4626 13466
rect 4626 13414 4636 13466
rect 4660 13414 4690 13466
rect 4690 13414 4716 13466
rect 4420 13412 4476 13414
rect 4500 13412 4556 13414
rect 4580 13412 4636 13414
rect 4660 13412 4716 13414
rect 9748 13466 9804 13468
rect 9828 13466 9884 13468
rect 9908 13466 9964 13468
rect 9988 13466 10044 13468
rect 9748 13414 9774 13466
rect 9774 13414 9804 13466
rect 9828 13414 9838 13466
rect 9838 13414 9884 13466
rect 9908 13414 9954 13466
rect 9954 13414 9964 13466
rect 9988 13414 10018 13466
rect 10018 13414 10044 13466
rect 9748 13412 9804 13414
rect 9828 13412 9884 13414
rect 9908 13412 9964 13414
rect 9988 13412 10044 13414
rect 15076 13466 15132 13468
rect 15156 13466 15212 13468
rect 15236 13466 15292 13468
rect 15316 13466 15372 13468
rect 15076 13414 15102 13466
rect 15102 13414 15132 13466
rect 15156 13414 15166 13466
rect 15166 13414 15212 13466
rect 15236 13414 15282 13466
rect 15282 13414 15292 13466
rect 15316 13414 15346 13466
rect 15346 13414 15372 13466
rect 15076 13412 15132 13414
rect 15156 13412 15212 13414
rect 15236 13412 15292 13414
rect 15316 13412 15372 13414
rect 20404 13466 20460 13468
rect 20484 13466 20540 13468
rect 20564 13466 20620 13468
rect 20644 13466 20700 13468
rect 20404 13414 20430 13466
rect 20430 13414 20460 13466
rect 20484 13414 20494 13466
rect 20494 13414 20540 13466
rect 20564 13414 20610 13466
rect 20610 13414 20620 13466
rect 20644 13414 20674 13466
rect 20674 13414 20700 13466
rect 20404 13412 20460 13414
rect 20484 13412 20540 13414
rect 20564 13412 20620 13414
rect 20644 13412 20700 13414
rect 7084 12922 7140 12924
rect 7164 12922 7220 12924
rect 7244 12922 7300 12924
rect 7324 12922 7380 12924
rect 7084 12870 7110 12922
rect 7110 12870 7140 12922
rect 7164 12870 7174 12922
rect 7174 12870 7220 12922
rect 7244 12870 7290 12922
rect 7290 12870 7300 12922
rect 7324 12870 7354 12922
rect 7354 12870 7380 12922
rect 7084 12868 7140 12870
rect 7164 12868 7220 12870
rect 7244 12868 7300 12870
rect 7324 12868 7380 12870
rect 12412 12922 12468 12924
rect 12492 12922 12548 12924
rect 12572 12922 12628 12924
rect 12652 12922 12708 12924
rect 12412 12870 12438 12922
rect 12438 12870 12468 12922
rect 12492 12870 12502 12922
rect 12502 12870 12548 12922
rect 12572 12870 12618 12922
rect 12618 12870 12628 12922
rect 12652 12870 12682 12922
rect 12682 12870 12708 12922
rect 12412 12868 12468 12870
rect 12492 12868 12548 12870
rect 12572 12868 12628 12870
rect 12652 12868 12708 12870
rect 17740 12922 17796 12924
rect 17820 12922 17876 12924
rect 17900 12922 17956 12924
rect 17980 12922 18036 12924
rect 17740 12870 17766 12922
rect 17766 12870 17796 12922
rect 17820 12870 17830 12922
rect 17830 12870 17876 12922
rect 17900 12870 17946 12922
rect 17946 12870 17956 12922
rect 17980 12870 18010 12922
rect 18010 12870 18036 12922
rect 17740 12868 17796 12870
rect 17820 12868 17876 12870
rect 17900 12868 17956 12870
rect 17980 12868 18036 12870
rect 4420 12378 4476 12380
rect 4500 12378 4556 12380
rect 4580 12378 4636 12380
rect 4660 12378 4716 12380
rect 4420 12326 4446 12378
rect 4446 12326 4476 12378
rect 4500 12326 4510 12378
rect 4510 12326 4556 12378
rect 4580 12326 4626 12378
rect 4626 12326 4636 12378
rect 4660 12326 4690 12378
rect 4690 12326 4716 12378
rect 4420 12324 4476 12326
rect 4500 12324 4556 12326
rect 4580 12324 4636 12326
rect 4660 12324 4716 12326
rect 9748 12378 9804 12380
rect 9828 12378 9884 12380
rect 9908 12378 9964 12380
rect 9988 12378 10044 12380
rect 9748 12326 9774 12378
rect 9774 12326 9804 12378
rect 9828 12326 9838 12378
rect 9838 12326 9884 12378
rect 9908 12326 9954 12378
rect 9954 12326 9964 12378
rect 9988 12326 10018 12378
rect 10018 12326 10044 12378
rect 9748 12324 9804 12326
rect 9828 12324 9884 12326
rect 9908 12324 9964 12326
rect 9988 12324 10044 12326
rect 15076 12378 15132 12380
rect 15156 12378 15212 12380
rect 15236 12378 15292 12380
rect 15316 12378 15372 12380
rect 15076 12326 15102 12378
rect 15102 12326 15132 12378
rect 15156 12326 15166 12378
rect 15166 12326 15212 12378
rect 15236 12326 15282 12378
rect 15282 12326 15292 12378
rect 15316 12326 15346 12378
rect 15346 12326 15372 12378
rect 15076 12324 15132 12326
rect 15156 12324 15212 12326
rect 15236 12324 15292 12326
rect 15316 12324 15372 12326
rect 20404 12378 20460 12380
rect 20484 12378 20540 12380
rect 20564 12378 20620 12380
rect 20644 12378 20700 12380
rect 20404 12326 20430 12378
rect 20430 12326 20460 12378
rect 20484 12326 20494 12378
rect 20494 12326 20540 12378
rect 20564 12326 20610 12378
rect 20610 12326 20620 12378
rect 20644 12326 20674 12378
rect 20674 12326 20700 12378
rect 20404 12324 20460 12326
rect 20484 12324 20540 12326
rect 20564 12324 20620 12326
rect 20644 12324 20700 12326
rect 7084 11834 7140 11836
rect 7164 11834 7220 11836
rect 7244 11834 7300 11836
rect 7324 11834 7380 11836
rect 7084 11782 7110 11834
rect 7110 11782 7140 11834
rect 7164 11782 7174 11834
rect 7174 11782 7220 11834
rect 7244 11782 7290 11834
rect 7290 11782 7300 11834
rect 7324 11782 7354 11834
rect 7354 11782 7380 11834
rect 7084 11780 7140 11782
rect 7164 11780 7220 11782
rect 7244 11780 7300 11782
rect 7324 11780 7380 11782
rect 12412 11834 12468 11836
rect 12492 11834 12548 11836
rect 12572 11834 12628 11836
rect 12652 11834 12708 11836
rect 12412 11782 12438 11834
rect 12438 11782 12468 11834
rect 12492 11782 12502 11834
rect 12502 11782 12548 11834
rect 12572 11782 12618 11834
rect 12618 11782 12628 11834
rect 12652 11782 12682 11834
rect 12682 11782 12708 11834
rect 12412 11780 12468 11782
rect 12492 11780 12548 11782
rect 12572 11780 12628 11782
rect 12652 11780 12708 11782
rect 17740 11834 17796 11836
rect 17820 11834 17876 11836
rect 17900 11834 17956 11836
rect 17980 11834 18036 11836
rect 17740 11782 17766 11834
rect 17766 11782 17796 11834
rect 17820 11782 17830 11834
rect 17830 11782 17876 11834
rect 17900 11782 17946 11834
rect 17946 11782 17956 11834
rect 17980 11782 18010 11834
rect 18010 11782 18036 11834
rect 17740 11780 17796 11782
rect 17820 11780 17876 11782
rect 17900 11780 17956 11782
rect 17980 11780 18036 11782
rect 4420 11290 4476 11292
rect 4500 11290 4556 11292
rect 4580 11290 4636 11292
rect 4660 11290 4716 11292
rect 4420 11238 4446 11290
rect 4446 11238 4476 11290
rect 4500 11238 4510 11290
rect 4510 11238 4556 11290
rect 4580 11238 4626 11290
rect 4626 11238 4636 11290
rect 4660 11238 4690 11290
rect 4690 11238 4716 11290
rect 4420 11236 4476 11238
rect 4500 11236 4556 11238
rect 4580 11236 4636 11238
rect 4660 11236 4716 11238
rect 9748 11290 9804 11292
rect 9828 11290 9884 11292
rect 9908 11290 9964 11292
rect 9988 11290 10044 11292
rect 9748 11238 9774 11290
rect 9774 11238 9804 11290
rect 9828 11238 9838 11290
rect 9838 11238 9884 11290
rect 9908 11238 9954 11290
rect 9954 11238 9964 11290
rect 9988 11238 10018 11290
rect 10018 11238 10044 11290
rect 9748 11236 9804 11238
rect 9828 11236 9884 11238
rect 9908 11236 9964 11238
rect 9988 11236 10044 11238
rect 15076 11290 15132 11292
rect 15156 11290 15212 11292
rect 15236 11290 15292 11292
rect 15316 11290 15372 11292
rect 15076 11238 15102 11290
rect 15102 11238 15132 11290
rect 15156 11238 15166 11290
rect 15166 11238 15212 11290
rect 15236 11238 15282 11290
rect 15282 11238 15292 11290
rect 15316 11238 15346 11290
rect 15346 11238 15372 11290
rect 15076 11236 15132 11238
rect 15156 11236 15212 11238
rect 15236 11236 15292 11238
rect 15316 11236 15372 11238
rect 20404 11290 20460 11292
rect 20484 11290 20540 11292
rect 20564 11290 20620 11292
rect 20644 11290 20700 11292
rect 20404 11238 20430 11290
rect 20430 11238 20460 11290
rect 20484 11238 20494 11290
rect 20494 11238 20540 11290
rect 20564 11238 20610 11290
rect 20610 11238 20620 11290
rect 20644 11238 20674 11290
rect 20674 11238 20700 11290
rect 20404 11236 20460 11238
rect 20484 11236 20540 11238
rect 20564 11236 20620 11238
rect 20644 11236 20700 11238
rect 7084 10746 7140 10748
rect 7164 10746 7220 10748
rect 7244 10746 7300 10748
rect 7324 10746 7380 10748
rect 7084 10694 7110 10746
rect 7110 10694 7140 10746
rect 7164 10694 7174 10746
rect 7174 10694 7220 10746
rect 7244 10694 7290 10746
rect 7290 10694 7300 10746
rect 7324 10694 7354 10746
rect 7354 10694 7380 10746
rect 7084 10692 7140 10694
rect 7164 10692 7220 10694
rect 7244 10692 7300 10694
rect 7324 10692 7380 10694
rect 12412 10746 12468 10748
rect 12492 10746 12548 10748
rect 12572 10746 12628 10748
rect 12652 10746 12708 10748
rect 12412 10694 12438 10746
rect 12438 10694 12468 10746
rect 12492 10694 12502 10746
rect 12502 10694 12548 10746
rect 12572 10694 12618 10746
rect 12618 10694 12628 10746
rect 12652 10694 12682 10746
rect 12682 10694 12708 10746
rect 12412 10692 12468 10694
rect 12492 10692 12548 10694
rect 12572 10692 12628 10694
rect 12652 10692 12708 10694
rect 17740 10746 17796 10748
rect 17820 10746 17876 10748
rect 17900 10746 17956 10748
rect 17980 10746 18036 10748
rect 17740 10694 17766 10746
rect 17766 10694 17796 10746
rect 17820 10694 17830 10746
rect 17830 10694 17876 10746
rect 17900 10694 17946 10746
rect 17946 10694 17956 10746
rect 17980 10694 18010 10746
rect 18010 10694 18036 10746
rect 17740 10692 17796 10694
rect 17820 10692 17876 10694
rect 17900 10692 17956 10694
rect 17980 10692 18036 10694
rect 4420 10202 4476 10204
rect 4500 10202 4556 10204
rect 4580 10202 4636 10204
rect 4660 10202 4716 10204
rect 4420 10150 4446 10202
rect 4446 10150 4476 10202
rect 4500 10150 4510 10202
rect 4510 10150 4556 10202
rect 4580 10150 4626 10202
rect 4626 10150 4636 10202
rect 4660 10150 4690 10202
rect 4690 10150 4716 10202
rect 4420 10148 4476 10150
rect 4500 10148 4556 10150
rect 4580 10148 4636 10150
rect 4660 10148 4716 10150
rect 9748 10202 9804 10204
rect 9828 10202 9884 10204
rect 9908 10202 9964 10204
rect 9988 10202 10044 10204
rect 9748 10150 9774 10202
rect 9774 10150 9804 10202
rect 9828 10150 9838 10202
rect 9838 10150 9884 10202
rect 9908 10150 9954 10202
rect 9954 10150 9964 10202
rect 9988 10150 10018 10202
rect 10018 10150 10044 10202
rect 9748 10148 9804 10150
rect 9828 10148 9884 10150
rect 9908 10148 9964 10150
rect 9988 10148 10044 10150
rect 15076 10202 15132 10204
rect 15156 10202 15212 10204
rect 15236 10202 15292 10204
rect 15316 10202 15372 10204
rect 15076 10150 15102 10202
rect 15102 10150 15132 10202
rect 15156 10150 15166 10202
rect 15166 10150 15212 10202
rect 15236 10150 15282 10202
rect 15282 10150 15292 10202
rect 15316 10150 15346 10202
rect 15346 10150 15372 10202
rect 15076 10148 15132 10150
rect 15156 10148 15212 10150
rect 15236 10148 15292 10150
rect 15316 10148 15372 10150
rect 20404 10202 20460 10204
rect 20484 10202 20540 10204
rect 20564 10202 20620 10204
rect 20644 10202 20700 10204
rect 20404 10150 20430 10202
rect 20430 10150 20460 10202
rect 20484 10150 20494 10202
rect 20494 10150 20540 10202
rect 20564 10150 20610 10202
rect 20610 10150 20620 10202
rect 20644 10150 20674 10202
rect 20674 10150 20700 10202
rect 20404 10148 20460 10150
rect 20484 10148 20540 10150
rect 20564 10148 20620 10150
rect 20644 10148 20700 10150
rect 7084 9658 7140 9660
rect 7164 9658 7220 9660
rect 7244 9658 7300 9660
rect 7324 9658 7380 9660
rect 7084 9606 7110 9658
rect 7110 9606 7140 9658
rect 7164 9606 7174 9658
rect 7174 9606 7220 9658
rect 7244 9606 7290 9658
rect 7290 9606 7300 9658
rect 7324 9606 7354 9658
rect 7354 9606 7380 9658
rect 7084 9604 7140 9606
rect 7164 9604 7220 9606
rect 7244 9604 7300 9606
rect 7324 9604 7380 9606
rect 12412 9658 12468 9660
rect 12492 9658 12548 9660
rect 12572 9658 12628 9660
rect 12652 9658 12708 9660
rect 12412 9606 12438 9658
rect 12438 9606 12468 9658
rect 12492 9606 12502 9658
rect 12502 9606 12548 9658
rect 12572 9606 12618 9658
rect 12618 9606 12628 9658
rect 12652 9606 12682 9658
rect 12682 9606 12708 9658
rect 12412 9604 12468 9606
rect 12492 9604 12548 9606
rect 12572 9604 12628 9606
rect 12652 9604 12708 9606
rect 17740 9658 17796 9660
rect 17820 9658 17876 9660
rect 17900 9658 17956 9660
rect 17980 9658 18036 9660
rect 17740 9606 17766 9658
rect 17766 9606 17796 9658
rect 17820 9606 17830 9658
rect 17830 9606 17876 9658
rect 17900 9606 17946 9658
rect 17946 9606 17956 9658
rect 17980 9606 18010 9658
rect 18010 9606 18036 9658
rect 17740 9604 17796 9606
rect 17820 9604 17876 9606
rect 17900 9604 17956 9606
rect 17980 9604 18036 9606
rect 4420 9114 4476 9116
rect 4500 9114 4556 9116
rect 4580 9114 4636 9116
rect 4660 9114 4716 9116
rect 4420 9062 4446 9114
rect 4446 9062 4476 9114
rect 4500 9062 4510 9114
rect 4510 9062 4556 9114
rect 4580 9062 4626 9114
rect 4626 9062 4636 9114
rect 4660 9062 4690 9114
rect 4690 9062 4716 9114
rect 4420 9060 4476 9062
rect 4500 9060 4556 9062
rect 4580 9060 4636 9062
rect 4660 9060 4716 9062
rect 9748 9114 9804 9116
rect 9828 9114 9884 9116
rect 9908 9114 9964 9116
rect 9988 9114 10044 9116
rect 9748 9062 9774 9114
rect 9774 9062 9804 9114
rect 9828 9062 9838 9114
rect 9838 9062 9884 9114
rect 9908 9062 9954 9114
rect 9954 9062 9964 9114
rect 9988 9062 10018 9114
rect 10018 9062 10044 9114
rect 9748 9060 9804 9062
rect 9828 9060 9884 9062
rect 9908 9060 9964 9062
rect 9988 9060 10044 9062
rect 15076 9114 15132 9116
rect 15156 9114 15212 9116
rect 15236 9114 15292 9116
rect 15316 9114 15372 9116
rect 15076 9062 15102 9114
rect 15102 9062 15132 9114
rect 15156 9062 15166 9114
rect 15166 9062 15212 9114
rect 15236 9062 15282 9114
rect 15282 9062 15292 9114
rect 15316 9062 15346 9114
rect 15346 9062 15372 9114
rect 15076 9060 15132 9062
rect 15156 9060 15212 9062
rect 15236 9060 15292 9062
rect 15316 9060 15372 9062
rect 20404 9114 20460 9116
rect 20484 9114 20540 9116
rect 20564 9114 20620 9116
rect 20644 9114 20700 9116
rect 20404 9062 20430 9114
rect 20430 9062 20460 9114
rect 20484 9062 20494 9114
rect 20494 9062 20540 9114
rect 20564 9062 20610 9114
rect 20610 9062 20620 9114
rect 20644 9062 20674 9114
rect 20674 9062 20700 9114
rect 20404 9060 20460 9062
rect 20484 9060 20540 9062
rect 20564 9060 20620 9062
rect 20644 9060 20700 9062
rect 2474 8720 2530 8776
rect 7084 8570 7140 8572
rect 7164 8570 7220 8572
rect 7244 8570 7300 8572
rect 7324 8570 7380 8572
rect 7084 8518 7110 8570
rect 7110 8518 7140 8570
rect 7164 8518 7174 8570
rect 7174 8518 7220 8570
rect 7244 8518 7290 8570
rect 7290 8518 7300 8570
rect 7324 8518 7354 8570
rect 7354 8518 7380 8570
rect 7084 8516 7140 8518
rect 7164 8516 7220 8518
rect 7244 8516 7300 8518
rect 7324 8516 7380 8518
rect 12412 8570 12468 8572
rect 12492 8570 12548 8572
rect 12572 8570 12628 8572
rect 12652 8570 12708 8572
rect 12412 8518 12438 8570
rect 12438 8518 12468 8570
rect 12492 8518 12502 8570
rect 12502 8518 12548 8570
rect 12572 8518 12618 8570
rect 12618 8518 12628 8570
rect 12652 8518 12682 8570
rect 12682 8518 12708 8570
rect 12412 8516 12468 8518
rect 12492 8516 12548 8518
rect 12572 8516 12628 8518
rect 12652 8516 12708 8518
rect 17740 8570 17796 8572
rect 17820 8570 17876 8572
rect 17900 8570 17956 8572
rect 17980 8570 18036 8572
rect 17740 8518 17766 8570
rect 17766 8518 17796 8570
rect 17820 8518 17830 8570
rect 17830 8518 17876 8570
rect 17900 8518 17946 8570
rect 17946 8518 17956 8570
rect 17980 8518 18010 8570
rect 18010 8518 18036 8570
rect 17740 8516 17796 8518
rect 17820 8516 17876 8518
rect 17900 8516 17956 8518
rect 17980 8516 18036 8518
rect 4420 8026 4476 8028
rect 4500 8026 4556 8028
rect 4580 8026 4636 8028
rect 4660 8026 4716 8028
rect 4420 7974 4446 8026
rect 4446 7974 4476 8026
rect 4500 7974 4510 8026
rect 4510 7974 4556 8026
rect 4580 7974 4626 8026
rect 4626 7974 4636 8026
rect 4660 7974 4690 8026
rect 4690 7974 4716 8026
rect 4420 7972 4476 7974
rect 4500 7972 4556 7974
rect 4580 7972 4636 7974
rect 4660 7972 4716 7974
rect 9748 8026 9804 8028
rect 9828 8026 9884 8028
rect 9908 8026 9964 8028
rect 9988 8026 10044 8028
rect 9748 7974 9774 8026
rect 9774 7974 9804 8026
rect 9828 7974 9838 8026
rect 9838 7974 9884 8026
rect 9908 7974 9954 8026
rect 9954 7974 9964 8026
rect 9988 7974 10018 8026
rect 10018 7974 10044 8026
rect 9748 7972 9804 7974
rect 9828 7972 9884 7974
rect 9908 7972 9964 7974
rect 9988 7972 10044 7974
rect 15076 8026 15132 8028
rect 15156 8026 15212 8028
rect 15236 8026 15292 8028
rect 15316 8026 15372 8028
rect 15076 7974 15102 8026
rect 15102 7974 15132 8026
rect 15156 7974 15166 8026
rect 15166 7974 15212 8026
rect 15236 7974 15282 8026
rect 15282 7974 15292 8026
rect 15316 7974 15346 8026
rect 15346 7974 15372 8026
rect 15076 7972 15132 7974
rect 15156 7972 15212 7974
rect 15236 7972 15292 7974
rect 15316 7972 15372 7974
rect 20404 8026 20460 8028
rect 20484 8026 20540 8028
rect 20564 8026 20620 8028
rect 20644 8026 20700 8028
rect 20404 7974 20430 8026
rect 20430 7974 20460 8026
rect 20484 7974 20494 8026
rect 20494 7974 20540 8026
rect 20564 7974 20610 8026
rect 20610 7974 20620 8026
rect 20644 7974 20674 8026
rect 20674 7974 20700 8026
rect 20404 7972 20460 7974
rect 20484 7972 20540 7974
rect 20564 7972 20620 7974
rect 20644 7972 20700 7974
rect 7084 7482 7140 7484
rect 7164 7482 7220 7484
rect 7244 7482 7300 7484
rect 7324 7482 7380 7484
rect 7084 7430 7110 7482
rect 7110 7430 7140 7482
rect 7164 7430 7174 7482
rect 7174 7430 7220 7482
rect 7244 7430 7290 7482
rect 7290 7430 7300 7482
rect 7324 7430 7354 7482
rect 7354 7430 7380 7482
rect 7084 7428 7140 7430
rect 7164 7428 7220 7430
rect 7244 7428 7300 7430
rect 7324 7428 7380 7430
rect 12412 7482 12468 7484
rect 12492 7482 12548 7484
rect 12572 7482 12628 7484
rect 12652 7482 12708 7484
rect 12412 7430 12438 7482
rect 12438 7430 12468 7482
rect 12492 7430 12502 7482
rect 12502 7430 12548 7482
rect 12572 7430 12618 7482
rect 12618 7430 12628 7482
rect 12652 7430 12682 7482
rect 12682 7430 12708 7482
rect 12412 7428 12468 7430
rect 12492 7428 12548 7430
rect 12572 7428 12628 7430
rect 12652 7428 12708 7430
rect 17740 7482 17796 7484
rect 17820 7482 17876 7484
rect 17900 7482 17956 7484
rect 17980 7482 18036 7484
rect 17740 7430 17766 7482
rect 17766 7430 17796 7482
rect 17820 7430 17830 7482
rect 17830 7430 17876 7482
rect 17900 7430 17946 7482
rect 17946 7430 17956 7482
rect 17980 7430 18010 7482
rect 18010 7430 18036 7482
rect 17740 7428 17796 7430
rect 17820 7428 17876 7430
rect 17900 7428 17956 7430
rect 17980 7428 18036 7430
rect 4420 6938 4476 6940
rect 4500 6938 4556 6940
rect 4580 6938 4636 6940
rect 4660 6938 4716 6940
rect 4420 6886 4446 6938
rect 4446 6886 4476 6938
rect 4500 6886 4510 6938
rect 4510 6886 4556 6938
rect 4580 6886 4626 6938
rect 4626 6886 4636 6938
rect 4660 6886 4690 6938
rect 4690 6886 4716 6938
rect 4420 6884 4476 6886
rect 4500 6884 4556 6886
rect 4580 6884 4636 6886
rect 4660 6884 4716 6886
rect 9748 6938 9804 6940
rect 9828 6938 9884 6940
rect 9908 6938 9964 6940
rect 9988 6938 10044 6940
rect 9748 6886 9774 6938
rect 9774 6886 9804 6938
rect 9828 6886 9838 6938
rect 9838 6886 9884 6938
rect 9908 6886 9954 6938
rect 9954 6886 9964 6938
rect 9988 6886 10018 6938
rect 10018 6886 10044 6938
rect 9748 6884 9804 6886
rect 9828 6884 9884 6886
rect 9908 6884 9964 6886
rect 9988 6884 10044 6886
rect 15076 6938 15132 6940
rect 15156 6938 15212 6940
rect 15236 6938 15292 6940
rect 15316 6938 15372 6940
rect 15076 6886 15102 6938
rect 15102 6886 15132 6938
rect 15156 6886 15166 6938
rect 15166 6886 15212 6938
rect 15236 6886 15282 6938
rect 15282 6886 15292 6938
rect 15316 6886 15346 6938
rect 15346 6886 15372 6938
rect 15076 6884 15132 6886
rect 15156 6884 15212 6886
rect 15236 6884 15292 6886
rect 15316 6884 15372 6886
rect 20404 6938 20460 6940
rect 20484 6938 20540 6940
rect 20564 6938 20620 6940
rect 20644 6938 20700 6940
rect 20404 6886 20430 6938
rect 20430 6886 20460 6938
rect 20484 6886 20494 6938
rect 20494 6886 20540 6938
rect 20564 6886 20610 6938
rect 20610 6886 20620 6938
rect 20644 6886 20674 6938
rect 20674 6886 20700 6938
rect 20404 6884 20460 6886
rect 20484 6884 20540 6886
rect 20564 6884 20620 6886
rect 20644 6884 20700 6886
rect 7084 6394 7140 6396
rect 7164 6394 7220 6396
rect 7244 6394 7300 6396
rect 7324 6394 7380 6396
rect 7084 6342 7110 6394
rect 7110 6342 7140 6394
rect 7164 6342 7174 6394
rect 7174 6342 7220 6394
rect 7244 6342 7290 6394
rect 7290 6342 7300 6394
rect 7324 6342 7354 6394
rect 7354 6342 7380 6394
rect 7084 6340 7140 6342
rect 7164 6340 7220 6342
rect 7244 6340 7300 6342
rect 7324 6340 7380 6342
rect 12412 6394 12468 6396
rect 12492 6394 12548 6396
rect 12572 6394 12628 6396
rect 12652 6394 12708 6396
rect 12412 6342 12438 6394
rect 12438 6342 12468 6394
rect 12492 6342 12502 6394
rect 12502 6342 12548 6394
rect 12572 6342 12618 6394
rect 12618 6342 12628 6394
rect 12652 6342 12682 6394
rect 12682 6342 12708 6394
rect 12412 6340 12468 6342
rect 12492 6340 12548 6342
rect 12572 6340 12628 6342
rect 12652 6340 12708 6342
rect 17740 6394 17796 6396
rect 17820 6394 17876 6396
rect 17900 6394 17956 6396
rect 17980 6394 18036 6396
rect 17740 6342 17766 6394
rect 17766 6342 17796 6394
rect 17820 6342 17830 6394
rect 17830 6342 17876 6394
rect 17900 6342 17946 6394
rect 17946 6342 17956 6394
rect 17980 6342 18010 6394
rect 18010 6342 18036 6394
rect 17740 6340 17796 6342
rect 17820 6340 17876 6342
rect 17900 6340 17956 6342
rect 17980 6340 18036 6342
rect 4420 5850 4476 5852
rect 4500 5850 4556 5852
rect 4580 5850 4636 5852
rect 4660 5850 4716 5852
rect 4420 5798 4446 5850
rect 4446 5798 4476 5850
rect 4500 5798 4510 5850
rect 4510 5798 4556 5850
rect 4580 5798 4626 5850
rect 4626 5798 4636 5850
rect 4660 5798 4690 5850
rect 4690 5798 4716 5850
rect 4420 5796 4476 5798
rect 4500 5796 4556 5798
rect 4580 5796 4636 5798
rect 4660 5796 4716 5798
rect 9748 5850 9804 5852
rect 9828 5850 9884 5852
rect 9908 5850 9964 5852
rect 9988 5850 10044 5852
rect 9748 5798 9774 5850
rect 9774 5798 9804 5850
rect 9828 5798 9838 5850
rect 9838 5798 9884 5850
rect 9908 5798 9954 5850
rect 9954 5798 9964 5850
rect 9988 5798 10018 5850
rect 10018 5798 10044 5850
rect 9748 5796 9804 5798
rect 9828 5796 9884 5798
rect 9908 5796 9964 5798
rect 9988 5796 10044 5798
rect 15076 5850 15132 5852
rect 15156 5850 15212 5852
rect 15236 5850 15292 5852
rect 15316 5850 15372 5852
rect 15076 5798 15102 5850
rect 15102 5798 15132 5850
rect 15156 5798 15166 5850
rect 15166 5798 15212 5850
rect 15236 5798 15282 5850
rect 15282 5798 15292 5850
rect 15316 5798 15346 5850
rect 15346 5798 15372 5850
rect 15076 5796 15132 5798
rect 15156 5796 15212 5798
rect 15236 5796 15292 5798
rect 15316 5796 15372 5798
rect 20404 5850 20460 5852
rect 20484 5850 20540 5852
rect 20564 5850 20620 5852
rect 20644 5850 20700 5852
rect 20404 5798 20430 5850
rect 20430 5798 20460 5850
rect 20484 5798 20494 5850
rect 20494 5798 20540 5850
rect 20564 5798 20610 5850
rect 20610 5798 20620 5850
rect 20644 5798 20674 5850
rect 20674 5798 20700 5850
rect 20404 5796 20460 5798
rect 20484 5796 20540 5798
rect 20564 5796 20620 5798
rect 20644 5796 20700 5798
rect 7084 5306 7140 5308
rect 7164 5306 7220 5308
rect 7244 5306 7300 5308
rect 7324 5306 7380 5308
rect 7084 5254 7110 5306
rect 7110 5254 7140 5306
rect 7164 5254 7174 5306
rect 7174 5254 7220 5306
rect 7244 5254 7290 5306
rect 7290 5254 7300 5306
rect 7324 5254 7354 5306
rect 7354 5254 7380 5306
rect 7084 5252 7140 5254
rect 7164 5252 7220 5254
rect 7244 5252 7300 5254
rect 7324 5252 7380 5254
rect 12412 5306 12468 5308
rect 12492 5306 12548 5308
rect 12572 5306 12628 5308
rect 12652 5306 12708 5308
rect 12412 5254 12438 5306
rect 12438 5254 12468 5306
rect 12492 5254 12502 5306
rect 12502 5254 12548 5306
rect 12572 5254 12618 5306
rect 12618 5254 12628 5306
rect 12652 5254 12682 5306
rect 12682 5254 12708 5306
rect 12412 5252 12468 5254
rect 12492 5252 12548 5254
rect 12572 5252 12628 5254
rect 12652 5252 12708 5254
rect 17740 5306 17796 5308
rect 17820 5306 17876 5308
rect 17900 5306 17956 5308
rect 17980 5306 18036 5308
rect 17740 5254 17766 5306
rect 17766 5254 17796 5306
rect 17820 5254 17830 5306
rect 17830 5254 17876 5306
rect 17900 5254 17946 5306
rect 17946 5254 17956 5306
rect 17980 5254 18010 5306
rect 18010 5254 18036 5306
rect 17740 5252 17796 5254
rect 17820 5252 17876 5254
rect 17900 5252 17956 5254
rect 17980 5252 18036 5254
rect 4420 4762 4476 4764
rect 4500 4762 4556 4764
rect 4580 4762 4636 4764
rect 4660 4762 4716 4764
rect 4420 4710 4446 4762
rect 4446 4710 4476 4762
rect 4500 4710 4510 4762
rect 4510 4710 4556 4762
rect 4580 4710 4626 4762
rect 4626 4710 4636 4762
rect 4660 4710 4690 4762
rect 4690 4710 4716 4762
rect 4420 4708 4476 4710
rect 4500 4708 4556 4710
rect 4580 4708 4636 4710
rect 4660 4708 4716 4710
rect 9748 4762 9804 4764
rect 9828 4762 9884 4764
rect 9908 4762 9964 4764
rect 9988 4762 10044 4764
rect 9748 4710 9774 4762
rect 9774 4710 9804 4762
rect 9828 4710 9838 4762
rect 9838 4710 9884 4762
rect 9908 4710 9954 4762
rect 9954 4710 9964 4762
rect 9988 4710 10018 4762
rect 10018 4710 10044 4762
rect 9748 4708 9804 4710
rect 9828 4708 9884 4710
rect 9908 4708 9964 4710
rect 9988 4708 10044 4710
rect 15076 4762 15132 4764
rect 15156 4762 15212 4764
rect 15236 4762 15292 4764
rect 15316 4762 15372 4764
rect 15076 4710 15102 4762
rect 15102 4710 15132 4762
rect 15156 4710 15166 4762
rect 15166 4710 15212 4762
rect 15236 4710 15282 4762
rect 15282 4710 15292 4762
rect 15316 4710 15346 4762
rect 15346 4710 15372 4762
rect 15076 4708 15132 4710
rect 15156 4708 15212 4710
rect 15236 4708 15292 4710
rect 15316 4708 15372 4710
rect 20404 4762 20460 4764
rect 20484 4762 20540 4764
rect 20564 4762 20620 4764
rect 20644 4762 20700 4764
rect 20404 4710 20430 4762
rect 20430 4710 20460 4762
rect 20484 4710 20494 4762
rect 20494 4710 20540 4762
rect 20564 4710 20610 4762
rect 20610 4710 20620 4762
rect 20644 4710 20674 4762
rect 20674 4710 20700 4762
rect 20404 4708 20460 4710
rect 20484 4708 20540 4710
rect 20564 4708 20620 4710
rect 20644 4708 20700 4710
rect 7084 4218 7140 4220
rect 7164 4218 7220 4220
rect 7244 4218 7300 4220
rect 7324 4218 7380 4220
rect 7084 4166 7110 4218
rect 7110 4166 7140 4218
rect 7164 4166 7174 4218
rect 7174 4166 7220 4218
rect 7244 4166 7290 4218
rect 7290 4166 7300 4218
rect 7324 4166 7354 4218
rect 7354 4166 7380 4218
rect 7084 4164 7140 4166
rect 7164 4164 7220 4166
rect 7244 4164 7300 4166
rect 7324 4164 7380 4166
rect 12412 4218 12468 4220
rect 12492 4218 12548 4220
rect 12572 4218 12628 4220
rect 12652 4218 12708 4220
rect 12412 4166 12438 4218
rect 12438 4166 12468 4218
rect 12492 4166 12502 4218
rect 12502 4166 12548 4218
rect 12572 4166 12618 4218
rect 12618 4166 12628 4218
rect 12652 4166 12682 4218
rect 12682 4166 12708 4218
rect 12412 4164 12468 4166
rect 12492 4164 12548 4166
rect 12572 4164 12628 4166
rect 12652 4164 12708 4166
rect 17740 4218 17796 4220
rect 17820 4218 17876 4220
rect 17900 4218 17956 4220
rect 17980 4218 18036 4220
rect 17740 4166 17766 4218
rect 17766 4166 17796 4218
rect 17820 4166 17830 4218
rect 17830 4166 17876 4218
rect 17900 4166 17946 4218
rect 17946 4166 17956 4218
rect 17980 4166 18010 4218
rect 18010 4166 18036 4218
rect 17740 4164 17796 4166
rect 17820 4164 17876 4166
rect 17900 4164 17956 4166
rect 17980 4164 18036 4166
rect 4420 3674 4476 3676
rect 4500 3674 4556 3676
rect 4580 3674 4636 3676
rect 4660 3674 4716 3676
rect 4420 3622 4446 3674
rect 4446 3622 4476 3674
rect 4500 3622 4510 3674
rect 4510 3622 4556 3674
rect 4580 3622 4626 3674
rect 4626 3622 4636 3674
rect 4660 3622 4690 3674
rect 4690 3622 4716 3674
rect 4420 3620 4476 3622
rect 4500 3620 4556 3622
rect 4580 3620 4636 3622
rect 4660 3620 4716 3622
rect 9748 3674 9804 3676
rect 9828 3674 9884 3676
rect 9908 3674 9964 3676
rect 9988 3674 10044 3676
rect 9748 3622 9774 3674
rect 9774 3622 9804 3674
rect 9828 3622 9838 3674
rect 9838 3622 9884 3674
rect 9908 3622 9954 3674
rect 9954 3622 9964 3674
rect 9988 3622 10018 3674
rect 10018 3622 10044 3674
rect 9748 3620 9804 3622
rect 9828 3620 9884 3622
rect 9908 3620 9964 3622
rect 9988 3620 10044 3622
rect 15076 3674 15132 3676
rect 15156 3674 15212 3676
rect 15236 3674 15292 3676
rect 15316 3674 15372 3676
rect 15076 3622 15102 3674
rect 15102 3622 15132 3674
rect 15156 3622 15166 3674
rect 15166 3622 15212 3674
rect 15236 3622 15282 3674
rect 15282 3622 15292 3674
rect 15316 3622 15346 3674
rect 15346 3622 15372 3674
rect 15076 3620 15132 3622
rect 15156 3620 15212 3622
rect 15236 3620 15292 3622
rect 15316 3620 15372 3622
rect 20404 3674 20460 3676
rect 20484 3674 20540 3676
rect 20564 3674 20620 3676
rect 20644 3674 20700 3676
rect 20404 3622 20430 3674
rect 20430 3622 20460 3674
rect 20484 3622 20494 3674
rect 20494 3622 20540 3674
rect 20564 3622 20610 3674
rect 20610 3622 20620 3674
rect 20644 3622 20674 3674
rect 20674 3622 20700 3674
rect 20404 3620 20460 3622
rect 20484 3620 20540 3622
rect 20564 3620 20620 3622
rect 20644 3620 20700 3622
rect 7084 3130 7140 3132
rect 7164 3130 7220 3132
rect 7244 3130 7300 3132
rect 7324 3130 7380 3132
rect 7084 3078 7110 3130
rect 7110 3078 7140 3130
rect 7164 3078 7174 3130
rect 7174 3078 7220 3130
rect 7244 3078 7290 3130
rect 7290 3078 7300 3130
rect 7324 3078 7354 3130
rect 7354 3078 7380 3130
rect 7084 3076 7140 3078
rect 7164 3076 7220 3078
rect 7244 3076 7300 3078
rect 7324 3076 7380 3078
rect 12412 3130 12468 3132
rect 12492 3130 12548 3132
rect 12572 3130 12628 3132
rect 12652 3130 12708 3132
rect 12412 3078 12438 3130
rect 12438 3078 12468 3130
rect 12492 3078 12502 3130
rect 12502 3078 12548 3130
rect 12572 3078 12618 3130
rect 12618 3078 12628 3130
rect 12652 3078 12682 3130
rect 12682 3078 12708 3130
rect 12412 3076 12468 3078
rect 12492 3076 12548 3078
rect 12572 3076 12628 3078
rect 12652 3076 12708 3078
rect 17740 3130 17796 3132
rect 17820 3130 17876 3132
rect 17900 3130 17956 3132
rect 17980 3130 18036 3132
rect 17740 3078 17766 3130
rect 17766 3078 17796 3130
rect 17820 3078 17830 3130
rect 17830 3078 17876 3130
rect 17900 3078 17946 3130
rect 17946 3078 17956 3130
rect 17980 3078 18010 3130
rect 18010 3078 18036 3130
rect 17740 3076 17796 3078
rect 17820 3076 17876 3078
rect 17900 3076 17956 3078
rect 17980 3076 18036 3078
rect 4420 2586 4476 2588
rect 4500 2586 4556 2588
rect 4580 2586 4636 2588
rect 4660 2586 4716 2588
rect 4420 2534 4446 2586
rect 4446 2534 4476 2586
rect 4500 2534 4510 2586
rect 4510 2534 4556 2586
rect 4580 2534 4626 2586
rect 4626 2534 4636 2586
rect 4660 2534 4690 2586
rect 4690 2534 4716 2586
rect 4420 2532 4476 2534
rect 4500 2532 4556 2534
rect 4580 2532 4636 2534
rect 4660 2532 4716 2534
rect 9748 2586 9804 2588
rect 9828 2586 9884 2588
rect 9908 2586 9964 2588
rect 9988 2586 10044 2588
rect 9748 2534 9774 2586
rect 9774 2534 9804 2586
rect 9828 2534 9838 2586
rect 9838 2534 9884 2586
rect 9908 2534 9954 2586
rect 9954 2534 9964 2586
rect 9988 2534 10018 2586
rect 10018 2534 10044 2586
rect 9748 2532 9804 2534
rect 9828 2532 9884 2534
rect 9908 2532 9964 2534
rect 9988 2532 10044 2534
rect 15076 2586 15132 2588
rect 15156 2586 15212 2588
rect 15236 2586 15292 2588
rect 15316 2586 15372 2588
rect 15076 2534 15102 2586
rect 15102 2534 15132 2586
rect 15156 2534 15166 2586
rect 15166 2534 15212 2586
rect 15236 2534 15282 2586
rect 15282 2534 15292 2586
rect 15316 2534 15346 2586
rect 15346 2534 15372 2586
rect 15076 2532 15132 2534
rect 15156 2532 15212 2534
rect 15236 2532 15292 2534
rect 15316 2532 15372 2534
rect 20404 2586 20460 2588
rect 20484 2586 20540 2588
rect 20564 2586 20620 2588
rect 20644 2586 20700 2588
rect 20404 2534 20430 2586
rect 20430 2534 20460 2586
rect 20484 2534 20494 2586
rect 20494 2534 20540 2586
rect 20564 2534 20610 2586
rect 20610 2534 20620 2586
rect 20644 2534 20674 2586
rect 20674 2534 20700 2586
rect 20404 2532 20460 2534
rect 20484 2532 20540 2534
rect 20564 2532 20620 2534
rect 20644 2532 20700 2534
rect 7084 2042 7140 2044
rect 7164 2042 7220 2044
rect 7244 2042 7300 2044
rect 7324 2042 7380 2044
rect 7084 1990 7110 2042
rect 7110 1990 7140 2042
rect 7164 1990 7174 2042
rect 7174 1990 7220 2042
rect 7244 1990 7290 2042
rect 7290 1990 7300 2042
rect 7324 1990 7354 2042
rect 7354 1990 7380 2042
rect 7084 1988 7140 1990
rect 7164 1988 7220 1990
rect 7244 1988 7300 1990
rect 7324 1988 7380 1990
rect 12412 2042 12468 2044
rect 12492 2042 12548 2044
rect 12572 2042 12628 2044
rect 12652 2042 12708 2044
rect 12412 1990 12438 2042
rect 12438 1990 12468 2042
rect 12492 1990 12502 2042
rect 12502 1990 12548 2042
rect 12572 1990 12618 2042
rect 12618 1990 12628 2042
rect 12652 1990 12682 2042
rect 12682 1990 12708 2042
rect 12412 1988 12468 1990
rect 12492 1988 12548 1990
rect 12572 1988 12628 1990
rect 12652 1988 12708 1990
rect 17740 2042 17796 2044
rect 17820 2042 17876 2044
rect 17900 2042 17956 2044
rect 17980 2042 18036 2044
rect 17740 1990 17766 2042
rect 17766 1990 17796 2042
rect 17820 1990 17830 2042
rect 17830 1990 17876 2042
rect 17900 1990 17946 2042
rect 17946 1990 17956 2042
rect 17980 1990 18010 2042
rect 18010 1990 18036 2042
rect 17740 1988 17796 1990
rect 17820 1988 17876 1990
rect 17900 1988 17956 1990
rect 17980 1988 18036 1990
rect 4420 1498 4476 1500
rect 4500 1498 4556 1500
rect 4580 1498 4636 1500
rect 4660 1498 4716 1500
rect 4420 1446 4446 1498
rect 4446 1446 4476 1498
rect 4500 1446 4510 1498
rect 4510 1446 4556 1498
rect 4580 1446 4626 1498
rect 4626 1446 4636 1498
rect 4660 1446 4690 1498
rect 4690 1446 4716 1498
rect 4420 1444 4476 1446
rect 4500 1444 4556 1446
rect 4580 1444 4636 1446
rect 4660 1444 4716 1446
rect 9748 1498 9804 1500
rect 9828 1498 9884 1500
rect 9908 1498 9964 1500
rect 9988 1498 10044 1500
rect 9748 1446 9774 1498
rect 9774 1446 9804 1498
rect 9828 1446 9838 1498
rect 9838 1446 9884 1498
rect 9908 1446 9954 1498
rect 9954 1446 9964 1498
rect 9988 1446 10018 1498
rect 10018 1446 10044 1498
rect 9748 1444 9804 1446
rect 9828 1444 9884 1446
rect 9908 1444 9964 1446
rect 9988 1444 10044 1446
rect 15076 1498 15132 1500
rect 15156 1498 15212 1500
rect 15236 1498 15292 1500
rect 15316 1498 15372 1500
rect 15076 1446 15102 1498
rect 15102 1446 15132 1498
rect 15156 1446 15166 1498
rect 15166 1446 15212 1498
rect 15236 1446 15282 1498
rect 15282 1446 15292 1498
rect 15316 1446 15346 1498
rect 15346 1446 15372 1498
rect 15076 1444 15132 1446
rect 15156 1444 15212 1446
rect 15236 1444 15292 1446
rect 15316 1444 15372 1446
rect 20404 1498 20460 1500
rect 20484 1498 20540 1500
rect 20564 1498 20620 1500
rect 20644 1498 20700 1500
rect 20404 1446 20430 1498
rect 20430 1446 20460 1498
rect 20484 1446 20494 1498
rect 20494 1446 20540 1498
rect 20564 1446 20610 1498
rect 20610 1446 20620 1498
rect 20644 1446 20674 1498
rect 20674 1446 20700 1498
rect 20404 1444 20460 1446
rect 20484 1444 20540 1446
rect 20564 1444 20620 1446
rect 20644 1444 20700 1446
rect 2290 1104 2346 1160
rect 2934 1140 2936 1160
rect 2936 1140 2988 1160
rect 2988 1140 2990 1160
rect 2934 1104 2990 1140
rect 7084 954 7140 956
rect 7164 954 7220 956
rect 7244 954 7300 956
rect 7324 954 7380 956
rect 7084 902 7110 954
rect 7110 902 7140 954
rect 7164 902 7174 954
rect 7174 902 7220 954
rect 7244 902 7290 954
rect 7290 902 7300 954
rect 7324 902 7354 954
rect 7354 902 7380 954
rect 7084 900 7140 902
rect 7164 900 7220 902
rect 7244 900 7300 902
rect 7324 900 7380 902
rect 12412 954 12468 956
rect 12492 954 12548 956
rect 12572 954 12628 956
rect 12652 954 12708 956
rect 12412 902 12438 954
rect 12438 902 12468 954
rect 12492 902 12502 954
rect 12502 902 12548 954
rect 12572 902 12618 954
rect 12618 902 12628 954
rect 12652 902 12682 954
rect 12682 902 12708 954
rect 12412 900 12468 902
rect 12492 900 12548 902
rect 12572 900 12628 902
rect 12652 900 12708 902
rect 17740 954 17796 956
rect 17820 954 17876 956
rect 17900 954 17956 956
rect 17980 954 18036 956
rect 17740 902 17766 954
rect 17766 902 17796 954
rect 17820 902 17830 954
rect 17830 902 17876 954
rect 17900 902 17946 954
rect 17946 902 17956 954
rect 17980 902 18010 954
rect 18010 902 18036 954
rect 17740 900 17796 902
rect 17820 900 17876 902
rect 17900 900 17956 902
rect 17980 900 18036 902
<< metal3 >>
rect 1917 22378 1983 22381
rect 830 22376 1983 22378
rect 830 22320 1922 22376
rect 1978 22320 1983 22376
rect 830 22318 1983 22320
rect 830 22136 890 22318
rect 1917 22315 1983 22318
rect 4408 22176 4728 22177
rect 800 22016 920 22136
rect 4408 22112 4416 22176
rect 4480 22112 4496 22176
rect 4560 22112 4576 22176
rect 4640 22112 4656 22176
rect 4720 22112 4728 22176
rect 4408 22111 4728 22112
rect 9736 22176 10056 22177
rect 9736 22112 9744 22176
rect 9808 22112 9824 22176
rect 9888 22112 9904 22176
rect 9968 22112 9984 22176
rect 10048 22112 10056 22176
rect 9736 22111 10056 22112
rect 15064 22176 15384 22177
rect 15064 22112 15072 22176
rect 15136 22112 15152 22176
rect 15216 22112 15232 22176
rect 15296 22112 15312 22176
rect 15376 22112 15384 22176
rect 15064 22111 15384 22112
rect 20392 22176 20712 22177
rect 20392 22112 20400 22176
rect 20464 22112 20480 22176
rect 20544 22112 20560 22176
rect 20624 22112 20640 22176
rect 20704 22112 20712 22176
rect 20392 22111 20712 22112
rect 2469 21834 2535 21837
rect 830 21832 2535 21834
rect 830 21776 2474 21832
rect 2530 21776 2535 21832
rect 830 21774 2535 21776
rect 830 21592 890 21774
rect 2469 21771 2535 21774
rect 7072 21632 7392 21633
rect 800 21472 920 21592
rect 7072 21568 7080 21632
rect 7144 21568 7160 21632
rect 7224 21568 7240 21632
rect 7304 21568 7320 21632
rect 7384 21568 7392 21632
rect 7072 21567 7392 21568
rect 12400 21632 12720 21633
rect 12400 21568 12408 21632
rect 12472 21568 12488 21632
rect 12552 21568 12568 21632
rect 12632 21568 12648 21632
rect 12712 21568 12720 21632
rect 12400 21567 12720 21568
rect 17728 21632 18048 21633
rect 17728 21568 17736 21632
rect 17800 21568 17816 21632
rect 17880 21568 17896 21632
rect 17960 21568 17976 21632
rect 18040 21568 18048 21632
rect 17728 21567 18048 21568
rect 2469 21290 2535 21293
rect 830 21288 2535 21290
rect 830 21232 2474 21288
rect 2530 21232 2535 21288
rect 830 21230 2535 21232
rect 830 21048 890 21230
rect 2469 21227 2535 21230
rect 4408 21088 4728 21089
rect 800 20928 920 21048
rect 4408 21024 4416 21088
rect 4480 21024 4496 21088
rect 4560 21024 4576 21088
rect 4640 21024 4656 21088
rect 4720 21024 4728 21088
rect 4408 21023 4728 21024
rect 9736 21088 10056 21089
rect 9736 21024 9744 21088
rect 9808 21024 9824 21088
rect 9888 21024 9904 21088
rect 9968 21024 9984 21088
rect 10048 21024 10056 21088
rect 9736 21023 10056 21024
rect 15064 21088 15384 21089
rect 15064 21024 15072 21088
rect 15136 21024 15152 21088
rect 15216 21024 15232 21088
rect 15296 21024 15312 21088
rect 15376 21024 15384 21088
rect 15064 21023 15384 21024
rect 20392 21088 20712 21089
rect 20392 21024 20400 21088
rect 20464 21024 20480 21088
rect 20544 21024 20560 21088
rect 20624 21024 20640 21088
rect 20704 21024 20712 21088
rect 20392 21023 20712 21024
rect 7072 20544 7392 20545
rect 7072 20480 7080 20544
rect 7144 20480 7160 20544
rect 7224 20480 7240 20544
rect 7304 20480 7320 20544
rect 7384 20480 7392 20544
rect 7072 20479 7392 20480
rect 12400 20544 12720 20545
rect 12400 20480 12408 20544
rect 12472 20480 12488 20544
rect 12552 20480 12568 20544
rect 12632 20480 12648 20544
rect 12712 20480 12720 20544
rect 12400 20479 12720 20480
rect 17728 20544 18048 20545
rect 17728 20480 17736 20544
rect 17800 20480 17816 20544
rect 17880 20480 17896 20544
rect 17960 20480 17976 20544
rect 18040 20480 18048 20544
rect 17728 20479 18048 20480
rect 2469 20202 2535 20205
rect 830 20200 2535 20202
rect 830 20144 2474 20200
rect 2530 20144 2535 20200
rect 830 20142 2535 20144
rect 830 19960 890 20142
rect 2469 20139 2535 20142
rect 4408 20000 4728 20001
rect 800 19840 920 19960
rect 4408 19936 4416 20000
rect 4480 19936 4496 20000
rect 4560 19936 4576 20000
rect 4640 19936 4656 20000
rect 4720 19936 4728 20000
rect 4408 19935 4728 19936
rect 9736 20000 10056 20001
rect 9736 19936 9744 20000
rect 9808 19936 9824 20000
rect 9888 19936 9904 20000
rect 9968 19936 9984 20000
rect 10048 19936 10056 20000
rect 9736 19935 10056 19936
rect 15064 20000 15384 20001
rect 15064 19936 15072 20000
rect 15136 19936 15152 20000
rect 15216 19936 15232 20000
rect 15296 19936 15312 20000
rect 15376 19936 15384 20000
rect 15064 19935 15384 19936
rect 20392 20000 20712 20001
rect 20392 19936 20400 20000
rect 20464 19936 20480 20000
rect 20544 19936 20560 20000
rect 20624 19936 20640 20000
rect 20704 19936 20712 20000
rect 20392 19935 20712 19936
rect 7072 19456 7392 19457
rect 7072 19392 7080 19456
rect 7144 19392 7160 19456
rect 7224 19392 7240 19456
rect 7304 19392 7320 19456
rect 7384 19392 7392 19456
rect 7072 19391 7392 19392
rect 12400 19456 12720 19457
rect 12400 19392 12408 19456
rect 12472 19392 12488 19456
rect 12552 19392 12568 19456
rect 12632 19392 12648 19456
rect 12712 19392 12720 19456
rect 12400 19391 12720 19392
rect 17728 19456 18048 19457
rect 17728 19392 17736 19456
rect 17800 19392 17816 19456
rect 17880 19392 17896 19456
rect 17960 19392 17976 19456
rect 18040 19392 18048 19456
rect 17728 19391 18048 19392
rect 2469 19114 2535 19117
rect 830 19112 2535 19114
rect 830 19056 2474 19112
rect 2530 19056 2535 19112
rect 830 19054 2535 19056
rect 830 18872 890 19054
rect 2469 19051 2535 19054
rect 4408 18912 4728 18913
rect 800 18752 920 18872
rect 4408 18848 4416 18912
rect 4480 18848 4496 18912
rect 4560 18848 4576 18912
rect 4640 18848 4656 18912
rect 4720 18848 4728 18912
rect 4408 18847 4728 18848
rect 9736 18912 10056 18913
rect 9736 18848 9744 18912
rect 9808 18848 9824 18912
rect 9888 18848 9904 18912
rect 9968 18848 9984 18912
rect 10048 18848 10056 18912
rect 9736 18847 10056 18848
rect 15064 18912 15384 18913
rect 15064 18848 15072 18912
rect 15136 18848 15152 18912
rect 15216 18848 15232 18912
rect 15296 18848 15312 18912
rect 15376 18848 15384 18912
rect 15064 18847 15384 18848
rect 20392 18912 20712 18913
rect 20392 18848 20400 18912
rect 20464 18848 20480 18912
rect 20544 18848 20560 18912
rect 20624 18848 20640 18912
rect 20704 18848 20712 18912
rect 20392 18847 20712 18848
rect 7072 18368 7392 18369
rect 7072 18304 7080 18368
rect 7144 18304 7160 18368
rect 7224 18304 7240 18368
rect 7304 18304 7320 18368
rect 7384 18304 7392 18368
rect 7072 18303 7392 18304
rect 12400 18368 12720 18369
rect 12400 18304 12408 18368
rect 12472 18304 12488 18368
rect 12552 18304 12568 18368
rect 12632 18304 12648 18368
rect 12712 18304 12720 18368
rect 12400 18303 12720 18304
rect 17728 18368 18048 18369
rect 17728 18304 17736 18368
rect 17800 18304 17816 18368
rect 17880 18304 17896 18368
rect 17960 18304 17976 18368
rect 18040 18304 18048 18368
rect 17728 18303 18048 18304
rect 2469 18026 2535 18029
rect 830 18024 2535 18026
rect 830 17968 2474 18024
rect 2530 17968 2535 18024
rect 830 17966 2535 17968
rect 830 17784 890 17966
rect 2469 17963 2535 17966
rect 4408 17824 4728 17825
rect 800 17664 920 17784
rect 4408 17760 4416 17824
rect 4480 17760 4496 17824
rect 4560 17760 4576 17824
rect 4640 17760 4656 17824
rect 4720 17760 4728 17824
rect 4408 17759 4728 17760
rect 9736 17824 10056 17825
rect 9736 17760 9744 17824
rect 9808 17760 9824 17824
rect 9888 17760 9904 17824
rect 9968 17760 9984 17824
rect 10048 17760 10056 17824
rect 9736 17759 10056 17760
rect 15064 17824 15384 17825
rect 15064 17760 15072 17824
rect 15136 17760 15152 17824
rect 15216 17760 15232 17824
rect 15296 17760 15312 17824
rect 15376 17760 15384 17824
rect 15064 17759 15384 17760
rect 20392 17824 20712 17825
rect 20392 17760 20400 17824
rect 20464 17760 20480 17824
rect 20544 17760 20560 17824
rect 20624 17760 20640 17824
rect 20704 17760 20712 17824
rect 20392 17759 20712 17760
rect 7072 17280 7392 17281
rect 7072 17216 7080 17280
rect 7144 17216 7160 17280
rect 7224 17216 7240 17280
rect 7304 17216 7320 17280
rect 7384 17216 7392 17280
rect 7072 17215 7392 17216
rect 12400 17280 12720 17281
rect 12400 17216 12408 17280
rect 12472 17216 12488 17280
rect 12552 17216 12568 17280
rect 12632 17216 12648 17280
rect 12712 17216 12720 17280
rect 12400 17215 12720 17216
rect 17728 17280 18048 17281
rect 17728 17216 17736 17280
rect 17800 17216 17816 17280
rect 17880 17216 17896 17280
rect 17960 17216 17976 17280
rect 18040 17216 18048 17280
rect 17728 17215 18048 17216
rect 4408 16736 4728 16737
rect 800 16576 920 16696
rect 4408 16672 4416 16736
rect 4480 16672 4496 16736
rect 4560 16672 4576 16736
rect 4640 16672 4656 16736
rect 4720 16672 4728 16736
rect 4408 16671 4728 16672
rect 9736 16736 10056 16737
rect 9736 16672 9744 16736
rect 9808 16672 9824 16736
rect 9888 16672 9904 16736
rect 9968 16672 9984 16736
rect 10048 16672 10056 16736
rect 9736 16671 10056 16672
rect 15064 16736 15384 16737
rect 15064 16672 15072 16736
rect 15136 16672 15152 16736
rect 15216 16672 15232 16736
rect 15296 16672 15312 16736
rect 15376 16672 15384 16736
rect 15064 16671 15384 16672
rect 20392 16736 20712 16737
rect 20392 16672 20400 16736
rect 20464 16672 20480 16736
rect 20544 16672 20560 16736
rect 20624 16672 20640 16736
rect 20704 16672 20712 16736
rect 20392 16671 20712 16672
rect 830 16394 890 16576
rect 2469 16394 2535 16397
rect 830 16392 2535 16394
rect 830 16336 2474 16392
rect 2530 16336 2535 16392
rect 830 16334 2535 16336
rect 2469 16331 2535 16334
rect 7072 16192 7392 16193
rect 7072 16128 7080 16192
rect 7144 16128 7160 16192
rect 7224 16128 7240 16192
rect 7304 16128 7320 16192
rect 7384 16128 7392 16192
rect 7072 16127 7392 16128
rect 12400 16192 12720 16193
rect 12400 16128 12408 16192
rect 12472 16128 12488 16192
rect 12552 16128 12568 16192
rect 12632 16128 12648 16192
rect 12712 16128 12720 16192
rect 12400 16127 12720 16128
rect 17728 16192 18048 16193
rect 17728 16128 17736 16192
rect 17800 16128 17816 16192
rect 17880 16128 17896 16192
rect 17960 16128 17976 16192
rect 18040 16128 18048 16192
rect 17728 16127 18048 16128
rect 2469 15850 2535 15853
rect 830 15848 2535 15850
rect 830 15792 2474 15848
rect 2530 15792 2535 15848
rect 830 15790 2535 15792
rect 830 15608 890 15790
rect 2469 15787 2535 15790
rect 4408 15648 4728 15649
rect 800 15488 920 15608
rect 4408 15584 4416 15648
rect 4480 15584 4496 15648
rect 4560 15584 4576 15648
rect 4640 15584 4656 15648
rect 4720 15584 4728 15648
rect 4408 15583 4728 15584
rect 9736 15648 10056 15649
rect 9736 15584 9744 15648
rect 9808 15584 9824 15648
rect 9888 15584 9904 15648
rect 9968 15584 9984 15648
rect 10048 15584 10056 15648
rect 9736 15583 10056 15584
rect 15064 15648 15384 15649
rect 15064 15584 15072 15648
rect 15136 15584 15152 15648
rect 15216 15584 15232 15648
rect 15296 15584 15312 15648
rect 15376 15584 15384 15648
rect 15064 15583 15384 15584
rect 20392 15648 20712 15649
rect 20392 15584 20400 15648
rect 20464 15584 20480 15648
rect 20544 15584 20560 15648
rect 20624 15584 20640 15648
rect 20704 15584 20712 15648
rect 20392 15583 20712 15584
rect 7072 15104 7392 15105
rect 7072 15040 7080 15104
rect 7144 15040 7160 15104
rect 7224 15040 7240 15104
rect 7304 15040 7320 15104
rect 7384 15040 7392 15104
rect 7072 15039 7392 15040
rect 12400 15104 12720 15105
rect 12400 15040 12408 15104
rect 12472 15040 12488 15104
rect 12552 15040 12568 15104
rect 12632 15040 12648 15104
rect 12712 15040 12720 15104
rect 12400 15039 12720 15040
rect 17728 15104 18048 15105
rect 17728 15040 17736 15104
rect 17800 15040 17816 15104
rect 17880 15040 17896 15104
rect 17960 15040 17976 15104
rect 18040 15040 18048 15104
rect 17728 15039 18048 15040
rect 4408 14560 4728 14561
rect 4408 14496 4416 14560
rect 4480 14496 4496 14560
rect 4560 14496 4576 14560
rect 4640 14496 4656 14560
rect 4720 14496 4728 14560
rect 4408 14495 4728 14496
rect 9736 14560 10056 14561
rect 9736 14496 9744 14560
rect 9808 14496 9824 14560
rect 9888 14496 9904 14560
rect 9968 14496 9984 14560
rect 10048 14496 10056 14560
rect 9736 14495 10056 14496
rect 15064 14560 15384 14561
rect 15064 14496 15072 14560
rect 15136 14496 15152 14560
rect 15216 14496 15232 14560
rect 15296 14496 15312 14560
rect 15376 14496 15384 14560
rect 15064 14495 15384 14496
rect 20392 14560 20712 14561
rect 20392 14496 20400 14560
rect 20464 14496 20480 14560
rect 20544 14496 20560 14560
rect 20624 14496 20640 14560
rect 20704 14496 20712 14560
rect 20392 14495 20712 14496
rect 7072 14016 7392 14017
rect 7072 13952 7080 14016
rect 7144 13952 7160 14016
rect 7224 13952 7240 14016
rect 7304 13952 7320 14016
rect 7384 13952 7392 14016
rect 7072 13951 7392 13952
rect 12400 14016 12720 14017
rect 12400 13952 12408 14016
rect 12472 13952 12488 14016
rect 12552 13952 12568 14016
rect 12632 13952 12648 14016
rect 12712 13952 12720 14016
rect 12400 13951 12720 13952
rect 17728 14016 18048 14017
rect 17728 13952 17736 14016
rect 17800 13952 17816 14016
rect 17880 13952 17896 14016
rect 17960 13952 17976 14016
rect 18040 13952 18048 14016
rect 17728 13951 18048 13952
rect 2469 13674 2535 13677
rect 830 13672 2535 13674
rect 830 13616 2474 13672
rect 2530 13616 2535 13672
rect 830 13614 2535 13616
rect 830 13432 890 13614
rect 2469 13611 2535 13614
rect 4408 13472 4728 13473
rect 800 13312 920 13432
rect 4408 13408 4416 13472
rect 4480 13408 4496 13472
rect 4560 13408 4576 13472
rect 4640 13408 4656 13472
rect 4720 13408 4728 13472
rect 4408 13407 4728 13408
rect 9736 13472 10056 13473
rect 9736 13408 9744 13472
rect 9808 13408 9824 13472
rect 9888 13408 9904 13472
rect 9968 13408 9984 13472
rect 10048 13408 10056 13472
rect 9736 13407 10056 13408
rect 15064 13472 15384 13473
rect 15064 13408 15072 13472
rect 15136 13408 15152 13472
rect 15216 13408 15232 13472
rect 15296 13408 15312 13472
rect 15376 13408 15384 13472
rect 15064 13407 15384 13408
rect 20392 13472 20712 13473
rect 20392 13408 20400 13472
rect 20464 13408 20480 13472
rect 20544 13408 20560 13472
rect 20624 13408 20640 13472
rect 20704 13408 20712 13472
rect 20392 13407 20712 13408
rect 7072 12928 7392 12929
rect 7072 12864 7080 12928
rect 7144 12864 7160 12928
rect 7224 12864 7240 12928
rect 7304 12864 7320 12928
rect 7384 12864 7392 12928
rect 7072 12863 7392 12864
rect 12400 12928 12720 12929
rect 12400 12864 12408 12928
rect 12472 12864 12488 12928
rect 12552 12864 12568 12928
rect 12632 12864 12648 12928
rect 12712 12864 12720 12928
rect 12400 12863 12720 12864
rect 17728 12928 18048 12929
rect 17728 12864 17736 12928
rect 17800 12864 17816 12928
rect 17880 12864 17896 12928
rect 17960 12864 17976 12928
rect 18040 12864 18048 12928
rect 17728 12863 18048 12864
rect 4408 12384 4728 12385
rect 4408 12320 4416 12384
rect 4480 12320 4496 12384
rect 4560 12320 4576 12384
rect 4640 12320 4656 12384
rect 4720 12320 4728 12384
rect 4408 12319 4728 12320
rect 9736 12384 10056 12385
rect 9736 12320 9744 12384
rect 9808 12320 9824 12384
rect 9888 12320 9904 12384
rect 9968 12320 9984 12384
rect 10048 12320 10056 12384
rect 9736 12319 10056 12320
rect 15064 12384 15384 12385
rect 15064 12320 15072 12384
rect 15136 12320 15152 12384
rect 15216 12320 15232 12384
rect 15296 12320 15312 12384
rect 15376 12320 15384 12384
rect 15064 12319 15384 12320
rect 20392 12384 20712 12385
rect 20392 12320 20400 12384
rect 20464 12320 20480 12384
rect 20544 12320 20560 12384
rect 20624 12320 20640 12384
rect 20704 12320 20712 12384
rect 20392 12319 20712 12320
rect 7072 11840 7392 11841
rect 7072 11776 7080 11840
rect 7144 11776 7160 11840
rect 7224 11776 7240 11840
rect 7304 11776 7320 11840
rect 7384 11776 7392 11840
rect 7072 11775 7392 11776
rect 12400 11840 12720 11841
rect 12400 11776 12408 11840
rect 12472 11776 12488 11840
rect 12552 11776 12568 11840
rect 12632 11776 12648 11840
rect 12712 11776 12720 11840
rect 12400 11775 12720 11776
rect 17728 11840 18048 11841
rect 17728 11776 17736 11840
rect 17800 11776 17816 11840
rect 17880 11776 17896 11840
rect 17960 11776 17976 11840
rect 18040 11776 18048 11840
rect 17728 11775 18048 11776
rect 4408 11296 4728 11297
rect 4408 11232 4416 11296
rect 4480 11232 4496 11296
rect 4560 11232 4576 11296
rect 4640 11232 4656 11296
rect 4720 11232 4728 11296
rect 4408 11231 4728 11232
rect 9736 11296 10056 11297
rect 9736 11232 9744 11296
rect 9808 11232 9824 11296
rect 9888 11232 9904 11296
rect 9968 11232 9984 11296
rect 10048 11232 10056 11296
rect 9736 11231 10056 11232
rect 15064 11296 15384 11297
rect 15064 11232 15072 11296
rect 15136 11232 15152 11296
rect 15216 11232 15232 11296
rect 15296 11232 15312 11296
rect 15376 11232 15384 11296
rect 15064 11231 15384 11232
rect 20392 11296 20712 11297
rect 20392 11232 20400 11296
rect 20464 11232 20480 11296
rect 20544 11232 20560 11296
rect 20624 11232 20640 11296
rect 20704 11232 20712 11296
rect 20392 11231 20712 11232
rect 7072 10752 7392 10753
rect 7072 10688 7080 10752
rect 7144 10688 7160 10752
rect 7224 10688 7240 10752
rect 7304 10688 7320 10752
rect 7384 10688 7392 10752
rect 7072 10687 7392 10688
rect 12400 10752 12720 10753
rect 12400 10688 12408 10752
rect 12472 10688 12488 10752
rect 12552 10688 12568 10752
rect 12632 10688 12648 10752
rect 12712 10688 12720 10752
rect 12400 10687 12720 10688
rect 17728 10752 18048 10753
rect 17728 10688 17736 10752
rect 17800 10688 17816 10752
rect 17880 10688 17896 10752
rect 17960 10688 17976 10752
rect 18040 10688 18048 10752
rect 17728 10687 18048 10688
rect 4408 10208 4728 10209
rect 4408 10144 4416 10208
rect 4480 10144 4496 10208
rect 4560 10144 4576 10208
rect 4640 10144 4656 10208
rect 4720 10144 4728 10208
rect 4408 10143 4728 10144
rect 9736 10208 10056 10209
rect 9736 10144 9744 10208
rect 9808 10144 9824 10208
rect 9888 10144 9904 10208
rect 9968 10144 9984 10208
rect 10048 10144 10056 10208
rect 9736 10143 10056 10144
rect 15064 10208 15384 10209
rect 15064 10144 15072 10208
rect 15136 10144 15152 10208
rect 15216 10144 15232 10208
rect 15296 10144 15312 10208
rect 15376 10144 15384 10208
rect 15064 10143 15384 10144
rect 20392 10208 20712 10209
rect 20392 10144 20400 10208
rect 20464 10144 20480 10208
rect 20544 10144 20560 10208
rect 20624 10144 20640 10208
rect 20704 10144 20712 10208
rect 20392 10143 20712 10144
rect 7072 9664 7392 9665
rect 7072 9600 7080 9664
rect 7144 9600 7160 9664
rect 7224 9600 7240 9664
rect 7304 9600 7320 9664
rect 7384 9600 7392 9664
rect 7072 9599 7392 9600
rect 12400 9664 12720 9665
rect 12400 9600 12408 9664
rect 12472 9600 12488 9664
rect 12552 9600 12568 9664
rect 12632 9600 12648 9664
rect 12712 9600 12720 9664
rect 12400 9599 12720 9600
rect 17728 9664 18048 9665
rect 17728 9600 17736 9664
rect 17800 9600 17816 9664
rect 17880 9600 17896 9664
rect 17960 9600 17976 9664
rect 18040 9600 18048 9664
rect 17728 9599 18048 9600
rect 4408 9120 4728 9121
rect 800 8960 920 9080
rect 4408 9056 4416 9120
rect 4480 9056 4496 9120
rect 4560 9056 4576 9120
rect 4640 9056 4656 9120
rect 4720 9056 4728 9120
rect 4408 9055 4728 9056
rect 9736 9120 10056 9121
rect 9736 9056 9744 9120
rect 9808 9056 9824 9120
rect 9888 9056 9904 9120
rect 9968 9056 9984 9120
rect 10048 9056 10056 9120
rect 9736 9055 10056 9056
rect 15064 9120 15384 9121
rect 15064 9056 15072 9120
rect 15136 9056 15152 9120
rect 15216 9056 15232 9120
rect 15296 9056 15312 9120
rect 15376 9056 15384 9120
rect 15064 9055 15384 9056
rect 20392 9120 20712 9121
rect 20392 9056 20400 9120
rect 20464 9056 20480 9120
rect 20544 9056 20560 9120
rect 20624 9056 20640 9120
rect 20704 9056 20712 9120
rect 20392 9055 20712 9056
rect 830 8778 890 8960
rect 2469 8778 2535 8781
rect 830 8776 2535 8778
rect 830 8720 2474 8776
rect 2530 8720 2535 8776
rect 830 8718 2535 8720
rect 2469 8715 2535 8718
rect 7072 8576 7392 8577
rect 7072 8512 7080 8576
rect 7144 8512 7160 8576
rect 7224 8512 7240 8576
rect 7304 8512 7320 8576
rect 7384 8512 7392 8576
rect 7072 8511 7392 8512
rect 12400 8576 12720 8577
rect 12400 8512 12408 8576
rect 12472 8512 12488 8576
rect 12552 8512 12568 8576
rect 12632 8512 12648 8576
rect 12712 8512 12720 8576
rect 12400 8511 12720 8512
rect 17728 8576 18048 8577
rect 17728 8512 17736 8576
rect 17800 8512 17816 8576
rect 17880 8512 17896 8576
rect 17960 8512 17976 8576
rect 18040 8512 18048 8576
rect 17728 8511 18048 8512
rect 4408 8032 4728 8033
rect 4408 7968 4416 8032
rect 4480 7968 4496 8032
rect 4560 7968 4576 8032
rect 4640 7968 4656 8032
rect 4720 7968 4728 8032
rect 4408 7967 4728 7968
rect 9736 8032 10056 8033
rect 9736 7968 9744 8032
rect 9808 7968 9824 8032
rect 9888 7968 9904 8032
rect 9968 7968 9984 8032
rect 10048 7968 10056 8032
rect 9736 7967 10056 7968
rect 15064 8032 15384 8033
rect 15064 7968 15072 8032
rect 15136 7968 15152 8032
rect 15216 7968 15232 8032
rect 15296 7968 15312 8032
rect 15376 7968 15384 8032
rect 15064 7967 15384 7968
rect 20392 8032 20712 8033
rect 20392 7968 20400 8032
rect 20464 7968 20480 8032
rect 20544 7968 20560 8032
rect 20624 7968 20640 8032
rect 20704 7968 20712 8032
rect 20392 7967 20712 7968
rect 7072 7488 7392 7489
rect 7072 7424 7080 7488
rect 7144 7424 7160 7488
rect 7224 7424 7240 7488
rect 7304 7424 7320 7488
rect 7384 7424 7392 7488
rect 7072 7423 7392 7424
rect 12400 7488 12720 7489
rect 12400 7424 12408 7488
rect 12472 7424 12488 7488
rect 12552 7424 12568 7488
rect 12632 7424 12648 7488
rect 12712 7424 12720 7488
rect 12400 7423 12720 7424
rect 17728 7488 18048 7489
rect 17728 7424 17736 7488
rect 17800 7424 17816 7488
rect 17880 7424 17896 7488
rect 17960 7424 17976 7488
rect 18040 7424 18048 7488
rect 17728 7423 18048 7424
rect 4408 6944 4728 6945
rect 4408 6880 4416 6944
rect 4480 6880 4496 6944
rect 4560 6880 4576 6944
rect 4640 6880 4656 6944
rect 4720 6880 4728 6944
rect 4408 6879 4728 6880
rect 9736 6944 10056 6945
rect 9736 6880 9744 6944
rect 9808 6880 9824 6944
rect 9888 6880 9904 6944
rect 9968 6880 9984 6944
rect 10048 6880 10056 6944
rect 9736 6879 10056 6880
rect 15064 6944 15384 6945
rect 15064 6880 15072 6944
rect 15136 6880 15152 6944
rect 15216 6880 15232 6944
rect 15296 6880 15312 6944
rect 15376 6880 15384 6944
rect 15064 6879 15384 6880
rect 20392 6944 20712 6945
rect 20392 6880 20400 6944
rect 20464 6880 20480 6944
rect 20544 6880 20560 6944
rect 20624 6880 20640 6944
rect 20704 6880 20712 6944
rect 20392 6879 20712 6880
rect 7072 6400 7392 6401
rect 7072 6336 7080 6400
rect 7144 6336 7160 6400
rect 7224 6336 7240 6400
rect 7304 6336 7320 6400
rect 7384 6336 7392 6400
rect 7072 6335 7392 6336
rect 12400 6400 12720 6401
rect 12400 6336 12408 6400
rect 12472 6336 12488 6400
rect 12552 6336 12568 6400
rect 12632 6336 12648 6400
rect 12712 6336 12720 6400
rect 12400 6335 12720 6336
rect 17728 6400 18048 6401
rect 17728 6336 17736 6400
rect 17800 6336 17816 6400
rect 17880 6336 17896 6400
rect 17960 6336 17976 6400
rect 18040 6336 18048 6400
rect 17728 6335 18048 6336
rect 4408 5856 4728 5857
rect 4408 5792 4416 5856
rect 4480 5792 4496 5856
rect 4560 5792 4576 5856
rect 4640 5792 4656 5856
rect 4720 5792 4728 5856
rect 4408 5791 4728 5792
rect 9736 5856 10056 5857
rect 9736 5792 9744 5856
rect 9808 5792 9824 5856
rect 9888 5792 9904 5856
rect 9968 5792 9984 5856
rect 10048 5792 10056 5856
rect 9736 5791 10056 5792
rect 15064 5856 15384 5857
rect 15064 5792 15072 5856
rect 15136 5792 15152 5856
rect 15216 5792 15232 5856
rect 15296 5792 15312 5856
rect 15376 5792 15384 5856
rect 15064 5791 15384 5792
rect 20392 5856 20712 5857
rect 20392 5792 20400 5856
rect 20464 5792 20480 5856
rect 20544 5792 20560 5856
rect 20624 5792 20640 5856
rect 20704 5792 20712 5856
rect 20392 5791 20712 5792
rect 7072 5312 7392 5313
rect 7072 5248 7080 5312
rect 7144 5248 7160 5312
rect 7224 5248 7240 5312
rect 7304 5248 7320 5312
rect 7384 5248 7392 5312
rect 7072 5247 7392 5248
rect 12400 5312 12720 5313
rect 12400 5248 12408 5312
rect 12472 5248 12488 5312
rect 12552 5248 12568 5312
rect 12632 5248 12648 5312
rect 12712 5248 12720 5312
rect 12400 5247 12720 5248
rect 17728 5312 18048 5313
rect 17728 5248 17736 5312
rect 17800 5248 17816 5312
rect 17880 5248 17896 5312
rect 17960 5248 17976 5312
rect 18040 5248 18048 5312
rect 17728 5247 18048 5248
rect 4408 4768 4728 4769
rect 4408 4704 4416 4768
rect 4480 4704 4496 4768
rect 4560 4704 4576 4768
rect 4640 4704 4656 4768
rect 4720 4704 4728 4768
rect 4408 4703 4728 4704
rect 9736 4768 10056 4769
rect 9736 4704 9744 4768
rect 9808 4704 9824 4768
rect 9888 4704 9904 4768
rect 9968 4704 9984 4768
rect 10048 4704 10056 4768
rect 9736 4703 10056 4704
rect 15064 4768 15384 4769
rect 15064 4704 15072 4768
rect 15136 4704 15152 4768
rect 15216 4704 15232 4768
rect 15296 4704 15312 4768
rect 15376 4704 15384 4768
rect 15064 4703 15384 4704
rect 20392 4768 20712 4769
rect 20392 4704 20400 4768
rect 20464 4704 20480 4768
rect 20544 4704 20560 4768
rect 20624 4704 20640 4768
rect 20704 4704 20712 4768
rect 20392 4703 20712 4704
rect 7072 4224 7392 4225
rect 7072 4160 7080 4224
rect 7144 4160 7160 4224
rect 7224 4160 7240 4224
rect 7304 4160 7320 4224
rect 7384 4160 7392 4224
rect 7072 4159 7392 4160
rect 12400 4224 12720 4225
rect 12400 4160 12408 4224
rect 12472 4160 12488 4224
rect 12552 4160 12568 4224
rect 12632 4160 12648 4224
rect 12712 4160 12720 4224
rect 12400 4159 12720 4160
rect 17728 4224 18048 4225
rect 17728 4160 17736 4224
rect 17800 4160 17816 4224
rect 17880 4160 17896 4224
rect 17960 4160 17976 4224
rect 18040 4160 18048 4224
rect 17728 4159 18048 4160
rect 4408 3680 4728 3681
rect 4408 3616 4416 3680
rect 4480 3616 4496 3680
rect 4560 3616 4576 3680
rect 4640 3616 4656 3680
rect 4720 3616 4728 3680
rect 4408 3615 4728 3616
rect 9736 3680 10056 3681
rect 9736 3616 9744 3680
rect 9808 3616 9824 3680
rect 9888 3616 9904 3680
rect 9968 3616 9984 3680
rect 10048 3616 10056 3680
rect 9736 3615 10056 3616
rect 15064 3680 15384 3681
rect 15064 3616 15072 3680
rect 15136 3616 15152 3680
rect 15216 3616 15232 3680
rect 15296 3616 15312 3680
rect 15376 3616 15384 3680
rect 15064 3615 15384 3616
rect 20392 3680 20712 3681
rect 20392 3616 20400 3680
rect 20464 3616 20480 3680
rect 20544 3616 20560 3680
rect 20624 3616 20640 3680
rect 20704 3616 20712 3680
rect 20392 3615 20712 3616
rect 7072 3136 7392 3137
rect 7072 3072 7080 3136
rect 7144 3072 7160 3136
rect 7224 3072 7240 3136
rect 7304 3072 7320 3136
rect 7384 3072 7392 3136
rect 7072 3071 7392 3072
rect 12400 3136 12720 3137
rect 12400 3072 12408 3136
rect 12472 3072 12488 3136
rect 12552 3072 12568 3136
rect 12632 3072 12648 3136
rect 12712 3072 12720 3136
rect 12400 3071 12720 3072
rect 17728 3136 18048 3137
rect 17728 3072 17736 3136
rect 17800 3072 17816 3136
rect 17880 3072 17896 3136
rect 17960 3072 17976 3136
rect 18040 3072 18048 3136
rect 17728 3071 18048 3072
rect 4408 2592 4728 2593
rect 4408 2528 4416 2592
rect 4480 2528 4496 2592
rect 4560 2528 4576 2592
rect 4640 2528 4656 2592
rect 4720 2528 4728 2592
rect 4408 2527 4728 2528
rect 9736 2592 10056 2593
rect 9736 2528 9744 2592
rect 9808 2528 9824 2592
rect 9888 2528 9904 2592
rect 9968 2528 9984 2592
rect 10048 2528 10056 2592
rect 9736 2527 10056 2528
rect 15064 2592 15384 2593
rect 15064 2528 15072 2592
rect 15136 2528 15152 2592
rect 15216 2528 15232 2592
rect 15296 2528 15312 2592
rect 15376 2528 15384 2592
rect 15064 2527 15384 2528
rect 20392 2592 20712 2593
rect 20392 2528 20400 2592
rect 20464 2528 20480 2592
rect 20544 2528 20560 2592
rect 20624 2528 20640 2592
rect 20704 2528 20712 2592
rect 20392 2527 20712 2528
rect 7072 2048 7392 2049
rect 7072 1984 7080 2048
rect 7144 1984 7160 2048
rect 7224 1984 7240 2048
rect 7304 1984 7320 2048
rect 7384 1984 7392 2048
rect 7072 1983 7392 1984
rect 12400 2048 12720 2049
rect 12400 1984 12408 2048
rect 12472 1984 12488 2048
rect 12552 1984 12568 2048
rect 12632 1984 12648 2048
rect 12712 1984 12720 2048
rect 12400 1983 12720 1984
rect 17728 2048 18048 2049
rect 17728 1984 17736 2048
rect 17800 1984 17816 2048
rect 17880 1984 17896 2048
rect 17960 1984 17976 2048
rect 18040 1984 18048 2048
rect 17728 1983 18048 1984
rect 4408 1504 4728 1505
rect 4408 1440 4416 1504
rect 4480 1440 4496 1504
rect 4560 1440 4576 1504
rect 4640 1440 4656 1504
rect 4720 1440 4728 1504
rect 4408 1439 4728 1440
rect 9736 1504 10056 1505
rect 9736 1440 9744 1504
rect 9808 1440 9824 1504
rect 9888 1440 9904 1504
rect 9968 1440 9984 1504
rect 10048 1440 10056 1504
rect 9736 1439 10056 1440
rect 15064 1504 15384 1505
rect 15064 1440 15072 1504
rect 15136 1440 15152 1504
rect 15216 1440 15232 1504
rect 15296 1440 15312 1504
rect 15376 1440 15384 1504
rect 15064 1439 15384 1440
rect 20392 1504 20712 1505
rect 20392 1440 20400 1504
rect 20464 1440 20480 1504
rect 20544 1440 20560 1504
rect 20624 1440 20640 1504
rect 20704 1440 20712 1504
rect 20392 1439 20712 1440
rect 2285 1162 2351 1165
rect 2929 1162 2995 1165
rect 830 1160 2995 1162
rect 830 1104 2290 1160
rect 2346 1104 2934 1160
rect 2990 1104 2995 1160
rect 830 1102 2995 1104
rect 830 920 890 1102
rect 2285 1099 2351 1102
rect 2929 1099 2995 1102
rect 7072 960 7392 961
rect 800 800 920 920
rect 7072 896 7080 960
rect 7144 896 7160 960
rect 7224 896 7240 960
rect 7304 896 7320 960
rect 7384 896 7392 960
rect 7072 895 7392 896
rect 12400 960 12720 961
rect 12400 896 12408 960
rect 12472 896 12488 960
rect 12552 896 12568 960
rect 12632 896 12648 960
rect 12712 896 12720 960
rect 12400 895 12720 896
rect 17728 960 18048 961
rect 17728 896 17736 960
rect 17800 896 17816 960
rect 17880 896 17896 960
rect 17960 896 17976 960
rect 18040 896 18048 960
rect 17728 895 18048 896
<< via3 >>
rect 4416 22172 4480 22176
rect 4416 22116 4420 22172
rect 4420 22116 4476 22172
rect 4476 22116 4480 22172
rect 4416 22112 4480 22116
rect 4496 22172 4560 22176
rect 4496 22116 4500 22172
rect 4500 22116 4556 22172
rect 4556 22116 4560 22172
rect 4496 22112 4560 22116
rect 4576 22172 4640 22176
rect 4576 22116 4580 22172
rect 4580 22116 4636 22172
rect 4636 22116 4640 22172
rect 4576 22112 4640 22116
rect 4656 22172 4720 22176
rect 4656 22116 4660 22172
rect 4660 22116 4716 22172
rect 4716 22116 4720 22172
rect 4656 22112 4720 22116
rect 9744 22172 9808 22176
rect 9744 22116 9748 22172
rect 9748 22116 9804 22172
rect 9804 22116 9808 22172
rect 9744 22112 9808 22116
rect 9824 22172 9888 22176
rect 9824 22116 9828 22172
rect 9828 22116 9884 22172
rect 9884 22116 9888 22172
rect 9824 22112 9888 22116
rect 9904 22172 9968 22176
rect 9904 22116 9908 22172
rect 9908 22116 9964 22172
rect 9964 22116 9968 22172
rect 9904 22112 9968 22116
rect 9984 22172 10048 22176
rect 9984 22116 9988 22172
rect 9988 22116 10044 22172
rect 10044 22116 10048 22172
rect 9984 22112 10048 22116
rect 15072 22172 15136 22176
rect 15072 22116 15076 22172
rect 15076 22116 15132 22172
rect 15132 22116 15136 22172
rect 15072 22112 15136 22116
rect 15152 22172 15216 22176
rect 15152 22116 15156 22172
rect 15156 22116 15212 22172
rect 15212 22116 15216 22172
rect 15152 22112 15216 22116
rect 15232 22172 15296 22176
rect 15232 22116 15236 22172
rect 15236 22116 15292 22172
rect 15292 22116 15296 22172
rect 15232 22112 15296 22116
rect 15312 22172 15376 22176
rect 15312 22116 15316 22172
rect 15316 22116 15372 22172
rect 15372 22116 15376 22172
rect 15312 22112 15376 22116
rect 20400 22172 20464 22176
rect 20400 22116 20404 22172
rect 20404 22116 20460 22172
rect 20460 22116 20464 22172
rect 20400 22112 20464 22116
rect 20480 22172 20544 22176
rect 20480 22116 20484 22172
rect 20484 22116 20540 22172
rect 20540 22116 20544 22172
rect 20480 22112 20544 22116
rect 20560 22172 20624 22176
rect 20560 22116 20564 22172
rect 20564 22116 20620 22172
rect 20620 22116 20624 22172
rect 20560 22112 20624 22116
rect 20640 22172 20704 22176
rect 20640 22116 20644 22172
rect 20644 22116 20700 22172
rect 20700 22116 20704 22172
rect 20640 22112 20704 22116
rect 7080 21628 7144 21632
rect 7080 21572 7084 21628
rect 7084 21572 7140 21628
rect 7140 21572 7144 21628
rect 7080 21568 7144 21572
rect 7160 21628 7224 21632
rect 7160 21572 7164 21628
rect 7164 21572 7220 21628
rect 7220 21572 7224 21628
rect 7160 21568 7224 21572
rect 7240 21628 7304 21632
rect 7240 21572 7244 21628
rect 7244 21572 7300 21628
rect 7300 21572 7304 21628
rect 7240 21568 7304 21572
rect 7320 21628 7384 21632
rect 7320 21572 7324 21628
rect 7324 21572 7380 21628
rect 7380 21572 7384 21628
rect 7320 21568 7384 21572
rect 12408 21628 12472 21632
rect 12408 21572 12412 21628
rect 12412 21572 12468 21628
rect 12468 21572 12472 21628
rect 12408 21568 12472 21572
rect 12488 21628 12552 21632
rect 12488 21572 12492 21628
rect 12492 21572 12548 21628
rect 12548 21572 12552 21628
rect 12488 21568 12552 21572
rect 12568 21628 12632 21632
rect 12568 21572 12572 21628
rect 12572 21572 12628 21628
rect 12628 21572 12632 21628
rect 12568 21568 12632 21572
rect 12648 21628 12712 21632
rect 12648 21572 12652 21628
rect 12652 21572 12708 21628
rect 12708 21572 12712 21628
rect 12648 21568 12712 21572
rect 17736 21628 17800 21632
rect 17736 21572 17740 21628
rect 17740 21572 17796 21628
rect 17796 21572 17800 21628
rect 17736 21568 17800 21572
rect 17816 21628 17880 21632
rect 17816 21572 17820 21628
rect 17820 21572 17876 21628
rect 17876 21572 17880 21628
rect 17816 21568 17880 21572
rect 17896 21628 17960 21632
rect 17896 21572 17900 21628
rect 17900 21572 17956 21628
rect 17956 21572 17960 21628
rect 17896 21568 17960 21572
rect 17976 21628 18040 21632
rect 17976 21572 17980 21628
rect 17980 21572 18036 21628
rect 18036 21572 18040 21628
rect 17976 21568 18040 21572
rect 4416 21084 4480 21088
rect 4416 21028 4420 21084
rect 4420 21028 4476 21084
rect 4476 21028 4480 21084
rect 4416 21024 4480 21028
rect 4496 21084 4560 21088
rect 4496 21028 4500 21084
rect 4500 21028 4556 21084
rect 4556 21028 4560 21084
rect 4496 21024 4560 21028
rect 4576 21084 4640 21088
rect 4576 21028 4580 21084
rect 4580 21028 4636 21084
rect 4636 21028 4640 21084
rect 4576 21024 4640 21028
rect 4656 21084 4720 21088
rect 4656 21028 4660 21084
rect 4660 21028 4716 21084
rect 4716 21028 4720 21084
rect 4656 21024 4720 21028
rect 9744 21084 9808 21088
rect 9744 21028 9748 21084
rect 9748 21028 9804 21084
rect 9804 21028 9808 21084
rect 9744 21024 9808 21028
rect 9824 21084 9888 21088
rect 9824 21028 9828 21084
rect 9828 21028 9884 21084
rect 9884 21028 9888 21084
rect 9824 21024 9888 21028
rect 9904 21084 9968 21088
rect 9904 21028 9908 21084
rect 9908 21028 9964 21084
rect 9964 21028 9968 21084
rect 9904 21024 9968 21028
rect 9984 21084 10048 21088
rect 9984 21028 9988 21084
rect 9988 21028 10044 21084
rect 10044 21028 10048 21084
rect 9984 21024 10048 21028
rect 15072 21084 15136 21088
rect 15072 21028 15076 21084
rect 15076 21028 15132 21084
rect 15132 21028 15136 21084
rect 15072 21024 15136 21028
rect 15152 21084 15216 21088
rect 15152 21028 15156 21084
rect 15156 21028 15212 21084
rect 15212 21028 15216 21084
rect 15152 21024 15216 21028
rect 15232 21084 15296 21088
rect 15232 21028 15236 21084
rect 15236 21028 15292 21084
rect 15292 21028 15296 21084
rect 15232 21024 15296 21028
rect 15312 21084 15376 21088
rect 15312 21028 15316 21084
rect 15316 21028 15372 21084
rect 15372 21028 15376 21084
rect 15312 21024 15376 21028
rect 20400 21084 20464 21088
rect 20400 21028 20404 21084
rect 20404 21028 20460 21084
rect 20460 21028 20464 21084
rect 20400 21024 20464 21028
rect 20480 21084 20544 21088
rect 20480 21028 20484 21084
rect 20484 21028 20540 21084
rect 20540 21028 20544 21084
rect 20480 21024 20544 21028
rect 20560 21084 20624 21088
rect 20560 21028 20564 21084
rect 20564 21028 20620 21084
rect 20620 21028 20624 21084
rect 20560 21024 20624 21028
rect 20640 21084 20704 21088
rect 20640 21028 20644 21084
rect 20644 21028 20700 21084
rect 20700 21028 20704 21084
rect 20640 21024 20704 21028
rect 7080 20540 7144 20544
rect 7080 20484 7084 20540
rect 7084 20484 7140 20540
rect 7140 20484 7144 20540
rect 7080 20480 7144 20484
rect 7160 20540 7224 20544
rect 7160 20484 7164 20540
rect 7164 20484 7220 20540
rect 7220 20484 7224 20540
rect 7160 20480 7224 20484
rect 7240 20540 7304 20544
rect 7240 20484 7244 20540
rect 7244 20484 7300 20540
rect 7300 20484 7304 20540
rect 7240 20480 7304 20484
rect 7320 20540 7384 20544
rect 7320 20484 7324 20540
rect 7324 20484 7380 20540
rect 7380 20484 7384 20540
rect 7320 20480 7384 20484
rect 12408 20540 12472 20544
rect 12408 20484 12412 20540
rect 12412 20484 12468 20540
rect 12468 20484 12472 20540
rect 12408 20480 12472 20484
rect 12488 20540 12552 20544
rect 12488 20484 12492 20540
rect 12492 20484 12548 20540
rect 12548 20484 12552 20540
rect 12488 20480 12552 20484
rect 12568 20540 12632 20544
rect 12568 20484 12572 20540
rect 12572 20484 12628 20540
rect 12628 20484 12632 20540
rect 12568 20480 12632 20484
rect 12648 20540 12712 20544
rect 12648 20484 12652 20540
rect 12652 20484 12708 20540
rect 12708 20484 12712 20540
rect 12648 20480 12712 20484
rect 17736 20540 17800 20544
rect 17736 20484 17740 20540
rect 17740 20484 17796 20540
rect 17796 20484 17800 20540
rect 17736 20480 17800 20484
rect 17816 20540 17880 20544
rect 17816 20484 17820 20540
rect 17820 20484 17876 20540
rect 17876 20484 17880 20540
rect 17816 20480 17880 20484
rect 17896 20540 17960 20544
rect 17896 20484 17900 20540
rect 17900 20484 17956 20540
rect 17956 20484 17960 20540
rect 17896 20480 17960 20484
rect 17976 20540 18040 20544
rect 17976 20484 17980 20540
rect 17980 20484 18036 20540
rect 18036 20484 18040 20540
rect 17976 20480 18040 20484
rect 4416 19996 4480 20000
rect 4416 19940 4420 19996
rect 4420 19940 4476 19996
rect 4476 19940 4480 19996
rect 4416 19936 4480 19940
rect 4496 19996 4560 20000
rect 4496 19940 4500 19996
rect 4500 19940 4556 19996
rect 4556 19940 4560 19996
rect 4496 19936 4560 19940
rect 4576 19996 4640 20000
rect 4576 19940 4580 19996
rect 4580 19940 4636 19996
rect 4636 19940 4640 19996
rect 4576 19936 4640 19940
rect 4656 19996 4720 20000
rect 4656 19940 4660 19996
rect 4660 19940 4716 19996
rect 4716 19940 4720 19996
rect 4656 19936 4720 19940
rect 9744 19996 9808 20000
rect 9744 19940 9748 19996
rect 9748 19940 9804 19996
rect 9804 19940 9808 19996
rect 9744 19936 9808 19940
rect 9824 19996 9888 20000
rect 9824 19940 9828 19996
rect 9828 19940 9884 19996
rect 9884 19940 9888 19996
rect 9824 19936 9888 19940
rect 9904 19996 9968 20000
rect 9904 19940 9908 19996
rect 9908 19940 9964 19996
rect 9964 19940 9968 19996
rect 9904 19936 9968 19940
rect 9984 19996 10048 20000
rect 9984 19940 9988 19996
rect 9988 19940 10044 19996
rect 10044 19940 10048 19996
rect 9984 19936 10048 19940
rect 15072 19996 15136 20000
rect 15072 19940 15076 19996
rect 15076 19940 15132 19996
rect 15132 19940 15136 19996
rect 15072 19936 15136 19940
rect 15152 19996 15216 20000
rect 15152 19940 15156 19996
rect 15156 19940 15212 19996
rect 15212 19940 15216 19996
rect 15152 19936 15216 19940
rect 15232 19996 15296 20000
rect 15232 19940 15236 19996
rect 15236 19940 15292 19996
rect 15292 19940 15296 19996
rect 15232 19936 15296 19940
rect 15312 19996 15376 20000
rect 15312 19940 15316 19996
rect 15316 19940 15372 19996
rect 15372 19940 15376 19996
rect 15312 19936 15376 19940
rect 20400 19996 20464 20000
rect 20400 19940 20404 19996
rect 20404 19940 20460 19996
rect 20460 19940 20464 19996
rect 20400 19936 20464 19940
rect 20480 19996 20544 20000
rect 20480 19940 20484 19996
rect 20484 19940 20540 19996
rect 20540 19940 20544 19996
rect 20480 19936 20544 19940
rect 20560 19996 20624 20000
rect 20560 19940 20564 19996
rect 20564 19940 20620 19996
rect 20620 19940 20624 19996
rect 20560 19936 20624 19940
rect 20640 19996 20704 20000
rect 20640 19940 20644 19996
rect 20644 19940 20700 19996
rect 20700 19940 20704 19996
rect 20640 19936 20704 19940
rect 7080 19452 7144 19456
rect 7080 19396 7084 19452
rect 7084 19396 7140 19452
rect 7140 19396 7144 19452
rect 7080 19392 7144 19396
rect 7160 19452 7224 19456
rect 7160 19396 7164 19452
rect 7164 19396 7220 19452
rect 7220 19396 7224 19452
rect 7160 19392 7224 19396
rect 7240 19452 7304 19456
rect 7240 19396 7244 19452
rect 7244 19396 7300 19452
rect 7300 19396 7304 19452
rect 7240 19392 7304 19396
rect 7320 19452 7384 19456
rect 7320 19396 7324 19452
rect 7324 19396 7380 19452
rect 7380 19396 7384 19452
rect 7320 19392 7384 19396
rect 12408 19452 12472 19456
rect 12408 19396 12412 19452
rect 12412 19396 12468 19452
rect 12468 19396 12472 19452
rect 12408 19392 12472 19396
rect 12488 19452 12552 19456
rect 12488 19396 12492 19452
rect 12492 19396 12548 19452
rect 12548 19396 12552 19452
rect 12488 19392 12552 19396
rect 12568 19452 12632 19456
rect 12568 19396 12572 19452
rect 12572 19396 12628 19452
rect 12628 19396 12632 19452
rect 12568 19392 12632 19396
rect 12648 19452 12712 19456
rect 12648 19396 12652 19452
rect 12652 19396 12708 19452
rect 12708 19396 12712 19452
rect 12648 19392 12712 19396
rect 17736 19452 17800 19456
rect 17736 19396 17740 19452
rect 17740 19396 17796 19452
rect 17796 19396 17800 19452
rect 17736 19392 17800 19396
rect 17816 19452 17880 19456
rect 17816 19396 17820 19452
rect 17820 19396 17876 19452
rect 17876 19396 17880 19452
rect 17816 19392 17880 19396
rect 17896 19452 17960 19456
rect 17896 19396 17900 19452
rect 17900 19396 17956 19452
rect 17956 19396 17960 19452
rect 17896 19392 17960 19396
rect 17976 19452 18040 19456
rect 17976 19396 17980 19452
rect 17980 19396 18036 19452
rect 18036 19396 18040 19452
rect 17976 19392 18040 19396
rect 4416 18908 4480 18912
rect 4416 18852 4420 18908
rect 4420 18852 4476 18908
rect 4476 18852 4480 18908
rect 4416 18848 4480 18852
rect 4496 18908 4560 18912
rect 4496 18852 4500 18908
rect 4500 18852 4556 18908
rect 4556 18852 4560 18908
rect 4496 18848 4560 18852
rect 4576 18908 4640 18912
rect 4576 18852 4580 18908
rect 4580 18852 4636 18908
rect 4636 18852 4640 18908
rect 4576 18848 4640 18852
rect 4656 18908 4720 18912
rect 4656 18852 4660 18908
rect 4660 18852 4716 18908
rect 4716 18852 4720 18908
rect 4656 18848 4720 18852
rect 9744 18908 9808 18912
rect 9744 18852 9748 18908
rect 9748 18852 9804 18908
rect 9804 18852 9808 18908
rect 9744 18848 9808 18852
rect 9824 18908 9888 18912
rect 9824 18852 9828 18908
rect 9828 18852 9884 18908
rect 9884 18852 9888 18908
rect 9824 18848 9888 18852
rect 9904 18908 9968 18912
rect 9904 18852 9908 18908
rect 9908 18852 9964 18908
rect 9964 18852 9968 18908
rect 9904 18848 9968 18852
rect 9984 18908 10048 18912
rect 9984 18852 9988 18908
rect 9988 18852 10044 18908
rect 10044 18852 10048 18908
rect 9984 18848 10048 18852
rect 15072 18908 15136 18912
rect 15072 18852 15076 18908
rect 15076 18852 15132 18908
rect 15132 18852 15136 18908
rect 15072 18848 15136 18852
rect 15152 18908 15216 18912
rect 15152 18852 15156 18908
rect 15156 18852 15212 18908
rect 15212 18852 15216 18908
rect 15152 18848 15216 18852
rect 15232 18908 15296 18912
rect 15232 18852 15236 18908
rect 15236 18852 15292 18908
rect 15292 18852 15296 18908
rect 15232 18848 15296 18852
rect 15312 18908 15376 18912
rect 15312 18852 15316 18908
rect 15316 18852 15372 18908
rect 15372 18852 15376 18908
rect 15312 18848 15376 18852
rect 20400 18908 20464 18912
rect 20400 18852 20404 18908
rect 20404 18852 20460 18908
rect 20460 18852 20464 18908
rect 20400 18848 20464 18852
rect 20480 18908 20544 18912
rect 20480 18852 20484 18908
rect 20484 18852 20540 18908
rect 20540 18852 20544 18908
rect 20480 18848 20544 18852
rect 20560 18908 20624 18912
rect 20560 18852 20564 18908
rect 20564 18852 20620 18908
rect 20620 18852 20624 18908
rect 20560 18848 20624 18852
rect 20640 18908 20704 18912
rect 20640 18852 20644 18908
rect 20644 18852 20700 18908
rect 20700 18852 20704 18908
rect 20640 18848 20704 18852
rect 7080 18364 7144 18368
rect 7080 18308 7084 18364
rect 7084 18308 7140 18364
rect 7140 18308 7144 18364
rect 7080 18304 7144 18308
rect 7160 18364 7224 18368
rect 7160 18308 7164 18364
rect 7164 18308 7220 18364
rect 7220 18308 7224 18364
rect 7160 18304 7224 18308
rect 7240 18364 7304 18368
rect 7240 18308 7244 18364
rect 7244 18308 7300 18364
rect 7300 18308 7304 18364
rect 7240 18304 7304 18308
rect 7320 18364 7384 18368
rect 7320 18308 7324 18364
rect 7324 18308 7380 18364
rect 7380 18308 7384 18364
rect 7320 18304 7384 18308
rect 12408 18364 12472 18368
rect 12408 18308 12412 18364
rect 12412 18308 12468 18364
rect 12468 18308 12472 18364
rect 12408 18304 12472 18308
rect 12488 18364 12552 18368
rect 12488 18308 12492 18364
rect 12492 18308 12548 18364
rect 12548 18308 12552 18364
rect 12488 18304 12552 18308
rect 12568 18364 12632 18368
rect 12568 18308 12572 18364
rect 12572 18308 12628 18364
rect 12628 18308 12632 18364
rect 12568 18304 12632 18308
rect 12648 18364 12712 18368
rect 12648 18308 12652 18364
rect 12652 18308 12708 18364
rect 12708 18308 12712 18364
rect 12648 18304 12712 18308
rect 17736 18364 17800 18368
rect 17736 18308 17740 18364
rect 17740 18308 17796 18364
rect 17796 18308 17800 18364
rect 17736 18304 17800 18308
rect 17816 18364 17880 18368
rect 17816 18308 17820 18364
rect 17820 18308 17876 18364
rect 17876 18308 17880 18364
rect 17816 18304 17880 18308
rect 17896 18364 17960 18368
rect 17896 18308 17900 18364
rect 17900 18308 17956 18364
rect 17956 18308 17960 18364
rect 17896 18304 17960 18308
rect 17976 18364 18040 18368
rect 17976 18308 17980 18364
rect 17980 18308 18036 18364
rect 18036 18308 18040 18364
rect 17976 18304 18040 18308
rect 4416 17820 4480 17824
rect 4416 17764 4420 17820
rect 4420 17764 4476 17820
rect 4476 17764 4480 17820
rect 4416 17760 4480 17764
rect 4496 17820 4560 17824
rect 4496 17764 4500 17820
rect 4500 17764 4556 17820
rect 4556 17764 4560 17820
rect 4496 17760 4560 17764
rect 4576 17820 4640 17824
rect 4576 17764 4580 17820
rect 4580 17764 4636 17820
rect 4636 17764 4640 17820
rect 4576 17760 4640 17764
rect 4656 17820 4720 17824
rect 4656 17764 4660 17820
rect 4660 17764 4716 17820
rect 4716 17764 4720 17820
rect 4656 17760 4720 17764
rect 9744 17820 9808 17824
rect 9744 17764 9748 17820
rect 9748 17764 9804 17820
rect 9804 17764 9808 17820
rect 9744 17760 9808 17764
rect 9824 17820 9888 17824
rect 9824 17764 9828 17820
rect 9828 17764 9884 17820
rect 9884 17764 9888 17820
rect 9824 17760 9888 17764
rect 9904 17820 9968 17824
rect 9904 17764 9908 17820
rect 9908 17764 9964 17820
rect 9964 17764 9968 17820
rect 9904 17760 9968 17764
rect 9984 17820 10048 17824
rect 9984 17764 9988 17820
rect 9988 17764 10044 17820
rect 10044 17764 10048 17820
rect 9984 17760 10048 17764
rect 15072 17820 15136 17824
rect 15072 17764 15076 17820
rect 15076 17764 15132 17820
rect 15132 17764 15136 17820
rect 15072 17760 15136 17764
rect 15152 17820 15216 17824
rect 15152 17764 15156 17820
rect 15156 17764 15212 17820
rect 15212 17764 15216 17820
rect 15152 17760 15216 17764
rect 15232 17820 15296 17824
rect 15232 17764 15236 17820
rect 15236 17764 15292 17820
rect 15292 17764 15296 17820
rect 15232 17760 15296 17764
rect 15312 17820 15376 17824
rect 15312 17764 15316 17820
rect 15316 17764 15372 17820
rect 15372 17764 15376 17820
rect 15312 17760 15376 17764
rect 20400 17820 20464 17824
rect 20400 17764 20404 17820
rect 20404 17764 20460 17820
rect 20460 17764 20464 17820
rect 20400 17760 20464 17764
rect 20480 17820 20544 17824
rect 20480 17764 20484 17820
rect 20484 17764 20540 17820
rect 20540 17764 20544 17820
rect 20480 17760 20544 17764
rect 20560 17820 20624 17824
rect 20560 17764 20564 17820
rect 20564 17764 20620 17820
rect 20620 17764 20624 17820
rect 20560 17760 20624 17764
rect 20640 17820 20704 17824
rect 20640 17764 20644 17820
rect 20644 17764 20700 17820
rect 20700 17764 20704 17820
rect 20640 17760 20704 17764
rect 7080 17276 7144 17280
rect 7080 17220 7084 17276
rect 7084 17220 7140 17276
rect 7140 17220 7144 17276
rect 7080 17216 7144 17220
rect 7160 17276 7224 17280
rect 7160 17220 7164 17276
rect 7164 17220 7220 17276
rect 7220 17220 7224 17276
rect 7160 17216 7224 17220
rect 7240 17276 7304 17280
rect 7240 17220 7244 17276
rect 7244 17220 7300 17276
rect 7300 17220 7304 17276
rect 7240 17216 7304 17220
rect 7320 17276 7384 17280
rect 7320 17220 7324 17276
rect 7324 17220 7380 17276
rect 7380 17220 7384 17276
rect 7320 17216 7384 17220
rect 12408 17276 12472 17280
rect 12408 17220 12412 17276
rect 12412 17220 12468 17276
rect 12468 17220 12472 17276
rect 12408 17216 12472 17220
rect 12488 17276 12552 17280
rect 12488 17220 12492 17276
rect 12492 17220 12548 17276
rect 12548 17220 12552 17276
rect 12488 17216 12552 17220
rect 12568 17276 12632 17280
rect 12568 17220 12572 17276
rect 12572 17220 12628 17276
rect 12628 17220 12632 17276
rect 12568 17216 12632 17220
rect 12648 17276 12712 17280
rect 12648 17220 12652 17276
rect 12652 17220 12708 17276
rect 12708 17220 12712 17276
rect 12648 17216 12712 17220
rect 17736 17276 17800 17280
rect 17736 17220 17740 17276
rect 17740 17220 17796 17276
rect 17796 17220 17800 17276
rect 17736 17216 17800 17220
rect 17816 17276 17880 17280
rect 17816 17220 17820 17276
rect 17820 17220 17876 17276
rect 17876 17220 17880 17276
rect 17816 17216 17880 17220
rect 17896 17276 17960 17280
rect 17896 17220 17900 17276
rect 17900 17220 17956 17276
rect 17956 17220 17960 17276
rect 17896 17216 17960 17220
rect 17976 17276 18040 17280
rect 17976 17220 17980 17276
rect 17980 17220 18036 17276
rect 18036 17220 18040 17276
rect 17976 17216 18040 17220
rect 4416 16732 4480 16736
rect 4416 16676 4420 16732
rect 4420 16676 4476 16732
rect 4476 16676 4480 16732
rect 4416 16672 4480 16676
rect 4496 16732 4560 16736
rect 4496 16676 4500 16732
rect 4500 16676 4556 16732
rect 4556 16676 4560 16732
rect 4496 16672 4560 16676
rect 4576 16732 4640 16736
rect 4576 16676 4580 16732
rect 4580 16676 4636 16732
rect 4636 16676 4640 16732
rect 4576 16672 4640 16676
rect 4656 16732 4720 16736
rect 4656 16676 4660 16732
rect 4660 16676 4716 16732
rect 4716 16676 4720 16732
rect 4656 16672 4720 16676
rect 9744 16732 9808 16736
rect 9744 16676 9748 16732
rect 9748 16676 9804 16732
rect 9804 16676 9808 16732
rect 9744 16672 9808 16676
rect 9824 16732 9888 16736
rect 9824 16676 9828 16732
rect 9828 16676 9884 16732
rect 9884 16676 9888 16732
rect 9824 16672 9888 16676
rect 9904 16732 9968 16736
rect 9904 16676 9908 16732
rect 9908 16676 9964 16732
rect 9964 16676 9968 16732
rect 9904 16672 9968 16676
rect 9984 16732 10048 16736
rect 9984 16676 9988 16732
rect 9988 16676 10044 16732
rect 10044 16676 10048 16732
rect 9984 16672 10048 16676
rect 15072 16732 15136 16736
rect 15072 16676 15076 16732
rect 15076 16676 15132 16732
rect 15132 16676 15136 16732
rect 15072 16672 15136 16676
rect 15152 16732 15216 16736
rect 15152 16676 15156 16732
rect 15156 16676 15212 16732
rect 15212 16676 15216 16732
rect 15152 16672 15216 16676
rect 15232 16732 15296 16736
rect 15232 16676 15236 16732
rect 15236 16676 15292 16732
rect 15292 16676 15296 16732
rect 15232 16672 15296 16676
rect 15312 16732 15376 16736
rect 15312 16676 15316 16732
rect 15316 16676 15372 16732
rect 15372 16676 15376 16732
rect 15312 16672 15376 16676
rect 20400 16732 20464 16736
rect 20400 16676 20404 16732
rect 20404 16676 20460 16732
rect 20460 16676 20464 16732
rect 20400 16672 20464 16676
rect 20480 16732 20544 16736
rect 20480 16676 20484 16732
rect 20484 16676 20540 16732
rect 20540 16676 20544 16732
rect 20480 16672 20544 16676
rect 20560 16732 20624 16736
rect 20560 16676 20564 16732
rect 20564 16676 20620 16732
rect 20620 16676 20624 16732
rect 20560 16672 20624 16676
rect 20640 16732 20704 16736
rect 20640 16676 20644 16732
rect 20644 16676 20700 16732
rect 20700 16676 20704 16732
rect 20640 16672 20704 16676
rect 7080 16188 7144 16192
rect 7080 16132 7084 16188
rect 7084 16132 7140 16188
rect 7140 16132 7144 16188
rect 7080 16128 7144 16132
rect 7160 16188 7224 16192
rect 7160 16132 7164 16188
rect 7164 16132 7220 16188
rect 7220 16132 7224 16188
rect 7160 16128 7224 16132
rect 7240 16188 7304 16192
rect 7240 16132 7244 16188
rect 7244 16132 7300 16188
rect 7300 16132 7304 16188
rect 7240 16128 7304 16132
rect 7320 16188 7384 16192
rect 7320 16132 7324 16188
rect 7324 16132 7380 16188
rect 7380 16132 7384 16188
rect 7320 16128 7384 16132
rect 12408 16188 12472 16192
rect 12408 16132 12412 16188
rect 12412 16132 12468 16188
rect 12468 16132 12472 16188
rect 12408 16128 12472 16132
rect 12488 16188 12552 16192
rect 12488 16132 12492 16188
rect 12492 16132 12548 16188
rect 12548 16132 12552 16188
rect 12488 16128 12552 16132
rect 12568 16188 12632 16192
rect 12568 16132 12572 16188
rect 12572 16132 12628 16188
rect 12628 16132 12632 16188
rect 12568 16128 12632 16132
rect 12648 16188 12712 16192
rect 12648 16132 12652 16188
rect 12652 16132 12708 16188
rect 12708 16132 12712 16188
rect 12648 16128 12712 16132
rect 17736 16188 17800 16192
rect 17736 16132 17740 16188
rect 17740 16132 17796 16188
rect 17796 16132 17800 16188
rect 17736 16128 17800 16132
rect 17816 16188 17880 16192
rect 17816 16132 17820 16188
rect 17820 16132 17876 16188
rect 17876 16132 17880 16188
rect 17816 16128 17880 16132
rect 17896 16188 17960 16192
rect 17896 16132 17900 16188
rect 17900 16132 17956 16188
rect 17956 16132 17960 16188
rect 17896 16128 17960 16132
rect 17976 16188 18040 16192
rect 17976 16132 17980 16188
rect 17980 16132 18036 16188
rect 18036 16132 18040 16188
rect 17976 16128 18040 16132
rect 4416 15644 4480 15648
rect 4416 15588 4420 15644
rect 4420 15588 4476 15644
rect 4476 15588 4480 15644
rect 4416 15584 4480 15588
rect 4496 15644 4560 15648
rect 4496 15588 4500 15644
rect 4500 15588 4556 15644
rect 4556 15588 4560 15644
rect 4496 15584 4560 15588
rect 4576 15644 4640 15648
rect 4576 15588 4580 15644
rect 4580 15588 4636 15644
rect 4636 15588 4640 15644
rect 4576 15584 4640 15588
rect 4656 15644 4720 15648
rect 4656 15588 4660 15644
rect 4660 15588 4716 15644
rect 4716 15588 4720 15644
rect 4656 15584 4720 15588
rect 9744 15644 9808 15648
rect 9744 15588 9748 15644
rect 9748 15588 9804 15644
rect 9804 15588 9808 15644
rect 9744 15584 9808 15588
rect 9824 15644 9888 15648
rect 9824 15588 9828 15644
rect 9828 15588 9884 15644
rect 9884 15588 9888 15644
rect 9824 15584 9888 15588
rect 9904 15644 9968 15648
rect 9904 15588 9908 15644
rect 9908 15588 9964 15644
rect 9964 15588 9968 15644
rect 9904 15584 9968 15588
rect 9984 15644 10048 15648
rect 9984 15588 9988 15644
rect 9988 15588 10044 15644
rect 10044 15588 10048 15644
rect 9984 15584 10048 15588
rect 15072 15644 15136 15648
rect 15072 15588 15076 15644
rect 15076 15588 15132 15644
rect 15132 15588 15136 15644
rect 15072 15584 15136 15588
rect 15152 15644 15216 15648
rect 15152 15588 15156 15644
rect 15156 15588 15212 15644
rect 15212 15588 15216 15644
rect 15152 15584 15216 15588
rect 15232 15644 15296 15648
rect 15232 15588 15236 15644
rect 15236 15588 15292 15644
rect 15292 15588 15296 15644
rect 15232 15584 15296 15588
rect 15312 15644 15376 15648
rect 15312 15588 15316 15644
rect 15316 15588 15372 15644
rect 15372 15588 15376 15644
rect 15312 15584 15376 15588
rect 20400 15644 20464 15648
rect 20400 15588 20404 15644
rect 20404 15588 20460 15644
rect 20460 15588 20464 15644
rect 20400 15584 20464 15588
rect 20480 15644 20544 15648
rect 20480 15588 20484 15644
rect 20484 15588 20540 15644
rect 20540 15588 20544 15644
rect 20480 15584 20544 15588
rect 20560 15644 20624 15648
rect 20560 15588 20564 15644
rect 20564 15588 20620 15644
rect 20620 15588 20624 15644
rect 20560 15584 20624 15588
rect 20640 15644 20704 15648
rect 20640 15588 20644 15644
rect 20644 15588 20700 15644
rect 20700 15588 20704 15644
rect 20640 15584 20704 15588
rect 7080 15100 7144 15104
rect 7080 15044 7084 15100
rect 7084 15044 7140 15100
rect 7140 15044 7144 15100
rect 7080 15040 7144 15044
rect 7160 15100 7224 15104
rect 7160 15044 7164 15100
rect 7164 15044 7220 15100
rect 7220 15044 7224 15100
rect 7160 15040 7224 15044
rect 7240 15100 7304 15104
rect 7240 15044 7244 15100
rect 7244 15044 7300 15100
rect 7300 15044 7304 15100
rect 7240 15040 7304 15044
rect 7320 15100 7384 15104
rect 7320 15044 7324 15100
rect 7324 15044 7380 15100
rect 7380 15044 7384 15100
rect 7320 15040 7384 15044
rect 12408 15100 12472 15104
rect 12408 15044 12412 15100
rect 12412 15044 12468 15100
rect 12468 15044 12472 15100
rect 12408 15040 12472 15044
rect 12488 15100 12552 15104
rect 12488 15044 12492 15100
rect 12492 15044 12548 15100
rect 12548 15044 12552 15100
rect 12488 15040 12552 15044
rect 12568 15100 12632 15104
rect 12568 15044 12572 15100
rect 12572 15044 12628 15100
rect 12628 15044 12632 15100
rect 12568 15040 12632 15044
rect 12648 15100 12712 15104
rect 12648 15044 12652 15100
rect 12652 15044 12708 15100
rect 12708 15044 12712 15100
rect 12648 15040 12712 15044
rect 17736 15100 17800 15104
rect 17736 15044 17740 15100
rect 17740 15044 17796 15100
rect 17796 15044 17800 15100
rect 17736 15040 17800 15044
rect 17816 15100 17880 15104
rect 17816 15044 17820 15100
rect 17820 15044 17876 15100
rect 17876 15044 17880 15100
rect 17816 15040 17880 15044
rect 17896 15100 17960 15104
rect 17896 15044 17900 15100
rect 17900 15044 17956 15100
rect 17956 15044 17960 15100
rect 17896 15040 17960 15044
rect 17976 15100 18040 15104
rect 17976 15044 17980 15100
rect 17980 15044 18036 15100
rect 18036 15044 18040 15100
rect 17976 15040 18040 15044
rect 4416 14556 4480 14560
rect 4416 14500 4420 14556
rect 4420 14500 4476 14556
rect 4476 14500 4480 14556
rect 4416 14496 4480 14500
rect 4496 14556 4560 14560
rect 4496 14500 4500 14556
rect 4500 14500 4556 14556
rect 4556 14500 4560 14556
rect 4496 14496 4560 14500
rect 4576 14556 4640 14560
rect 4576 14500 4580 14556
rect 4580 14500 4636 14556
rect 4636 14500 4640 14556
rect 4576 14496 4640 14500
rect 4656 14556 4720 14560
rect 4656 14500 4660 14556
rect 4660 14500 4716 14556
rect 4716 14500 4720 14556
rect 4656 14496 4720 14500
rect 9744 14556 9808 14560
rect 9744 14500 9748 14556
rect 9748 14500 9804 14556
rect 9804 14500 9808 14556
rect 9744 14496 9808 14500
rect 9824 14556 9888 14560
rect 9824 14500 9828 14556
rect 9828 14500 9884 14556
rect 9884 14500 9888 14556
rect 9824 14496 9888 14500
rect 9904 14556 9968 14560
rect 9904 14500 9908 14556
rect 9908 14500 9964 14556
rect 9964 14500 9968 14556
rect 9904 14496 9968 14500
rect 9984 14556 10048 14560
rect 9984 14500 9988 14556
rect 9988 14500 10044 14556
rect 10044 14500 10048 14556
rect 9984 14496 10048 14500
rect 15072 14556 15136 14560
rect 15072 14500 15076 14556
rect 15076 14500 15132 14556
rect 15132 14500 15136 14556
rect 15072 14496 15136 14500
rect 15152 14556 15216 14560
rect 15152 14500 15156 14556
rect 15156 14500 15212 14556
rect 15212 14500 15216 14556
rect 15152 14496 15216 14500
rect 15232 14556 15296 14560
rect 15232 14500 15236 14556
rect 15236 14500 15292 14556
rect 15292 14500 15296 14556
rect 15232 14496 15296 14500
rect 15312 14556 15376 14560
rect 15312 14500 15316 14556
rect 15316 14500 15372 14556
rect 15372 14500 15376 14556
rect 15312 14496 15376 14500
rect 20400 14556 20464 14560
rect 20400 14500 20404 14556
rect 20404 14500 20460 14556
rect 20460 14500 20464 14556
rect 20400 14496 20464 14500
rect 20480 14556 20544 14560
rect 20480 14500 20484 14556
rect 20484 14500 20540 14556
rect 20540 14500 20544 14556
rect 20480 14496 20544 14500
rect 20560 14556 20624 14560
rect 20560 14500 20564 14556
rect 20564 14500 20620 14556
rect 20620 14500 20624 14556
rect 20560 14496 20624 14500
rect 20640 14556 20704 14560
rect 20640 14500 20644 14556
rect 20644 14500 20700 14556
rect 20700 14500 20704 14556
rect 20640 14496 20704 14500
rect 7080 14012 7144 14016
rect 7080 13956 7084 14012
rect 7084 13956 7140 14012
rect 7140 13956 7144 14012
rect 7080 13952 7144 13956
rect 7160 14012 7224 14016
rect 7160 13956 7164 14012
rect 7164 13956 7220 14012
rect 7220 13956 7224 14012
rect 7160 13952 7224 13956
rect 7240 14012 7304 14016
rect 7240 13956 7244 14012
rect 7244 13956 7300 14012
rect 7300 13956 7304 14012
rect 7240 13952 7304 13956
rect 7320 14012 7384 14016
rect 7320 13956 7324 14012
rect 7324 13956 7380 14012
rect 7380 13956 7384 14012
rect 7320 13952 7384 13956
rect 12408 14012 12472 14016
rect 12408 13956 12412 14012
rect 12412 13956 12468 14012
rect 12468 13956 12472 14012
rect 12408 13952 12472 13956
rect 12488 14012 12552 14016
rect 12488 13956 12492 14012
rect 12492 13956 12548 14012
rect 12548 13956 12552 14012
rect 12488 13952 12552 13956
rect 12568 14012 12632 14016
rect 12568 13956 12572 14012
rect 12572 13956 12628 14012
rect 12628 13956 12632 14012
rect 12568 13952 12632 13956
rect 12648 14012 12712 14016
rect 12648 13956 12652 14012
rect 12652 13956 12708 14012
rect 12708 13956 12712 14012
rect 12648 13952 12712 13956
rect 17736 14012 17800 14016
rect 17736 13956 17740 14012
rect 17740 13956 17796 14012
rect 17796 13956 17800 14012
rect 17736 13952 17800 13956
rect 17816 14012 17880 14016
rect 17816 13956 17820 14012
rect 17820 13956 17876 14012
rect 17876 13956 17880 14012
rect 17816 13952 17880 13956
rect 17896 14012 17960 14016
rect 17896 13956 17900 14012
rect 17900 13956 17956 14012
rect 17956 13956 17960 14012
rect 17896 13952 17960 13956
rect 17976 14012 18040 14016
rect 17976 13956 17980 14012
rect 17980 13956 18036 14012
rect 18036 13956 18040 14012
rect 17976 13952 18040 13956
rect 4416 13468 4480 13472
rect 4416 13412 4420 13468
rect 4420 13412 4476 13468
rect 4476 13412 4480 13468
rect 4416 13408 4480 13412
rect 4496 13468 4560 13472
rect 4496 13412 4500 13468
rect 4500 13412 4556 13468
rect 4556 13412 4560 13468
rect 4496 13408 4560 13412
rect 4576 13468 4640 13472
rect 4576 13412 4580 13468
rect 4580 13412 4636 13468
rect 4636 13412 4640 13468
rect 4576 13408 4640 13412
rect 4656 13468 4720 13472
rect 4656 13412 4660 13468
rect 4660 13412 4716 13468
rect 4716 13412 4720 13468
rect 4656 13408 4720 13412
rect 9744 13468 9808 13472
rect 9744 13412 9748 13468
rect 9748 13412 9804 13468
rect 9804 13412 9808 13468
rect 9744 13408 9808 13412
rect 9824 13468 9888 13472
rect 9824 13412 9828 13468
rect 9828 13412 9884 13468
rect 9884 13412 9888 13468
rect 9824 13408 9888 13412
rect 9904 13468 9968 13472
rect 9904 13412 9908 13468
rect 9908 13412 9964 13468
rect 9964 13412 9968 13468
rect 9904 13408 9968 13412
rect 9984 13468 10048 13472
rect 9984 13412 9988 13468
rect 9988 13412 10044 13468
rect 10044 13412 10048 13468
rect 9984 13408 10048 13412
rect 15072 13468 15136 13472
rect 15072 13412 15076 13468
rect 15076 13412 15132 13468
rect 15132 13412 15136 13468
rect 15072 13408 15136 13412
rect 15152 13468 15216 13472
rect 15152 13412 15156 13468
rect 15156 13412 15212 13468
rect 15212 13412 15216 13468
rect 15152 13408 15216 13412
rect 15232 13468 15296 13472
rect 15232 13412 15236 13468
rect 15236 13412 15292 13468
rect 15292 13412 15296 13468
rect 15232 13408 15296 13412
rect 15312 13468 15376 13472
rect 15312 13412 15316 13468
rect 15316 13412 15372 13468
rect 15372 13412 15376 13468
rect 15312 13408 15376 13412
rect 20400 13468 20464 13472
rect 20400 13412 20404 13468
rect 20404 13412 20460 13468
rect 20460 13412 20464 13468
rect 20400 13408 20464 13412
rect 20480 13468 20544 13472
rect 20480 13412 20484 13468
rect 20484 13412 20540 13468
rect 20540 13412 20544 13468
rect 20480 13408 20544 13412
rect 20560 13468 20624 13472
rect 20560 13412 20564 13468
rect 20564 13412 20620 13468
rect 20620 13412 20624 13468
rect 20560 13408 20624 13412
rect 20640 13468 20704 13472
rect 20640 13412 20644 13468
rect 20644 13412 20700 13468
rect 20700 13412 20704 13468
rect 20640 13408 20704 13412
rect 7080 12924 7144 12928
rect 7080 12868 7084 12924
rect 7084 12868 7140 12924
rect 7140 12868 7144 12924
rect 7080 12864 7144 12868
rect 7160 12924 7224 12928
rect 7160 12868 7164 12924
rect 7164 12868 7220 12924
rect 7220 12868 7224 12924
rect 7160 12864 7224 12868
rect 7240 12924 7304 12928
rect 7240 12868 7244 12924
rect 7244 12868 7300 12924
rect 7300 12868 7304 12924
rect 7240 12864 7304 12868
rect 7320 12924 7384 12928
rect 7320 12868 7324 12924
rect 7324 12868 7380 12924
rect 7380 12868 7384 12924
rect 7320 12864 7384 12868
rect 12408 12924 12472 12928
rect 12408 12868 12412 12924
rect 12412 12868 12468 12924
rect 12468 12868 12472 12924
rect 12408 12864 12472 12868
rect 12488 12924 12552 12928
rect 12488 12868 12492 12924
rect 12492 12868 12548 12924
rect 12548 12868 12552 12924
rect 12488 12864 12552 12868
rect 12568 12924 12632 12928
rect 12568 12868 12572 12924
rect 12572 12868 12628 12924
rect 12628 12868 12632 12924
rect 12568 12864 12632 12868
rect 12648 12924 12712 12928
rect 12648 12868 12652 12924
rect 12652 12868 12708 12924
rect 12708 12868 12712 12924
rect 12648 12864 12712 12868
rect 17736 12924 17800 12928
rect 17736 12868 17740 12924
rect 17740 12868 17796 12924
rect 17796 12868 17800 12924
rect 17736 12864 17800 12868
rect 17816 12924 17880 12928
rect 17816 12868 17820 12924
rect 17820 12868 17876 12924
rect 17876 12868 17880 12924
rect 17816 12864 17880 12868
rect 17896 12924 17960 12928
rect 17896 12868 17900 12924
rect 17900 12868 17956 12924
rect 17956 12868 17960 12924
rect 17896 12864 17960 12868
rect 17976 12924 18040 12928
rect 17976 12868 17980 12924
rect 17980 12868 18036 12924
rect 18036 12868 18040 12924
rect 17976 12864 18040 12868
rect 4416 12380 4480 12384
rect 4416 12324 4420 12380
rect 4420 12324 4476 12380
rect 4476 12324 4480 12380
rect 4416 12320 4480 12324
rect 4496 12380 4560 12384
rect 4496 12324 4500 12380
rect 4500 12324 4556 12380
rect 4556 12324 4560 12380
rect 4496 12320 4560 12324
rect 4576 12380 4640 12384
rect 4576 12324 4580 12380
rect 4580 12324 4636 12380
rect 4636 12324 4640 12380
rect 4576 12320 4640 12324
rect 4656 12380 4720 12384
rect 4656 12324 4660 12380
rect 4660 12324 4716 12380
rect 4716 12324 4720 12380
rect 4656 12320 4720 12324
rect 9744 12380 9808 12384
rect 9744 12324 9748 12380
rect 9748 12324 9804 12380
rect 9804 12324 9808 12380
rect 9744 12320 9808 12324
rect 9824 12380 9888 12384
rect 9824 12324 9828 12380
rect 9828 12324 9884 12380
rect 9884 12324 9888 12380
rect 9824 12320 9888 12324
rect 9904 12380 9968 12384
rect 9904 12324 9908 12380
rect 9908 12324 9964 12380
rect 9964 12324 9968 12380
rect 9904 12320 9968 12324
rect 9984 12380 10048 12384
rect 9984 12324 9988 12380
rect 9988 12324 10044 12380
rect 10044 12324 10048 12380
rect 9984 12320 10048 12324
rect 15072 12380 15136 12384
rect 15072 12324 15076 12380
rect 15076 12324 15132 12380
rect 15132 12324 15136 12380
rect 15072 12320 15136 12324
rect 15152 12380 15216 12384
rect 15152 12324 15156 12380
rect 15156 12324 15212 12380
rect 15212 12324 15216 12380
rect 15152 12320 15216 12324
rect 15232 12380 15296 12384
rect 15232 12324 15236 12380
rect 15236 12324 15292 12380
rect 15292 12324 15296 12380
rect 15232 12320 15296 12324
rect 15312 12380 15376 12384
rect 15312 12324 15316 12380
rect 15316 12324 15372 12380
rect 15372 12324 15376 12380
rect 15312 12320 15376 12324
rect 20400 12380 20464 12384
rect 20400 12324 20404 12380
rect 20404 12324 20460 12380
rect 20460 12324 20464 12380
rect 20400 12320 20464 12324
rect 20480 12380 20544 12384
rect 20480 12324 20484 12380
rect 20484 12324 20540 12380
rect 20540 12324 20544 12380
rect 20480 12320 20544 12324
rect 20560 12380 20624 12384
rect 20560 12324 20564 12380
rect 20564 12324 20620 12380
rect 20620 12324 20624 12380
rect 20560 12320 20624 12324
rect 20640 12380 20704 12384
rect 20640 12324 20644 12380
rect 20644 12324 20700 12380
rect 20700 12324 20704 12380
rect 20640 12320 20704 12324
rect 7080 11836 7144 11840
rect 7080 11780 7084 11836
rect 7084 11780 7140 11836
rect 7140 11780 7144 11836
rect 7080 11776 7144 11780
rect 7160 11836 7224 11840
rect 7160 11780 7164 11836
rect 7164 11780 7220 11836
rect 7220 11780 7224 11836
rect 7160 11776 7224 11780
rect 7240 11836 7304 11840
rect 7240 11780 7244 11836
rect 7244 11780 7300 11836
rect 7300 11780 7304 11836
rect 7240 11776 7304 11780
rect 7320 11836 7384 11840
rect 7320 11780 7324 11836
rect 7324 11780 7380 11836
rect 7380 11780 7384 11836
rect 7320 11776 7384 11780
rect 12408 11836 12472 11840
rect 12408 11780 12412 11836
rect 12412 11780 12468 11836
rect 12468 11780 12472 11836
rect 12408 11776 12472 11780
rect 12488 11836 12552 11840
rect 12488 11780 12492 11836
rect 12492 11780 12548 11836
rect 12548 11780 12552 11836
rect 12488 11776 12552 11780
rect 12568 11836 12632 11840
rect 12568 11780 12572 11836
rect 12572 11780 12628 11836
rect 12628 11780 12632 11836
rect 12568 11776 12632 11780
rect 12648 11836 12712 11840
rect 12648 11780 12652 11836
rect 12652 11780 12708 11836
rect 12708 11780 12712 11836
rect 12648 11776 12712 11780
rect 17736 11836 17800 11840
rect 17736 11780 17740 11836
rect 17740 11780 17796 11836
rect 17796 11780 17800 11836
rect 17736 11776 17800 11780
rect 17816 11836 17880 11840
rect 17816 11780 17820 11836
rect 17820 11780 17876 11836
rect 17876 11780 17880 11836
rect 17816 11776 17880 11780
rect 17896 11836 17960 11840
rect 17896 11780 17900 11836
rect 17900 11780 17956 11836
rect 17956 11780 17960 11836
rect 17896 11776 17960 11780
rect 17976 11836 18040 11840
rect 17976 11780 17980 11836
rect 17980 11780 18036 11836
rect 18036 11780 18040 11836
rect 17976 11776 18040 11780
rect 4416 11292 4480 11296
rect 4416 11236 4420 11292
rect 4420 11236 4476 11292
rect 4476 11236 4480 11292
rect 4416 11232 4480 11236
rect 4496 11292 4560 11296
rect 4496 11236 4500 11292
rect 4500 11236 4556 11292
rect 4556 11236 4560 11292
rect 4496 11232 4560 11236
rect 4576 11292 4640 11296
rect 4576 11236 4580 11292
rect 4580 11236 4636 11292
rect 4636 11236 4640 11292
rect 4576 11232 4640 11236
rect 4656 11292 4720 11296
rect 4656 11236 4660 11292
rect 4660 11236 4716 11292
rect 4716 11236 4720 11292
rect 4656 11232 4720 11236
rect 9744 11292 9808 11296
rect 9744 11236 9748 11292
rect 9748 11236 9804 11292
rect 9804 11236 9808 11292
rect 9744 11232 9808 11236
rect 9824 11292 9888 11296
rect 9824 11236 9828 11292
rect 9828 11236 9884 11292
rect 9884 11236 9888 11292
rect 9824 11232 9888 11236
rect 9904 11292 9968 11296
rect 9904 11236 9908 11292
rect 9908 11236 9964 11292
rect 9964 11236 9968 11292
rect 9904 11232 9968 11236
rect 9984 11292 10048 11296
rect 9984 11236 9988 11292
rect 9988 11236 10044 11292
rect 10044 11236 10048 11292
rect 9984 11232 10048 11236
rect 15072 11292 15136 11296
rect 15072 11236 15076 11292
rect 15076 11236 15132 11292
rect 15132 11236 15136 11292
rect 15072 11232 15136 11236
rect 15152 11292 15216 11296
rect 15152 11236 15156 11292
rect 15156 11236 15212 11292
rect 15212 11236 15216 11292
rect 15152 11232 15216 11236
rect 15232 11292 15296 11296
rect 15232 11236 15236 11292
rect 15236 11236 15292 11292
rect 15292 11236 15296 11292
rect 15232 11232 15296 11236
rect 15312 11292 15376 11296
rect 15312 11236 15316 11292
rect 15316 11236 15372 11292
rect 15372 11236 15376 11292
rect 15312 11232 15376 11236
rect 20400 11292 20464 11296
rect 20400 11236 20404 11292
rect 20404 11236 20460 11292
rect 20460 11236 20464 11292
rect 20400 11232 20464 11236
rect 20480 11292 20544 11296
rect 20480 11236 20484 11292
rect 20484 11236 20540 11292
rect 20540 11236 20544 11292
rect 20480 11232 20544 11236
rect 20560 11292 20624 11296
rect 20560 11236 20564 11292
rect 20564 11236 20620 11292
rect 20620 11236 20624 11292
rect 20560 11232 20624 11236
rect 20640 11292 20704 11296
rect 20640 11236 20644 11292
rect 20644 11236 20700 11292
rect 20700 11236 20704 11292
rect 20640 11232 20704 11236
rect 7080 10748 7144 10752
rect 7080 10692 7084 10748
rect 7084 10692 7140 10748
rect 7140 10692 7144 10748
rect 7080 10688 7144 10692
rect 7160 10748 7224 10752
rect 7160 10692 7164 10748
rect 7164 10692 7220 10748
rect 7220 10692 7224 10748
rect 7160 10688 7224 10692
rect 7240 10748 7304 10752
rect 7240 10692 7244 10748
rect 7244 10692 7300 10748
rect 7300 10692 7304 10748
rect 7240 10688 7304 10692
rect 7320 10748 7384 10752
rect 7320 10692 7324 10748
rect 7324 10692 7380 10748
rect 7380 10692 7384 10748
rect 7320 10688 7384 10692
rect 12408 10748 12472 10752
rect 12408 10692 12412 10748
rect 12412 10692 12468 10748
rect 12468 10692 12472 10748
rect 12408 10688 12472 10692
rect 12488 10748 12552 10752
rect 12488 10692 12492 10748
rect 12492 10692 12548 10748
rect 12548 10692 12552 10748
rect 12488 10688 12552 10692
rect 12568 10748 12632 10752
rect 12568 10692 12572 10748
rect 12572 10692 12628 10748
rect 12628 10692 12632 10748
rect 12568 10688 12632 10692
rect 12648 10748 12712 10752
rect 12648 10692 12652 10748
rect 12652 10692 12708 10748
rect 12708 10692 12712 10748
rect 12648 10688 12712 10692
rect 17736 10748 17800 10752
rect 17736 10692 17740 10748
rect 17740 10692 17796 10748
rect 17796 10692 17800 10748
rect 17736 10688 17800 10692
rect 17816 10748 17880 10752
rect 17816 10692 17820 10748
rect 17820 10692 17876 10748
rect 17876 10692 17880 10748
rect 17816 10688 17880 10692
rect 17896 10748 17960 10752
rect 17896 10692 17900 10748
rect 17900 10692 17956 10748
rect 17956 10692 17960 10748
rect 17896 10688 17960 10692
rect 17976 10748 18040 10752
rect 17976 10692 17980 10748
rect 17980 10692 18036 10748
rect 18036 10692 18040 10748
rect 17976 10688 18040 10692
rect 4416 10204 4480 10208
rect 4416 10148 4420 10204
rect 4420 10148 4476 10204
rect 4476 10148 4480 10204
rect 4416 10144 4480 10148
rect 4496 10204 4560 10208
rect 4496 10148 4500 10204
rect 4500 10148 4556 10204
rect 4556 10148 4560 10204
rect 4496 10144 4560 10148
rect 4576 10204 4640 10208
rect 4576 10148 4580 10204
rect 4580 10148 4636 10204
rect 4636 10148 4640 10204
rect 4576 10144 4640 10148
rect 4656 10204 4720 10208
rect 4656 10148 4660 10204
rect 4660 10148 4716 10204
rect 4716 10148 4720 10204
rect 4656 10144 4720 10148
rect 9744 10204 9808 10208
rect 9744 10148 9748 10204
rect 9748 10148 9804 10204
rect 9804 10148 9808 10204
rect 9744 10144 9808 10148
rect 9824 10204 9888 10208
rect 9824 10148 9828 10204
rect 9828 10148 9884 10204
rect 9884 10148 9888 10204
rect 9824 10144 9888 10148
rect 9904 10204 9968 10208
rect 9904 10148 9908 10204
rect 9908 10148 9964 10204
rect 9964 10148 9968 10204
rect 9904 10144 9968 10148
rect 9984 10204 10048 10208
rect 9984 10148 9988 10204
rect 9988 10148 10044 10204
rect 10044 10148 10048 10204
rect 9984 10144 10048 10148
rect 15072 10204 15136 10208
rect 15072 10148 15076 10204
rect 15076 10148 15132 10204
rect 15132 10148 15136 10204
rect 15072 10144 15136 10148
rect 15152 10204 15216 10208
rect 15152 10148 15156 10204
rect 15156 10148 15212 10204
rect 15212 10148 15216 10204
rect 15152 10144 15216 10148
rect 15232 10204 15296 10208
rect 15232 10148 15236 10204
rect 15236 10148 15292 10204
rect 15292 10148 15296 10204
rect 15232 10144 15296 10148
rect 15312 10204 15376 10208
rect 15312 10148 15316 10204
rect 15316 10148 15372 10204
rect 15372 10148 15376 10204
rect 15312 10144 15376 10148
rect 20400 10204 20464 10208
rect 20400 10148 20404 10204
rect 20404 10148 20460 10204
rect 20460 10148 20464 10204
rect 20400 10144 20464 10148
rect 20480 10204 20544 10208
rect 20480 10148 20484 10204
rect 20484 10148 20540 10204
rect 20540 10148 20544 10204
rect 20480 10144 20544 10148
rect 20560 10204 20624 10208
rect 20560 10148 20564 10204
rect 20564 10148 20620 10204
rect 20620 10148 20624 10204
rect 20560 10144 20624 10148
rect 20640 10204 20704 10208
rect 20640 10148 20644 10204
rect 20644 10148 20700 10204
rect 20700 10148 20704 10204
rect 20640 10144 20704 10148
rect 7080 9660 7144 9664
rect 7080 9604 7084 9660
rect 7084 9604 7140 9660
rect 7140 9604 7144 9660
rect 7080 9600 7144 9604
rect 7160 9660 7224 9664
rect 7160 9604 7164 9660
rect 7164 9604 7220 9660
rect 7220 9604 7224 9660
rect 7160 9600 7224 9604
rect 7240 9660 7304 9664
rect 7240 9604 7244 9660
rect 7244 9604 7300 9660
rect 7300 9604 7304 9660
rect 7240 9600 7304 9604
rect 7320 9660 7384 9664
rect 7320 9604 7324 9660
rect 7324 9604 7380 9660
rect 7380 9604 7384 9660
rect 7320 9600 7384 9604
rect 12408 9660 12472 9664
rect 12408 9604 12412 9660
rect 12412 9604 12468 9660
rect 12468 9604 12472 9660
rect 12408 9600 12472 9604
rect 12488 9660 12552 9664
rect 12488 9604 12492 9660
rect 12492 9604 12548 9660
rect 12548 9604 12552 9660
rect 12488 9600 12552 9604
rect 12568 9660 12632 9664
rect 12568 9604 12572 9660
rect 12572 9604 12628 9660
rect 12628 9604 12632 9660
rect 12568 9600 12632 9604
rect 12648 9660 12712 9664
rect 12648 9604 12652 9660
rect 12652 9604 12708 9660
rect 12708 9604 12712 9660
rect 12648 9600 12712 9604
rect 17736 9660 17800 9664
rect 17736 9604 17740 9660
rect 17740 9604 17796 9660
rect 17796 9604 17800 9660
rect 17736 9600 17800 9604
rect 17816 9660 17880 9664
rect 17816 9604 17820 9660
rect 17820 9604 17876 9660
rect 17876 9604 17880 9660
rect 17816 9600 17880 9604
rect 17896 9660 17960 9664
rect 17896 9604 17900 9660
rect 17900 9604 17956 9660
rect 17956 9604 17960 9660
rect 17896 9600 17960 9604
rect 17976 9660 18040 9664
rect 17976 9604 17980 9660
rect 17980 9604 18036 9660
rect 18036 9604 18040 9660
rect 17976 9600 18040 9604
rect 4416 9116 4480 9120
rect 4416 9060 4420 9116
rect 4420 9060 4476 9116
rect 4476 9060 4480 9116
rect 4416 9056 4480 9060
rect 4496 9116 4560 9120
rect 4496 9060 4500 9116
rect 4500 9060 4556 9116
rect 4556 9060 4560 9116
rect 4496 9056 4560 9060
rect 4576 9116 4640 9120
rect 4576 9060 4580 9116
rect 4580 9060 4636 9116
rect 4636 9060 4640 9116
rect 4576 9056 4640 9060
rect 4656 9116 4720 9120
rect 4656 9060 4660 9116
rect 4660 9060 4716 9116
rect 4716 9060 4720 9116
rect 4656 9056 4720 9060
rect 9744 9116 9808 9120
rect 9744 9060 9748 9116
rect 9748 9060 9804 9116
rect 9804 9060 9808 9116
rect 9744 9056 9808 9060
rect 9824 9116 9888 9120
rect 9824 9060 9828 9116
rect 9828 9060 9884 9116
rect 9884 9060 9888 9116
rect 9824 9056 9888 9060
rect 9904 9116 9968 9120
rect 9904 9060 9908 9116
rect 9908 9060 9964 9116
rect 9964 9060 9968 9116
rect 9904 9056 9968 9060
rect 9984 9116 10048 9120
rect 9984 9060 9988 9116
rect 9988 9060 10044 9116
rect 10044 9060 10048 9116
rect 9984 9056 10048 9060
rect 15072 9116 15136 9120
rect 15072 9060 15076 9116
rect 15076 9060 15132 9116
rect 15132 9060 15136 9116
rect 15072 9056 15136 9060
rect 15152 9116 15216 9120
rect 15152 9060 15156 9116
rect 15156 9060 15212 9116
rect 15212 9060 15216 9116
rect 15152 9056 15216 9060
rect 15232 9116 15296 9120
rect 15232 9060 15236 9116
rect 15236 9060 15292 9116
rect 15292 9060 15296 9116
rect 15232 9056 15296 9060
rect 15312 9116 15376 9120
rect 15312 9060 15316 9116
rect 15316 9060 15372 9116
rect 15372 9060 15376 9116
rect 15312 9056 15376 9060
rect 20400 9116 20464 9120
rect 20400 9060 20404 9116
rect 20404 9060 20460 9116
rect 20460 9060 20464 9116
rect 20400 9056 20464 9060
rect 20480 9116 20544 9120
rect 20480 9060 20484 9116
rect 20484 9060 20540 9116
rect 20540 9060 20544 9116
rect 20480 9056 20544 9060
rect 20560 9116 20624 9120
rect 20560 9060 20564 9116
rect 20564 9060 20620 9116
rect 20620 9060 20624 9116
rect 20560 9056 20624 9060
rect 20640 9116 20704 9120
rect 20640 9060 20644 9116
rect 20644 9060 20700 9116
rect 20700 9060 20704 9116
rect 20640 9056 20704 9060
rect 7080 8572 7144 8576
rect 7080 8516 7084 8572
rect 7084 8516 7140 8572
rect 7140 8516 7144 8572
rect 7080 8512 7144 8516
rect 7160 8572 7224 8576
rect 7160 8516 7164 8572
rect 7164 8516 7220 8572
rect 7220 8516 7224 8572
rect 7160 8512 7224 8516
rect 7240 8572 7304 8576
rect 7240 8516 7244 8572
rect 7244 8516 7300 8572
rect 7300 8516 7304 8572
rect 7240 8512 7304 8516
rect 7320 8572 7384 8576
rect 7320 8516 7324 8572
rect 7324 8516 7380 8572
rect 7380 8516 7384 8572
rect 7320 8512 7384 8516
rect 12408 8572 12472 8576
rect 12408 8516 12412 8572
rect 12412 8516 12468 8572
rect 12468 8516 12472 8572
rect 12408 8512 12472 8516
rect 12488 8572 12552 8576
rect 12488 8516 12492 8572
rect 12492 8516 12548 8572
rect 12548 8516 12552 8572
rect 12488 8512 12552 8516
rect 12568 8572 12632 8576
rect 12568 8516 12572 8572
rect 12572 8516 12628 8572
rect 12628 8516 12632 8572
rect 12568 8512 12632 8516
rect 12648 8572 12712 8576
rect 12648 8516 12652 8572
rect 12652 8516 12708 8572
rect 12708 8516 12712 8572
rect 12648 8512 12712 8516
rect 17736 8572 17800 8576
rect 17736 8516 17740 8572
rect 17740 8516 17796 8572
rect 17796 8516 17800 8572
rect 17736 8512 17800 8516
rect 17816 8572 17880 8576
rect 17816 8516 17820 8572
rect 17820 8516 17876 8572
rect 17876 8516 17880 8572
rect 17816 8512 17880 8516
rect 17896 8572 17960 8576
rect 17896 8516 17900 8572
rect 17900 8516 17956 8572
rect 17956 8516 17960 8572
rect 17896 8512 17960 8516
rect 17976 8572 18040 8576
rect 17976 8516 17980 8572
rect 17980 8516 18036 8572
rect 18036 8516 18040 8572
rect 17976 8512 18040 8516
rect 4416 8028 4480 8032
rect 4416 7972 4420 8028
rect 4420 7972 4476 8028
rect 4476 7972 4480 8028
rect 4416 7968 4480 7972
rect 4496 8028 4560 8032
rect 4496 7972 4500 8028
rect 4500 7972 4556 8028
rect 4556 7972 4560 8028
rect 4496 7968 4560 7972
rect 4576 8028 4640 8032
rect 4576 7972 4580 8028
rect 4580 7972 4636 8028
rect 4636 7972 4640 8028
rect 4576 7968 4640 7972
rect 4656 8028 4720 8032
rect 4656 7972 4660 8028
rect 4660 7972 4716 8028
rect 4716 7972 4720 8028
rect 4656 7968 4720 7972
rect 9744 8028 9808 8032
rect 9744 7972 9748 8028
rect 9748 7972 9804 8028
rect 9804 7972 9808 8028
rect 9744 7968 9808 7972
rect 9824 8028 9888 8032
rect 9824 7972 9828 8028
rect 9828 7972 9884 8028
rect 9884 7972 9888 8028
rect 9824 7968 9888 7972
rect 9904 8028 9968 8032
rect 9904 7972 9908 8028
rect 9908 7972 9964 8028
rect 9964 7972 9968 8028
rect 9904 7968 9968 7972
rect 9984 8028 10048 8032
rect 9984 7972 9988 8028
rect 9988 7972 10044 8028
rect 10044 7972 10048 8028
rect 9984 7968 10048 7972
rect 15072 8028 15136 8032
rect 15072 7972 15076 8028
rect 15076 7972 15132 8028
rect 15132 7972 15136 8028
rect 15072 7968 15136 7972
rect 15152 8028 15216 8032
rect 15152 7972 15156 8028
rect 15156 7972 15212 8028
rect 15212 7972 15216 8028
rect 15152 7968 15216 7972
rect 15232 8028 15296 8032
rect 15232 7972 15236 8028
rect 15236 7972 15292 8028
rect 15292 7972 15296 8028
rect 15232 7968 15296 7972
rect 15312 8028 15376 8032
rect 15312 7972 15316 8028
rect 15316 7972 15372 8028
rect 15372 7972 15376 8028
rect 15312 7968 15376 7972
rect 20400 8028 20464 8032
rect 20400 7972 20404 8028
rect 20404 7972 20460 8028
rect 20460 7972 20464 8028
rect 20400 7968 20464 7972
rect 20480 8028 20544 8032
rect 20480 7972 20484 8028
rect 20484 7972 20540 8028
rect 20540 7972 20544 8028
rect 20480 7968 20544 7972
rect 20560 8028 20624 8032
rect 20560 7972 20564 8028
rect 20564 7972 20620 8028
rect 20620 7972 20624 8028
rect 20560 7968 20624 7972
rect 20640 8028 20704 8032
rect 20640 7972 20644 8028
rect 20644 7972 20700 8028
rect 20700 7972 20704 8028
rect 20640 7968 20704 7972
rect 7080 7484 7144 7488
rect 7080 7428 7084 7484
rect 7084 7428 7140 7484
rect 7140 7428 7144 7484
rect 7080 7424 7144 7428
rect 7160 7484 7224 7488
rect 7160 7428 7164 7484
rect 7164 7428 7220 7484
rect 7220 7428 7224 7484
rect 7160 7424 7224 7428
rect 7240 7484 7304 7488
rect 7240 7428 7244 7484
rect 7244 7428 7300 7484
rect 7300 7428 7304 7484
rect 7240 7424 7304 7428
rect 7320 7484 7384 7488
rect 7320 7428 7324 7484
rect 7324 7428 7380 7484
rect 7380 7428 7384 7484
rect 7320 7424 7384 7428
rect 12408 7484 12472 7488
rect 12408 7428 12412 7484
rect 12412 7428 12468 7484
rect 12468 7428 12472 7484
rect 12408 7424 12472 7428
rect 12488 7484 12552 7488
rect 12488 7428 12492 7484
rect 12492 7428 12548 7484
rect 12548 7428 12552 7484
rect 12488 7424 12552 7428
rect 12568 7484 12632 7488
rect 12568 7428 12572 7484
rect 12572 7428 12628 7484
rect 12628 7428 12632 7484
rect 12568 7424 12632 7428
rect 12648 7484 12712 7488
rect 12648 7428 12652 7484
rect 12652 7428 12708 7484
rect 12708 7428 12712 7484
rect 12648 7424 12712 7428
rect 17736 7484 17800 7488
rect 17736 7428 17740 7484
rect 17740 7428 17796 7484
rect 17796 7428 17800 7484
rect 17736 7424 17800 7428
rect 17816 7484 17880 7488
rect 17816 7428 17820 7484
rect 17820 7428 17876 7484
rect 17876 7428 17880 7484
rect 17816 7424 17880 7428
rect 17896 7484 17960 7488
rect 17896 7428 17900 7484
rect 17900 7428 17956 7484
rect 17956 7428 17960 7484
rect 17896 7424 17960 7428
rect 17976 7484 18040 7488
rect 17976 7428 17980 7484
rect 17980 7428 18036 7484
rect 18036 7428 18040 7484
rect 17976 7424 18040 7428
rect 4416 6940 4480 6944
rect 4416 6884 4420 6940
rect 4420 6884 4476 6940
rect 4476 6884 4480 6940
rect 4416 6880 4480 6884
rect 4496 6940 4560 6944
rect 4496 6884 4500 6940
rect 4500 6884 4556 6940
rect 4556 6884 4560 6940
rect 4496 6880 4560 6884
rect 4576 6940 4640 6944
rect 4576 6884 4580 6940
rect 4580 6884 4636 6940
rect 4636 6884 4640 6940
rect 4576 6880 4640 6884
rect 4656 6940 4720 6944
rect 4656 6884 4660 6940
rect 4660 6884 4716 6940
rect 4716 6884 4720 6940
rect 4656 6880 4720 6884
rect 9744 6940 9808 6944
rect 9744 6884 9748 6940
rect 9748 6884 9804 6940
rect 9804 6884 9808 6940
rect 9744 6880 9808 6884
rect 9824 6940 9888 6944
rect 9824 6884 9828 6940
rect 9828 6884 9884 6940
rect 9884 6884 9888 6940
rect 9824 6880 9888 6884
rect 9904 6940 9968 6944
rect 9904 6884 9908 6940
rect 9908 6884 9964 6940
rect 9964 6884 9968 6940
rect 9904 6880 9968 6884
rect 9984 6940 10048 6944
rect 9984 6884 9988 6940
rect 9988 6884 10044 6940
rect 10044 6884 10048 6940
rect 9984 6880 10048 6884
rect 15072 6940 15136 6944
rect 15072 6884 15076 6940
rect 15076 6884 15132 6940
rect 15132 6884 15136 6940
rect 15072 6880 15136 6884
rect 15152 6940 15216 6944
rect 15152 6884 15156 6940
rect 15156 6884 15212 6940
rect 15212 6884 15216 6940
rect 15152 6880 15216 6884
rect 15232 6940 15296 6944
rect 15232 6884 15236 6940
rect 15236 6884 15292 6940
rect 15292 6884 15296 6940
rect 15232 6880 15296 6884
rect 15312 6940 15376 6944
rect 15312 6884 15316 6940
rect 15316 6884 15372 6940
rect 15372 6884 15376 6940
rect 15312 6880 15376 6884
rect 20400 6940 20464 6944
rect 20400 6884 20404 6940
rect 20404 6884 20460 6940
rect 20460 6884 20464 6940
rect 20400 6880 20464 6884
rect 20480 6940 20544 6944
rect 20480 6884 20484 6940
rect 20484 6884 20540 6940
rect 20540 6884 20544 6940
rect 20480 6880 20544 6884
rect 20560 6940 20624 6944
rect 20560 6884 20564 6940
rect 20564 6884 20620 6940
rect 20620 6884 20624 6940
rect 20560 6880 20624 6884
rect 20640 6940 20704 6944
rect 20640 6884 20644 6940
rect 20644 6884 20700 6940
rect 20700 6884 20704 6940
rect 20640 6880 20704 6884
rect 7080 6396 7144 6400
rect 7080 6340 7084 6396
rect 7084 6340 7140 6396
rect 7140 6340 7144 6396
rect 7080 6336 7144 6340
rect 7160 6396 7224 6400
rect 7160 6340 7164 6396
rect 7164 6340 7220 6396
rect 7220 6340 7224 6396
rect 7160 6336 7224 6340
rect 7240 6396 7304 6400
rect 7240 6340 7244 6396
rect 7244 6340 7300 6396
rect 7300 6340 7304 6396
rect 7240 6336 7304 6340
rect 7320 6396 7384 6400
rect 7320 6340 7324 6396
rect 7324 6340 7380 6396
rect 7380 6340 7384 6396
rect 7320 6336 7384 6340
rect 12408 6396 12472 6400
rect 12408 6340 12412 6396
rect 12412 6340 12468 6396
rect 12468 6340 12472 6396
rect 12408 6336 12472 6340
rect 12488 6396 12552 6400
rect 12488 6340 12492 6396
rect 12492 6340 12548 6396
rect 12548 6340 12552 6396
rect 12488 6336 12552 6340
rect 12568 6396 12632 6400
rect 12568 6340 12572 6396
rect 12572 6340 12628 6396
rect 12628 6340 12632 6396
rect 12568 6336 12632 6340
rect 12648 6396 12712 6400
rect 12648 6340 12652 6396
rect 12652 6340 12708 6396
rect 12708 6340 12712 6396
rect 12648 6336 12712 6340
rect 17736 6396 17800 6400
rect 17736 6340 17740 6396
rect 17740 6340 17796 6396
rect 17796 6340 17800 6396
rect 17736 6336 17800 6340
rect 17816 6396 17880 6400
rect 17816 6340 17820 6396
rect 17820 6340 17876 6396
rect 17876 6340 17880 6396
rect 17816 6336 17880 6340
rect 17896 6396 17960 6400
rect 17896 6340 17900 6396
rect 17900 6340 17956 6396
rect 17956 6340 17960 6396
rect 17896 6336 17960 6340
rect 17976 6396 18040 6400
rect 17976 6340 17980 6396
rect 17980 6340 18036 6396
rect 18036 6340 18040 6396
rect 17976 6336 18040 6340
rect 4416 5852 4480 5856
rect 4416 5796 4420 5852
rect 4420 5796 4476 5852
rect 4476 5796 4480 5852
rect 4416 5792 4480 5796
rect 4496 5852 4560 5856
rect 4496 5796 4500 5852
rect 4500 5796 4556 5852
rect 4556 5796 4560 5852
rect 4496 5792 4560 5796
rect 4576 5852 4640 5856
rect 4576 5796 4580 5852
rect 4580 5796 4636 5852
rect 4636 5796 4640 5852
rect 4576 5792 4640 5796
rect 4656 5852 4720 5856
rect 4656 5796 4660 5852
rect 4660 5796 4716 5852
rect 4716 5796 4720 5852
rect 4656 5792 4720 5796
rect 9744 5852 9808 5856
rect 9744 5796 9748 5852
rect 9748 5796 9804 5852
rect 9804 5796 9808 5852
rect 9744 5792 9808 5796
rect 9824 5852 9888 5856
rect 9824 5796 9828 5852
rect 9828 5796 9884 5852
rect 9884 5796 9888 5852
rect 9824 5792 9888 5796
rect 9904 5852 9968 5856
rect 9904 5796 9908 5852
rect 9908 5796 9964 5852
rect 9964 5796 9968 5852
rect 9904 5792 9968 5796
rect 9984 5852 10048 5856
rect 9984 5796 9988 5852
rect 9988 5796 10044 5852
rect 10044 5796 10048 5852
rect 9984 5792 10048 5796
rect 15072 5852 15136 5856
rect 15072 5796 15076 5852
rect 15076 5796 15132 5852
rect 15132 5796 15136 5852
rect 15072 5792 15136 5796
rect 15152 5852 15216 5856
rect 15152 5796 15156 5852
rect 15156 5796 15212 5852
rect 15212 5796 15216 5852
rect 15152 5792 15216 5796
rect 15232 5852 15296 5856
rect 15232 5796 15236 5852
rect 15236 5796 15292 5852
rect 15292 5796 15296 5852
rect 15232 5792 15296 5796
rect 15312 5852 15376 5856
rect 15312 5796 15316 5852
rect 15316 5796 15372 5852
rect 15372 5796 15376 5852
rect 15312 5792 15376 5796
rect 20400 5852 20464 5856
rect 20400 5796 20404 5852
rect 20404 5796 20460 5852
rect 20460 5796 20464 5852
rect 20400 5792 20464 5796
rect 20480 5852 20544 5856
rect 20480 5796 20484 5852
rect 20484 5796 20540 5852
rect 20540 5796 20544 5852
rect 20480 5792 20544 5796
rect 20560 5852 20624 5856
rect 20560 5796 20564 5852
rect 20564 5796 20620 5852
rect 20620 5796 20624 5852
rect 20560 5792 20624 5796
rect 20640 5852 20704 5856
rect 20640 5796 20644 5852
rect 20644 5796 20700 5852
rect 20700 5796 20704 5852
rect 20640 5792 20704 5796
rect 7080 5308 7144 5312
rect 7080 5252 7084 5308
rect 7084 5252 7140 5308
rect 7140 5252 7144 5308
rect 7080 5248 7144 5252
rect 7160 5308 7224 5312
rect 7160 5252 7164 5308
rect 7164 5252 7220 5308
rect 7220 5252 7224 5308
rect 7160 5248 7224 5252
rect 7240 5308 7304 5312
rect 7240 5252 7244 5308
rect 7244 5252 7300 5308
rect 7300 5252 7304 5308
rect 7240 5248 7304 5252
rect 7320 5308 7384 5312
rect 7320 5252 7324 5308
rect 7324 5252 7380 5308
rect 7380 5252 7384 5308
rect 7320 5248 7384 5252
rect 12408 5308 12472 5312
rect 12408 5252 12412 5308
rect 12412 5252 12468 5308
rect 12468 5252 12472 5308
rect 12408 5248 12472 5252
rect 12488 5308 12552 5312
rect 12488 5252 12492 5308
rect 12492 5252 12548 5308
rect 12548 5252 12552 5308
rect 12488 5248 12552 5252
rect 12568 5308 12632 5312
rect 12568 5252 12572 5308
rect 12572 5252 12628 5308
rect 12628 5252 12632 5308
rect 12568 5248 12632 5252
rect 12648 5308 12712 5312
rect 12648 5252 12652 5308
rect 12652 5252 12708 5308
rect 12708 5252 12712 5308
rect 12648 5248 12712 5252
rect 17736 5308 17800 5312
rect 17736 5252 17740 5308
rect 17740 5252 17796 5308
rect 17796 5252 17800 5308
rect 17736 5248 17800 5252
rect 17816 5308 17880 5312
rect 17816 5252 17820 5308
rect 17820 5252 17876 5308
rect 17876 5252 17880 5308
rect 17816 5248 17880 5252
rect 17896 5308 17960 5312
rect 17896 5252 17900 5308
rect 17900 5252 17956 5308
rect 17956 5252 17960 5308
rect 17896 5248 17960 5252
rect 17976 5308 18040 5312
rect 17976 5252 17980 5308
rect 17980 5252 18036 5308
rect 18036 5252 18040 5308
rect 17976 5248 18040 5252
rect 4416 4764 4480 4768
rect 4416 4708 4420 4764
rect 4420 4708 4476 4764
rect 4476 4708 4480 4764
rect 4416 4704 4480 4708
rect 4496 4764 4560 4768
rect 4496 4708 4500 4764
rect 4500 4708 4556 4764
rect 4556 4708 4560 4764
rect 4496 4704 4560 4708
rect 4576 4764 4640 4768
rect 4576 4708 4580 4764
rect 4580 4708 4636 4764
rect 4636 4708 4640 4764
rect 4576 4704 4640 4708
rect 4656 4764 4720 4768
rect 4656 4708 4660 4764
rect 4660 4708 4716 4764
rect 4716 4708 4720 4764
rect 4656 4704 4720 4708
rect 9744 4764 9808 4768
rect 9744 4708 9748 4764
rect 9748 4708 9804 4764
rect 9804 4708 9808 4764
rect 9744 4704 9808 4708
rect 9824 4764 9888 4768
rect 9824 4708 9828 4764
rect 9828 4708 9884 4764
rect 9884 4708 9888 4764
rect 9824 4704 9888 4708
rect 9904 4764 9968 4768
rect 9904 4708 9908 4764
rect 9908 4708 9964 4764
rect 9964 4708 9968 4764
rect 9904 4704 9968 4708
rect 9984 4764 10048 4768
rect 9984 4708 9988 4764
rect 9988 4708 10044 4764
rect 10044 4708 10048 4764
rect 9984 4704 10048 4708
rect 15072 4764 15136 4768
rect 15072 4708 15076 4764
rect 15076 4708 15132 4764
rect 15132 4708 15136 4764
rect 15072 4704 15136 4708
rect 15152 4764 15216 4768
rect 15152 4708 15156 4764
rect 15156 4708 15212 4764
rect 15212 4708 15216 4764
rect 15152 4704 15216 4708
rect 15232 4764 15296 4768
rect 15232 4708 15236 4764
rect 15236 4708 15292 4764
rect 15292 4708 15296 4764
rect 15232 4704 15296 4708
rect 15312 4764 15376 4768
rect 15312 4708 15316 4764
rect 15316 4708 15372 4764
rect 15372 4708 15376 4764
rect 15312 4704 15376 4708
rect 20400 4764 20464 4768
rect 20400 4708 20404 4764
rect 20404 4708 20460 4764
rect 20460 4708 20464 4764
rect 20400 4704 20464 4708
rect 20480 4764 20544 4768
rect 20480 4708 20484 4764
rect 20484 4708 20540 4764
rect 20540 4708 20544 4764
rect 20480 4704 20544 4708
rect 20560 4764 20624 4768
rect 20560 4708 20564 4764
rect 20564 4708 20620 4764
rect 20620 4708 20624 4764
rect 20560 4704 20624 4708
rect 20640 4764 20704 4768
rect 20640 4708 20644 4764
rect 20644 4708 20700 4764
rect 20700 4708 20704 4764
rect 20640 4704 20704 4708
rect 7080 4220 7144 4224
rect 7080 4164 7084 4220
rect 7084 4164 7140 4220
rect 7140 4164 7144 4220
rect 7080 4160 7144 4164
rect 7160 4220 7224 4224
rect 7160 4164 7164 4220
rect 7164 4164 7220 4220
rect 7220 4164 7224 4220
rect 7160 4160 7224 4164
rect 7240 4220 7304 4224
rect 7240 4164 7244 4220
rect 7244 4164 7300 4220
rect 7300 4164 7304 4220
rect 7240 4160 7304 4164
rect 7320 4220 7384 4224
rect 7320 4164 7324 4220
rect 7324 4164 7380 4220
rect 7380 4164 7384 4220
rect 7320 4160 7384 4164
rect 12408 4220 12472 4224
rect 12408 4164 12412 4220
rect 12412 4164 12468 4220
rect 12468 4164 12472 4220
rect 12408 4160 12472 4164
rect 12488 4220 12552 4224
rect 12488 4164 12492 4220
rect 12492 4164 12548 4220
rect 12548 4164 12552 4220
rect 12488 4160 12552 4164
rect 12568 4220 12632 4224
rect 12568 4164 12572 4220
rect 12572 4164 12628 4220
rect 12628 4164 12632 4220
rect 12568 4160 12632 4164
rect 12648 4220 12712 4224
rect 12648 4164 12652 4220
rect 12652 4164 12708 4220
rect 12708 4164 12712 4220
rect 12648 4160 12712 4164
rect 17736 4220 17800 4224
rect 17736 4164 17740 4220
rect 17740 4164 17796 4220
rect 17796 4164 17800 4220
rect 17736 4160 17800 4164
rect 17816 4220 17880 4224
rect 17816 4164 17820 4220
rect 17820 4164 17876 4220
rect 17876 4164 17880 4220
rect 17816 4160 17880 4164
rect 17896 4220 17960 4224
rect 17896 4164 17900 4220
rect 17900 4164 17956 4220
rect 17956 4164 17960 4220
rect 17896 4160 17960 4164
rect 17976 4220 18040 4224
rect 17976 4164 17980 4220
rect 17980 4164 18036 4220
rect 18036 4164 18040 4220
rect 17976 4160 18040 4164
rect 4416 3676 4480 3680
rect 4416 3620 4420 3676
rect 4420 3620 4476 3676
rect 4476 3620 4480 3676
rect 4416 3616 4480 3620
rect 4496 3676 4560 3680
rect 4496 3620 4500 3676
rect 4500 3620 4556 3676
rect 4556 3620 4560 3676
rect 4496 3616 4560 3620
rect 4576 3676 4640 3680
rect 4576 3620 4580 3676
rect 4580 3620 4636 3676
rect 4636 3620 4640 3676
rect 4576 3616 4640 3620
rect 4656 3676 4720 3680
rect 4656 3620 4660 3676
rect 4660 3620 4716 3676
rect 4716 3620 4720 3676
rect 4656 3616 4720 3620
rect 9744 3676 9808 3680
rect 9744 3620 9748 3676
rect 9748 3620 9804 3676
rect 9804 3620 9808 3676
rect 9744 3616 9808 3620
rect 9824 3676 9888 3680
rect 9824 3620 9828 3676
rect 9828 3620 9884 3676
rect 9884 3620 9888 3676
rect 9824 3616 9888 3620
rect 9904 3676 9968 3680
rect 9904 3620 9908 3676
rect 9908 3620 9964 3676
rect 9964 3620 9968 3676
rect 9904 3616 9968 3620
rect 9984 3676 10048 3680
rect 9984 3620 9988 3676
rect 9988 3620 10044 3676
rect 10044 3620 10048 3676
rect 9984 3616 10048 3620
rect 15072 3676 15136 3680
rect 15072 3620 15076 3676
rect 15076 3620 15132 3676
rect 15132 3620 15136 3676
rect 15072 3616 15136 3620
rect 15152 3676 15216 3680
rect 15152 3620 15156 3676
rect 15156 3620 15212 3676
rect 15212 3620 15216 3676
rect 15152 3616 15216 3620
rect 15232 3676 15296 3680
rect 15232 3620 15236 3676
rect 15236 3620 15292 3676
rect 15292 3620 15296 3676
rect 15232 3616 15296 3620
rect 15312 3676 15376 3680
rect 15312 3620 15316 3676
rect 15316 3620 15372 3676
rect 15372 3620 15376 3676
rect 15312 3616 15376 3620
rect 20400 3676 20464 3680
rect 20400 3620 20404 3676
rect 20404 3620 20460 3676
rect 20460 3620 20464 3676
rect 20400 3616 20464 3620
rect 20480 3676 20544 3680
rect 20480 3620 20484 3676
rect 20484 3620 20540 3676
rect 20540 3620 20544 3676
rect 20480 3616 20544 3620
rect 20560 3676 20624 3680
rect 20560 3620 20564 3676
rect 20564 3620 20620 3676
rect 20620 3620 20624 3676
rect 20560 3616 20624 3620
rect 20640 3676 20704 3680
rect 20640 3620 20644 3676
rect 20644 3620 20700 3676
rect 20700 3620 20704 3676
rect 20640 3616 20704 3620
rect 7080 3132 7144 3136
rect 7080 3076 7084 3132
rect 7084 3076 7140 3132
rect 7140 3076 7144 3132
rect 7080 3072 7144 3076
rect 7160 3132 7224 3136
rect 7160 3076 7164 3132
rect 7164 3076 7220 3132
rect 7220 3076 7224 3132
rect 7160 3072 7224 3076
rect 7240 3132 7304 3136
rect 7240 3076 7244 3132
rect 7244 3076 7300 3132
rect 7300 3076 7304 3132
rect 7240 3072 7304 3076
rect 7320 3132 7384 3136
rect 7320 3076 7324 3132
rect 7324 3076 7380 3132
rect 7380 3076 7384 3132
rect 7320 3072 7384 3076
rect 12408 3132 12472 3136
rect 12408 3076 12412 3132
rect 12412 3076 12468 3132
rect 12468 3076 12472 3132
rect 12408 3072 12472 3076
rect 12488 3132 12552 3136
rect 12488 3076 12492 3132
rect 12492 3076 12548 3132
rect 12548 3076 12552 3132
rect 12488 3072 12552 3076
rect 12568 3132 12632 3136
rect 12568 3076 12572 3132
rect 12572 3076 12628 3132
rect 12628 3076 12632 3132
rect 12568 3072 12632 3076
rect 12648 3132 12712 3136
rect 12648 3076 12652 3132
rect 12652 3076 12708 3132
rect 12708 3076 12712 3132
rect 12648 3072 12712 3076
rect 17736 3132 17800 3136
rect 17736 3076 17740 3132
rect 17740 3076 17796 3132
rect 17796 3076 17800 3132
rect 17736 3072 17800 3076
rect 17816 3132 17880 3136
rect 17816 3076 17820 3132
rect 17820 3076 17876 3132
rect 17876 3076 17880 3132
rect 17816 3072 17880 3076
rect 17896 3132 17960 3136
rect 17896 3076 17900 3132
rect 17900 3076 17956 3132
rect 17956 3076 17960 3132
rect 17896 3072 17960 3076
rect 17976 3132 18040 3136
rect 17976 3076 17980 3132
rect 17980 3076 18036 3132
rect 18036 3076 18040 3132
rect 17976 3072 18040 3076
rect 4416 2588 4480 2592
rect 4416 2532 4420 2588
rect 4420 2532 4476 2588
rect 4476 2532 4480 2588
rect 4416 2528 4480 2532
rect 4496 2588 4560 2592
rect 4496 2532 4500 2588
rect 4500 2532 4556 2588
rect 4556 2532 4560 2588
rect 4496 2528 4560 2532
rect 4576 2588 4640 2592
rect 4576 2532 4580 2588
rect 4580 2532 4636 2588
rect 4636 2532 4640 2588
rect 4576 2528 4640 2532
rect 4656 2588 4720 2592
rect 4656 2532 4660 2588
rect 4660 2532 4716 2588
rect 4716 2532 4720 2588
rect 4656 2528 4720 2532
rect 9744 2588 9808 2592
rect 9744 2532 9748 2588
rect 9748 2532 9804 2588
rect 9804 2532 9808 2588
rect 9744 2528 9808 2532
rect 9824 2588 9888 2592
rect 9824 2532 9828 2588
rect 9828 2532 9884 2588
rect 9884 2532 9888 2588
rect 9824 2528 9888 2532
rect 9904 2588 9968 2592
rect 9904 2532 9908 2588
rect 9908 2532 9964 2588
rect 9964 2532 9968 2588
rect 9904 2528 9968 2532
rect 9984 2588 10048 2592
rect 9984 2532 9988 2588
rect 9988 2532 10044 2588
rect 10044 2532 10048 2588
rect 9984 2528 10048 2532
rect 15072 2588 15136 2592
rect 15072 2532 15076 2588
rect 15076 2532 15132 2588
rect 15132 2532 15136 2588
rect 15072 2528 15136 2532
rect 15152 2588 15216 2592
rect 15152 2532 15156 2588
rect 15156 2532 15212 2588
rect 15212 2532 15216 2588
rect 15152 2528 15216 2532
rect 15232 2588 15296 2592
rect 15232 2532 15236 2588
rect 15236 2532 15292 2588
rect 15292 2532 15296 2588
rect 15232 2528 15296 2532
rect 15312 2588 15376 2592
rect 15312 2532 15316 2588
rect 15316 2532 15372 2588
rect 15372 2532 15376 2588
rect 15312 2528 15376 2532
rect 20400 2588 20464 2592
rect 20400 2532 20404 2588
rect 20404 2532 20460 2588
rect 20460 2532 20464 2588
rect 20400 2528 20464 2532
rect 20480 2588 20544 2592
rect 20480 2532 20484 2588
rect 20484 2532 20540 2588
rect 20540 2532 20544 2588
rect 20480 2528 20544 2532
rect 20560 2588 20624 2592
rect 20560 2532 20564 2588
rect 20564 2532 20620 2588
rect 20620 2532 20624 2588
rect 20560 2528 20624 2532
rect 20640 2588 20704 2592
rect 20640 2532 20644 2588
rect 20644 2532 20700 2588
rect 20700 2532 20704 2588
rect 20640 2528 20704 2532
rect 7080 2044 7144 2048
rect 7080 1988 7084 2044
rect 7084 1988 7140 2044
rect 7140 1988 7144 2044
rect 7080 1984 7144 1988
rect 7160 2044 7224 2048
rect 7160 1988 7164 2044
rect 7164 1988 7220 2044
rect 7220 1988 7224 2044
rect 7160 1984 7224 1988
rect 7240 2044 7304 2048
rect 7240 1988 7244 2044
rect 7244 1988 7300 2044
rect 7300 1988 7304 2044
rect 7240 1984 7304 1988
rect 7320 2044 7384 2048
rect 7320 1988 7324 2044
rect 7324 1988 7380 2044
rect 7380 1988 7384 2044
rect 7320 1984 7384 1988
rect 12408 2044 12472 2048
rect 12408 1988 12412 2044
rect 12412 1988 12468 2044
rect 12468 1988 12472 2044
rect 12408 1984 12472 1988
rect 12488 2044 12552 2048
rect 12488 1988 12492 2044
rect 12492 1988 12548 2044
rect 12548 1988 12552 2044
rect 12488 1984 12552 1988
rect 12568 2044 12632 2048
rect 12568 1988 12572 2044
rect 12572 1988 12628 2044
rect 12628 1988 12632 2044
rect 12568 1984 12632 1988
rect 12648 2044 12712 2048
rect 12648 1988 12652 2044
rect 12652 1988 12708 2044
rect 12708 1988 12712 2044
rect 12648 1984 12712 1988
rect 17736 2044 17800 2048
rect 17736 1988 17740 2044
rect 17740 1988 17796 2044
rect 17796 1988 17800 2044
rect 17736 1984 17800 1988
rect 17816 2044 17880 2048
rect 17816 1988 17820 2044
rect 17820 1988 17876 2044
rect 17876 1988 17880 2044
rect 17816 1984 17880 1988
rect 17896 2044 17960 2048
rect 17896 1988 17900 2044
rect 17900 1988 17956 2044
rect 17956 1988 17960 2044
rect 17896 1984 17960 1988
rect 17976 2044 18040 2048
rect 17976 1988 17980 2044
rect 17980 1988 18036 2044
rect 18036 1988 18040 2044
rect 17976 1984 18040 1988
rect 4416 1500 4480 1504
rect 4416 1444 4420 1500
rect 4420 1444 4476 1500
rect 4476 1444 4480 1500
rect 4416 1440 4480 1444
rect 4496 1500 4560 1504
rect 4496 1444 4500 1500
rect 4500 1444 4556 1500
rect 4556 1444 4560 1500
rect 4496 1440 4560 1444
rect 4576 1500 4640 1504
rect 4576 1444 4580 1500
rect 4580 1444 4636 1500
rect 4636 1444 4640 1500
rect 4576 1440 4640 1444
rect 4656 1500 4720 1504
rect 4656 1444 4660 1500
rect 4660 1444 4716 1500
rect 4716 1444 4720 1500
rect 4656 1440 4720 1444
rect 9744 1500 9808 1504
rect 9744 1444 9748 1500
rect 9748 1444 9804 1500
rect 9804 1444 9808 1500
rect 9744 1440 9808 1444
rect 9824 1500 9888 1504
rect 9824 1444 9828 1500
rect 9828 1444 9884 1500
rect 9884 1444 9888 1500
rect 9824 1440 9888 1444
rect 9904 1500 9968 1504
rect 9904 1444 9908 1500
rect 9908 1444 9964 1500
rect 9964 1444 9968 1500
rect 9904 1440 9968 1444
rect 9984 1500 10048 1504
rect 9984 1444 9988 1500
rect 9988 1444 10044 1500
rect 10044 1444 10048 1500
rect 9984 1440 10048 1444
rect 15072 1500 15136 1504
rect 15072 1444 15076 1500
rect 15076 1444 15132 1500
rect 15132 1444 15136 1500
rect 15072 1440 15136 1444
rect 15152 1500 15216 1504
rect 15152 1444 15156 1500
rect 15156 1444 15212 1500
rect 15212 1444 15216 1500
rect 15152 1440 15216 1444
rect 15232 1500 15296 1504
rect 15232 1444 15236 1500
rect 15236 1444 15292 1500
rect 15292 1444 15296 1500
rect 15232 1440 15296 1444
rect 15312 1500 15376 1504
rect 15312 1444 15316 1500
rect 15316 1444 15372 1500
rect 15372 1444 15376 1500
rect 15312 1440 15376 1444
rect 20400 1500 20464 1504
rect 20400 1444 20404 1500
rect 20404 1444 20460 1500
rect 20460 1444 20464 1500
rect 20400 1440 20464 1444
rect 20480 1500 20544 1504
rect 20480 1444 20484 1500
rect 20484 1444 20540 1500
rect 20540 1444 20544 1500
rect 20480 1440 20544 1444
rect 20560 1500 20624 1504
rect 20560 1444 20564 1500
rect 20564 1444 20620 1500
rect 20620 1444 20624 1500
rect 20560 1440 20624 1444
rect 20640 1500 20704 1504
rect 20640 1444 20644 1500
rect 20644 1444 20700 1500
rect 20700 1444 20704 1500
rect 20640 1440 20704 1444
rect 7080 956 7144 960
rect 7080 900 7084 956
rect 7084 900 7140 956
rect 7140 900 7144 956
rect 7080 896 7144 900
rect 7160 956 7224 960
rect 7160 900 7164 956
rect 7164 900 7220 956
rect 7220 900 7224 956
rect 7160 896 7224 900
rect 7240 956 7304 960
rect 7240 900 7244 956
rect 7244 900 7300 956
rect 7300 900 7304 956
rect 7240 896 7304 900
rect 7320 956 7384 960
rect 7320 900 7324 956
rect 7324 900 7380 956
rect 7380 900 7384 956
rect 7320 896 7384 900
rect 12408 956 12472 960
rect 12408 900 12412 956
rect 12412 900 12468 956
rect 12468 900 12472 956
rect 12408 896 12472 900
rect 12488 956 12552 960
rect 12488 900 12492 956
rect 12492 900 12548 956
rect 12548 900 12552 956
rect 12488 896 12552 900
rect 12568 956 12632 960
rect 12568 900 12572 956
rect 12572 900 12628 956
rect 12628 900 12632 956
rect 12568 896 12632 900
rect 12648 956 12712 960
rect 12648 900 12652 956
rect 12652 900 12708 956
rect 12708 900 12712 956
rect 12648 896 12712 900
rect 17736 956 17800 960
rect 17736 900 17740 956
rect 17740 900 17796 956
rect 17796 900 17800 956
rect 17736 896 17800 900
rect 17816 956 17880 960
rect 17816 900 17820 956
rect 17820 900 17876 956
rect 17876 900 17880 956
rect 17816 896 17880 900
rect 17896 956 17960 960
rect 17896 900 17900 956
rect 17900 900 17956 956
rect 17956 900 17960 956
rect 17896 896 17960 900
rect 17976 956 18040 960
rect 17976 900 17980 956
rect 17980 900 18036 956
rect 18036 900 18040 956
rect 17976 896 18040 900
<< metal4 >>
rect 4408 22176 4728 22192
rect 4408 22112 4416 22176
rect 4480 22112 4496 22176
rect 4560 22112 4576 22176
rect 4640 22112 4656 22176
rect 4720 22112 4728 22176
rect 4408 21088 4728 22112
rect 4408 21024 4416 21088
rect 4480 21024 4496 21088
rect 4560 21024 4576 21088
rect 4640 21024 4656 21088
rect 4720 21024 4728 21088
rect 4408 20838 4728 21024
rect 4408 20602 4450 20838
rect 4686 20602 4728 20838
rect 4408 20000 4728 20602
rect 4408 19936 4416 20000
rect 4480 19936 4496 20000
rect 4560 19936 4576 20000
rect 4640 19936 4656 20000
rect 4720 19936 4728 20000
rect 4408 18912 4728 19936
rect 4408 18848 4416 18912
rect 4480 18848 4496 18912
rect 4560 18848 4576 18912
rect 4640 18848 4656 18912
rect 4720 18848 4728 18912
rect 4408 17824 4728 18848
rect 4408 17760 4416 17824
rect 4480 17760 4496 17824
rect 4560 17760 4576 17824
rect 4640 17760 4656 17824
rect 4720 17760 4728 17824
rect 4408 16736 4728 17760
rect 4408 16672 4416 16736
rect 4480 16672 4496 16736
rect 4560 16672 4576 16736
rect 4640 16672 4656 16736
rect 4720 16672 4728 16736
rect 4408 15648 4728 16672
rect 4408 15584 4416 15648
rect 4480 15584 4496 15648
rect 4560 15584 4576 15648
rect 4640 15584 4656 15648
rect 4720 15584 4728 15648
rect 4408 14560 4728 15584
rect 4408 14496 4416 14560
rect 4480 14496 4496 14560
rect 4560 14496 4576 14560
rect 4640 14496 4656 14560
rect 4720 14496 4728 14560
rect 4408 13472 4728 14496
rect 4408 13408 4416 13472
rect 4480 13408 4496 13472
rect 4560 13408 4576 13472
rect 4640 13408 4656 13472
rect 4720 13408 4728 13472
rect 4408 12384 4728 13408
rect 4408 12320 4416 12384
rect 4480 12320 4496 12384
rect 4560 12320 4576 12384
rect 4640 12320 4656 12384
rect 4720 12320 4728 12384
rect 4408 11296 4728 12320
rect 4408 11232 4416 11296
rect 4480 11232 4496 11296
rect 4560 11232 4576 11296
rect 4640 11232 4656 11296
rect 4720 11232 4728 11296
rect 4408 10208 4728 11232
rect 4408 10144 4416 10208
rect 4480 10144 4496 10208
rect 4560 10144 4576 10208
rect 4640 10144 4656 10208
rect 4720 10144 4728 10208
rect 4408 9120 4728 10144
rect 4408 9056 4416 9120
rect 4480 9056 4496 9120
rect 4560 9056 4576 9120
rect 4640 9056 4656 9120
rect 4720 9056 4728 9120
rect 4408 8032 4728 9056
rect 4408 7968 4416 8032
rect 4480 7968 4496 8032
rect 4560 7968 4576 8032
rect 4640 7968 4656 8032
rect 4720 7968 4728 8032
rect 4408 6944 4728 7968
rect 4408 6880 4416 6944
rect 4480 6880 4496 6944
rect 4560 6880 4576 6944
rect 4640 6880 4656 6944
rect 4720 6880 4728 6944
rect 4408 5856 4728 6880
rect 4408 5792 4416 5856
rect 4480 5792 4496 5856
rect 4560 5792 4576 5856
rect 4640 5792 4656 5856
rect 4720 5792 4728 5856
rect 4408 4768 4728 5792
rect 4408 4704 4416 4768
rect 4480 4704 4496 4768
rect 4560 4704 4576 4768
rect 4640 4704 4656 4768
rect 4720 4704 4728 4768
rect 4408 3680 4728 4704
rect 4408 3616 4416 3680
rect 4480 3616 4496 3680
rect 4560 3616 4576 3680
rect 4640 3616 4656 3680
rect 4720 3616 4728 3680
rect 4408 2592 4728 3616
rect 4408 2528 4416 2592
rect 4480 2528 4496 2592
rect 4560 2528 4576 2592
rect 4640 2528 4656 2592
rect 4720 2528 4728 2592
rect 4408 1504 4728 2528
rect 4408 1440 4416 1504
rect 4480 1440 4496 1504
rect 4560 1440 4576 1504
rect 4640 1440 4656 1504
rect 4720 1440 4728 1504
rect 4408 880 4728 1440
rect 7072 21632 7392 22192
rect 7072 21568 7080 21632
rect 7144 21568 7160 21632
rect 7224 21568 7240 21632
rect 7304 21568 7320 21632
rect 7384 21568 7392 21632
rect 7072 20544 7392 21568
rect 7072 20480 7080 20544
rect 7144 20480 7160 20544
rect 7224 20480 7240 20544
rect 7304 20480 7320 20544
rect 7384 20480 7392 20544
rect 7072 19456 7392 20480
rect 7072 19392 7080 19456
rect 7144 19392 7160 19456
rect 7224 19392 7240 19456
rect 7304 19392 7320 19456
rect 7384 19392 7392 19456
rect 7072 18368 7392 19392
rect 7072 18304 7080 18368
rect 7144 18304 7160 18368
rect 7224 18304 7240 18368
rect 7304 18304 7320 18368
rect 7384 18304 7392 18368
rect 7072 17280 7392 18304
rect 7072 17216 7080 17280
rect 7144 17216 7160 17280
rect 7224 17216 7240 17280
rect 7304 17216 7320 17280
rect 7384 17216 7392 17280
rect 7072 16192 7392 17216
rect 7072 16128 7080 16192
rect 7144 16128 7160 16192
rect 7224 16128 7240 16192
rect 7304 16128 7320 16192
rect 7384 16128 7392 16192
rect 7072 15104 7392 16128
rect 7072 15040 7080 15104
rect 7144 15040 7160 15104
rect 7224 15040 7240 15104
rect 7304 15040 7320 15104
rect 7384 15040 7392 15104
rect 7072 14016 7392 15040
rect 7072 13952 7080 14016
rect 7144 13952 7160 14016
rect 7224 13952 7240 14016
rect 7304 13952 7320 14016
rect 7384 13952 7392 14016
rect 7072 12928 7392 13952
rect 7072 12864 7080 12928
rect 7144 12864 7160 12928
rect 7224 12864 7240 12928
rect 7304 12864 7320 12928
rect 7384 12864 7392 12928
rect 7072 11840 7392 12864
rect 7072 11776 7080 11840
rect 7144 11776 7160 11840
rect 7224 11776 7240 11840
rect 7304 11776 7320 11840
rect 7384 11776 7392 11840
rect 7072 10752 7392 11776
rect 7072 10688 7080 10752
rect 7144 10688 7160 10752
rect 7224 10688 7240 10752
rect 7304 10688 7320 10752
rect 7384 10688 7392 10752
rect 7072 9664 7392 10688
rect 7072 9600 7080 9664
rect 7144 9600 7160 9664
rect 7224 9600 7240 9664
rect 7304 9600 7320 9664
rect 7384 9600 7392 9664
rect 7072 8576 7392 9600
rect 7072 8512 7080 8576
rect 7144 8512 7160 8576
rect 7224 8512 7240 8576
rect 7304 8512 7320 8576
rect 7384 8512 7392 8576
rect 7072 7488 7392 8512
rect 7072 7424 7080 7488
rect 7144 7424 7160 7488
rect 7224 7424 7240 7488
rect 7304 7424 7320 7488
rect 7384 7424 7392 7488
rect 7072 6400 7392 7424
rect 7072 6336 7080 6400
rect 7144 6336 7160 6400
rect 7224 6336 7240 6400
rect 7304 6336 7320 6400
rect 7384 6336 7392 6400
rect 7072 5312 7392 6336
rect 7072 5248 7080 5312
rect 7144 5248 7160 5312
rect 7224 5248 7240 5312
rect 7304 5248 7320 5312
rect 7384 5248 7392 5312
rect 7072 4224 7392 5248
rect 7072 4160 7080 4224
rect 7144 4160 7160 4224
rect 7224 4160 7240 4224
rect 7304 4160 7320 4224
rect 7384 4160 7392 4224
rect 7072 3136 7392 4160
rect 7072 3072 7080 3136
rect 7144 3072 7160 3136
rect 7224 3072 7240 3136
rect 7304 3072 7320 3136
rect 7384 3072 7392 3136
rect 7072 2838 7392 3072
rect 7072 2602 7114 2838
rect 7350 2602 7392 2838
rect 7072 2048 7392 2602
rect 7072 1984 7080 2048
rect 7144 1984 7160 2048
rect 7224 1984 7240 2048
rect 7304 1984 7320 2048
rect 7384 1984 7392 2048
rect 7072 960 7392 1984
rect 7072 896 7080 960
rect 7144 896 7160 960
rect 7224 896 7240 960
rect 7304 896 7320 960
rect 7384 896 7392 960
rect 7072 880 7392 896
rect 9736 22176 10056 22192
rect 9736 22112 9744 22176
rect 9808 22112 9824 22176
rect 9888 22112 9904 22176
rect 9968 22112 9984 22176
rect 10048 22112 10056 22176
rect 9736 21088 10056 22112
rect 9736 21024 9744 21088
rect 9808 21024 9824 21088
rect 9888 21024 9904 21088
rect 9968 21024 9984 21088
rect 10048 21024 10056 21088
rect 9736 20838 10056 21024
rect 9736 20602 9778 20838
rect 10014 20602 10056 20838
rect 9736 20000 10056 20602
rect 9736 19936 9744 20000
rect 9808 19936 9824 20000
rect 9888 19936 9904 20000
rect 9968 19936 9984 20000
rect 10048 19936 10056 20000
rect 9736 18912 10056 19936
rect 9736 18848 9744 18912
rect 9808 18848 9824 18912
rect 9888 18848 9904 18912
rect 9968 18848 9984 18912
rect 10048 18848 10056 18912
rect 9736 17824 10056 18848
rect 9736 17760 9744 17824
rect 9808 17760 9824 17824
rect 9888 17760 9904 17824
rect 9968 17760 9984 17824
rect 10048 17760 10056 17824
rect 9736 16736 10056 17760
rect 9736 16672 9744 16736
rect 9808 16672 9824 16736
rect 9888 16672 9904 16736
rect 9968 16672 9984 16736
rect 10048 16672 10056 16736
rect 9736 15648 10056 16672
rect 9736 15584 9744 15648
rect 9808 15584 9824 15648
rect 9888 15584 9904 15648
rect 9968 15584 9984 15648
rect 10048 15584 10056 15648
rect 9736 14560 10056 15584
rect 9736 14496 9744 14560
rect 9808 14496 9824 14560
rect 9888 14496 9904 14560
rect 9968 14496 9984 14560
rect 10048 14496 10056 14560
rect 9736 13472 10056 14496
rect 9736 13408 9744 13472
rect 9808 13408 9824 13472
rect 9888 13408 9904 13472
rect 9968 13408 9984 13472
rect 10048 13408 10056 13472
rect 9736 12384 10056 13408
rect 9736 12320 9744 12384
rect 9808 12320 9824 12384
rect 9888 12320 9904 12384
rect 9968 12320 9984 12384
rect 10048 12320 10056 12384
rect 9736 11296 10056 12320
rect 9736 11232 9744 11296
rect 9808 11232 9824 11296
rect 9888 11232 9904 11296
rect 9968 11232 9984 11296
rect 10048 11232 10056 11296
rect 9736 10208 10056 11232
rect 9736 10144 9744 10208
rect 9808 10144 9824 10208
rect 9888 10144 9904 10208
rect 9968 10144 9984 10208
rect 10048 10144 10056 10208
rect 9736 9120 10056 10144
rect 9736 9056 9744 9120
rect 9808 9056 9824 9120
rect 9888 9056 9904 9120
rect 9968 9056 9984 9120
rect 10048 9056 10056 9120
rect 9736 8032 10056 9056
rect 9736 7968 9744 8032
rect 9808 7968 9824 8032
rect 9888 7968 9904 8032
rect 9968 7968 9984 8032
rect 10048 7968 10056 8032
rect 9736 6944 10056 7968
rect 9736 6880 9744 6944
rect 9808 6880 9824 6944
rect 9888 6880 9904 6944
rect 9968 6880 9984 6944
rect 10048 6880 10056 6944
rect 9736 5856 10056 6880
rect 9736 5792 9744 5856
rect 9808 5792 9824 5856
rect 9888 5792 9904 5856
rect 9968 5792 9984 5856
rect 10048 5792 10056 5856
rect 9736 4768 10056 5792
rect 9736 4704 9744 4768
rect 9808 4704 9824 4768
rect 9888 4704 9904 4768
rect 9968 4704 9984 4768
rect 10048 4704 10056 4768
rect 9736 3680 10056 4704
rect 9736 3616 9744 3680
rect 9808 3616 9824 3680
rect 9888 3616 9904 3680
rect 9968 3616 9984 3680
rect 10048 3616 10056 3680
rect 9736 2592 10056 3616
rect 9736 2528 9744 2592
rect 9808 2528 9824 2592
rect 9888 2528 9904 2592
rect 9968 2528 9984 2592
rect 10048 2528 10056 2592
rect 9736 1504 10056 2528
rect 9736 1440 9744 1504
rect 9808 1440 9824 1504
rect 9888 1440 9904 1504
rect 9968 1440 9984 1504
rect 10048 1440 10056 1504
rect 9736 880 10056 1440
rect 12400 21632 12720 22192
rect 12400 21568 12408 21632
rect 12472 21568 12488 21632
rect 12552 21568 12568 21632
rect 12632 21568 12648 21632
rect 12712 21568 12720 21632
rect 12400 20544 12720 21568
rect 12400 20480 12408 20544
rect 12472 20480 12488 20544
rect 12552 20480 12568 20544
rect 12632 20480 12648 20544
rect 12712 20480 12720 20544
rect 12400 19456 12720 20480
rect 12400 19392 12408 19456
rect 12472 19392 12488 19456
rect 12552 19392 12568 19456
rect 12632 19392 12648 19456
rect 12712 19392 12720 19456
rect 12400 18368 12720 19392
rect 12400 18304 12408 18368
rect 12472 18304 12488 18368
rect 12552 18304 12568 18368
rect 12632 18304 12648 18368
rect 12712 18304 12720 18368
rect 12400 17280 12720 18304
rect 12400 17216 12408 17280
rect 12472 17216 12488 17280
rect 12552 17216 12568 17280
rect 12632 17216 12648 17280
rect 12712 17216 12720 17280
rect 12400 16192 12720 17216
rect 12400 16128 12408 16192
rect 12472 16128 12488 16192
rect 12552 16128 12568 16192
rect 12632 16128 12648 16192
rect 12712 16128 12720 16192
rect 12400 15104 12720 16128
rect 12400 15040 12408 15104
rect 12472 15040 12488 15104
rect 12552 15040 12568 15104
rect 12632 15040 12648 15104
rect 12712 15040 12720 15104
rect 12400 14016 12720 15040
rect 12400 13952 12408 14016
rect 12472 13952 12488 14016
rect 12552 13952 12568 14016
rect 12632 13952 12648 14016
rect 12712 13952 12720 14016
rect 12400 12928 12720 13952
rect 12400 12864 12408 12928
rect 12472 12864 12488 12928
rect 12552 12864 12568 12928
rect 12632 12864 12648 12928
rect 12712 12864 12720 12928
rect 12400 11840 12720 12864
rect 12400 11776 12408 11840
rect 12472 11776 12488 11840
rect 12552 11776 12568 11840
rect 12632 11776 12648 11840
rect 12712 11776 12720 11840
rect 12400 10752 12720 11776
rect 12400 10688 12408 10752
rect 12472 10688 12488 10752
rect 12552 10688 12568 10752
rect 12632 10688 12648 10752
rect 12712 10688 12720 10752
rect 12400 9664 12720 10688
rect 12400 9600 12408 9664
rect 12472 9600 12488 9664
rect 12552 9600 12568 9664
rect 12632 9600 12648 9664
rect 12712 9600 12720 9664
rect 12400 8576 12720 9600
rect 12400 8512 12408 8576
rect 12472 8512 12488 8576
rect 12552 8512 12568 8576
rect 12632 8512 12648 8576
rect 12712 8512 12720 8576
rect 12400 7488 12720 8512
rect 12400 7424 12408 7488
rect 12472 7424 12488 7488
rect 12552 7424 12568 7488
rect 12632 7424 12648 7488
rect 12712 7424 12720 7488
rect 12400 6400 12720 7424
rect 12400 6336 12408 6400
rect 12472 6336 12488 6400
rect 12552 6336 12568 6400
rect 12632 6336 12648 6400
rect 12712 6336 12720 6400
rect 12400 5312 12720 6336
rect 12400 5248 12408 5312
rect 12472 5248 12488 5312
rect 12552 5248 12568 5312
rect 12632 5248 12648 5312
rect 12712 5248 12720 5312
rect 12400 4224 12720 5248
rect 12400 4160 12408 4224
rect 12472 4160 12488 4224
rect 12552 4160 12568 4224
rect 12632 4160 12648 4224
rect 12712 4160 12720 4224
rect 12400 3136 12720 4160
rect 12400 3072 12408 3136
rect 12472 3072 12488 3136
rect 12552 3072 12568 3136
rect 12632 3072 12648 3136
rect 12712 3072 12720 3136
rect 12400 2838 12720 3072
rect 12400 2602 12442 2838
rect 12678 2602 12720 2838
rect 12400 2048 12720 2602
rect 12400 1984 12408 2048
rect 12472 1984 12488 2048
rect 12552 1984 12568 2048
rect 12632 1984 12648 2048
rect 12712 1984 12720 2048
rect 12400 960 12720 1984
rect 12400 896 12408 960
rect 12472 896 12488 960
rect 12552 896 12568 960
rect 12632 896 12648 960
rect 12712 896 12720 960
rect 12400 880 12720 896
rect 15064 22176 15384 22192
rect 15064 22112 15072 22176
rect 15136 22112 15152 22176
rect 15216 22112 15232 22176
rect 15296 22112 15312 22176
rect 15376 22112 15384 22176
rect 15064 21088 15384 22112
rect 15064 21024 15072 21088
rect 15136 21024 15152 21088
rect 15216 21024 15232 21088
rect 15296 21024 15312 21088
rect 15376 21024 15384 21088
rect 15064 20838 15384 21024
rect 15064 20602 15106 20838
rect 15342 20602 15384 20838
rect 15064 20000 15384 20602
rect 15064 19936 15072 20000
rect 15136 19936 15152 20000
rect 15216 19936 15232 20000
rect 15296 19936 15312 20000
rect 15376 19936 15384 20000
rect 15064 18912 15384 19936
rect 15064 18848 15072 18912
rect 15136 18848 15152 18912
rect 15216 18848 15232 18912
rect 15296 18848 15312 18912
rect 15376 18848 15384 18912
rect 15064 17824 15384 18848
rect 15064 17760 15072 17824
rect 15136 17760 15152 17824
rect 15216 17760 15232 17824
rect 15296 17760 15312 17824
rect 15376 17760 15384 17824
rect 15064 16736 15384 17760
rect 15064 16672 15072 16736
rect 15136 16672 15152 16736
rect 15216 16672 15232 16736
rect 15296 16672 15312 16736
rect 15376 16672 15384 16736
rect 15064 15648 15384 16672
rect 15064 15584 15072 15648
rect 15136 15584 15152 15648
rect 15216 15584 15232 15648
rect 15296 15584 15312 15648
rect 15376 15584 15384 15648
rect 15064 14560 15384 15584
rect 15064 14496 15072 14560
rect 15136 14496 15152 14560
rect 15216 14496 15232 14560
rect 15296 14496 15312 14560
rect 15376 14496 15384 14560
rect 15064 13472 15384 14496
rect 15064 13408 15072 13472
rect 15136 13408 15152 13472
rect 15216 13408 15232 13472
rect 15296 13408 15312 13472
rect 15376 13408 15384 13472
rect 15064 12384 15384 13408
rect 15064 12320 15072 12384
rect 15136 12320 15152 12384
rect 15216 12320 15232 12384
rect 15296 12320 15312 12384
rect 15376 12320 15384 12384
rect 15064 11296 15384 12320
rect 15064 11232 15072 11296
rect 15136 11232 15152 11296
rect 15216 11232 15232 11296
rect 15296 11232 15312 11296
rect 15376 11232 15384 11296
rect 15064 10208 15384 11232
rect 15064 10144 15072 10208
rect 15136 10144 15152 10208
rect 15216 10144 15232 10208
rect 15296 10144 15312 10208
rect 15376 10144 15384 10208
rect 15064 9120 15384 10144
rect 15064 9056 15072 9120
rect 15136 9056 15152 9120
rect 15216 9056 15232 9120
rect 15296 9056 15312 9120
rect 15376 9056 15384 9120
rect 15064 8032 15384 9056
rect 15064 7968 15072 8032
rect 15136 7968 15152 8032
rect 15216 7968 15232 8032
rect 15296 7968 15312 8032
rect 15376 7968 15384 8032
rect 15064 6944 15384 7968
rect 15064 6880 15072 6944
rect 15136 6880 15152 6944
rect 15216 6880 15232 6944
rect 15296 6880 15312 6944
rect 15376 6880 15384 6944
rect 15064 5856 15384 6880
rect 15064 5792 15072 5856
rect 15136 5792 15152 5856
rect 15216 5792 15232 5856
rect 15296 5792 15312 5856
rect 15376 5792 15384 5856
rect 15064 4768 15384 5792
rect 15064 4704 15072 4768
rect 15136 4704 15152 4768
rect 15216 4704 15232 4768
rect 15296 4704 15312 4768
rect 15376 4704 15384 4768
rect 15064 3680 15384 4704
rect 15064 3616 15072 3680
rect 15136 3616 15152 3680
rect 15216 3616 15232 3680
rect 15296 3616 15312 3680
rect 15376 3616 15384 3680
rect 15064 2592 15384 3616
rect 15064 2528 15072 2592
rect 15136 2528 15152 2592
rect 15216 2528 15232 2592
rect 15296 2528 15312 2592
rect 15376 2528 15384 2592
rect 15064 1504 15384 2528
rect 15064 1440 15072 1504
rect 15136 1440 15152 1504
rect 15216 1440 15232 1504
rect 15296 1440 15312 1504
rect 15376 1440 15384 1504
rect 15064 880 15384 1440
rect 17728 21632 18048 22192
rect 17728 21568 17736 21632
rect 17800 21568 17816 21632
rect 17880 21568 17896 21632
rect 17960 21568 17976 21632
rect 18040 21568 18048 21632
rect 17728 20544 18048 21568
rect 17728 20480 17736 20544
rect 17800 20480 17816 20544
rect 17880 20480 17896 20544
rect 17960 20480 17976 20544
rect 18040 20480 18048 20544
rect 17728 19456 18048 20480
rect 17728 19392 17736 19456
rect 17800 19392 17816 19456
rect 17880 19392 17896 19456
rect 17960 19392 17976 19456
rect 18040 19392 18048 19456
rect 17728 18368 18048 19392
rect 17728 18304 17736 18368
rect 17800 18304 17816 18368
rect 17880 18304 17896 18368
rect 17960 18304 17976 18368
rect 18040 18304 18048 18368
rect 17728 17280 18048 18304
rect 17728 17216 17736 17280
rect 17800 17216 17816 17280
rect 17880 17216 17896 17280
rect 17960 17216 17976 17280
rect 18040 17216 18048 17280
rect 17728 16192 18048 17216
rect 17728 16128 17736 16192
rect 17800 16128 17816 16192
rect 17880 16128 17896 16192
rect 17960 16128 17976 16192
rect 18040 16128 18048 16192
rect 17728 15104 18048 16128
rect 17728 15040 17736 15104
rect 17800 15040 17816 15104
rect 17880 15040 17896 15104
rect 17960 15040 17976 15104
rect 18040 15040 18048 15104
rect 17728 14016 18048 15040
rect 17728 13952 17736 14016
rect 17800 13952 17816 14016
rect 17880 13952 17896 14016
rect 17960 13952 17976 14016
rect 18040 13952 18048 14016
rect 17728 12928 18048 13952
rect 17728 12864 17736 12928
rect 17800 12864 17816 12928
rect 17880 12864 17896 12928
rect 17960 12864 17976 12928
rect 18040 12864 18048 12928
rect 17728 11840 18048 12864
rect 17728 11776 17736 11840
rect 17800 11776 17816 11840
rect 17880 11776 17896 11840
rect 17960 11776 17976 11840
rect 18040 11776 18048 11840
rect 17728 10752 18048 11776
rect 17728 10688 17736 10752
rect 17800 10688 17816 10752
rect 17880 10688 17896 10752
rect 17960 10688 17976 10752
rect 18040 10688 18048 10752
rect 17728 9664 18048 10688
rect 17728 9600 17736 9664
rect 17800 9600 17816 9664
rect 17880 9600 17896 9664
rect 17960 9600 17976 9664
rect 18040 9600 18048 9664
rect 17728 8576 18048 9600
rect 17728 8512 17736 8576
rect 17800 8512 17816 8576
rect 17880 8512 17896 8576
rect 17960 8512 17976 8576
rect 18040 8512 18048 8576
rect 17728 7488 18048 8512
rect 17728 7424 17736 7488
rect 17800 7424 17816 7488
rect 17880 7424 17896 7488
rect 17960 7424 17976 7488
rect 18040 7424 18048 7488
rect 17728 6400 18048 7424
rect 17728 6336 17736 6400
rect 17800 6336 17816 6400
rect 17880 6336 17896 6400
rect 17960 6336 17976 6400
rect 18040 6336 18048 6400
rect 17728 5312 18048 6336
rect 17728 5248 17736 5312
rect 17800 5248 17816 5312
rect 17880 5248 17896 5312
rect 17960 5248 17976 5312
rect 18040 5248 18048 5312
rect 17728 4224 18048 5248
rect 17728 4160 17736 4224
rect 17800 4160 17816 4224
rect 17880 4160 17896 4224
rect 17960 4160 17976 4224
rect 18040 4160 18048 4224
rect 17728 3136 18048 4160
rect 17728 3072 17736 3136
rect 17800 3072 17816 3136
rect 17880 3072 17896 3136
rect 17960 3072 17976 3136
rect 18040 3072 18048 3136
rect 17728 2838 18048 3072
rect 17728 2602 17770 2838
rect 18006 2602 18048 2838
rect 17728 2048 18048 2602
rect 17728 1984 17736 2048
rect 17800 1984 17816 2048
rect 17880 1984 17896 2048
rect 17960 1984 17976 2048
rect 18040 1984 18048 2048
rect 17728 960 18048 1984
rect 17728 896 17736 960
rect 17800 896 17816 960
rect 17880 896 17896 960
rect 17960 896 17976 960
rect 18040 896 18048 960
rect 17728 880 18048 896
rect 20392 22176 20712 22192
rect 20392 22112 20400 22176
rect 20464 22112 20480 22176
rect 20544 22112 20560 22176
rect 20624 22112 20640 22176
rect 20704 22112 20712 22176
rect 20392 21088 20712 22112
rect 20392 21024 20400 21088
rect 20464 21024 20480 21088
rect 20544 21024 20560 21088
rect 20624 21024 20640 21088
rect 20704 21024 20712 21088
rect 20392 20838 20712 21024
rect 20392 20602 20434 20838
rect 20670 20602 20712 20838
rect 20392 20000 20712 20602
rect 20392 19936 20400 20000
rect 20464 19936 20480 20000
rect 20544 19936 20560 20000
rect 20624 19936 20640 20000
rect 20704 19936 20712 20000
rect 20392 18912 20712 19936
rect 20392 18848 20400 18912
rect 20464 18848 20480 18912
rect 20544 18848 20560 18912
rect 20624 18848 20640 18912
rect 20704 18848 20712 18912
rect 20392 17824 20712 18848
rect 20392 17760 20400 17824
rect 20464 17760 20480 17824
rect 20544 17760 20560 17824
rect 20624 17760 20640 17824
rect 20704 17760 20712 17824
rect 20392 16736 20712 17760
rect 20392 16672 20400 16736
rect 20464 16672 20480 16736
rect 20544 16672 20560 16736
rect 20624 16672 20640 16736
rect 20704 16672 20712 16736
rect 20392 15648 20712 16672
rect 20392 15584 20400 15648
rect 20464 15584 20480 15648
rect 20544 15584 20560 15648
rect 20624 15584 20640 15648
rect 20704 15584 20712 15648
rect 20392 14560 20712 15584
rect 20392 14496 20400 14560
rect 20464 14496 20480 14560
rect 20544 14496 20560 14560
rect 20624 14496 20640 14560
rect 20704 14496 20712 14560
rect 20392 13472 20712 14496
rect 20392 13408 20400 13472
rect 20464 13408 20480 13472
rect 20544 13408 20560 13472
rect 20624 13408 20640 13472
rect 20704 13408 20712 13472
rect 20392 12384 20712 13408
rect 20392 12320 20400 12384
rect 20464 12320 20480 12384
rect 20544 12320 20560 12384
rect 20624 12320 20640 12384
rect 20704 12320 20712 12384
rect 20392 11296 20712 12320
rect 20392 11232 20400 11296
rect 20464 11232 20480 11296
rect 20544 11232 20560 11296
rect 20624 11232 20640 11296
rect 20704 11232 20712 11296
rect 20392 10208 20712 11232
rect 20392 10144 20400 10208
rect 20464 10144 20480 10208
rect 20544 10144 20560 10208
rect 20624 10144 20640 10208
rect 20704 10144 20712 10208
rect 20392 9120 20712 10144
rect 20392 9056 20400 9120
rect 20464 9056 20480 9120
rect 20544 9056 20560 9120
rect 20624 9056 20640 9120
rect 20704 9056 20712 9120
rect 20392 8032 20712 9056
rect 20392 7968 20400 8032
rect 20464 7968 20480 8032
rect 20544 7968 20560 8032
rect 20624 7968 20640 8032
rect 20704 7968 20712 8032
rect 20392 6944 20712 7968
rect 20392 6880 20400 6944
rect 20464 6880 20480 6944
rect 20544 6880 20560 6944
rect 20624 6880 20640 6944
rect 20704 6880 20712 6944
rect 20392 5856 20712 6880
rect 20392 5792 20400 5856
rect 20464 5792 20480 5856
rect 20544 5792 20560 5856
rect 20624 5792 20640 5856
rect 20704 5792 20712 5856
rect 20392 4768 20712 5792
rect 20392 4704 20400 4768
rect 20464 4704 20480 4768
rect 20544 4704 20560 4768
rect 20624 4704 20640 4768
rect 20704 4704 20712 4768
rect 20392 3680 20712 4704
rect 20392 3616 20400 3680
rect 20464 3616 20480 3680
rect 20544 3616 20560 3680
rect 20624 3616 20640 3680
rect 20704 3616 20712 3680
rect 20392 2592 20712 3616
rect 20392 2528 20400 2592
rect 20464 2528 20480 2592
rect 20544 2528 20560 2592
rect 20624 2528 20640 2592
rect 20704 2528 20712 2592
rect 20392 1504 20712 2528
rect 20392 1440 20400 1504
rect 20464 1440 20480 1504
rect 20544 1440 20560 1504
rect 20624 1440 20640 1504
rect 20704 1440 20712 1504
rect 20392 880 20712 1440
<< via4 >>
rect 4450 20602 4686 20838
rect 7114 2602 7350 2838
rect 9778 20602 10014 20838
rect 12442 2602 12678 2838
rect 15106 20602 15342 20838
rect 17770 2602 18006 2838
rect 20434 20602 20670 20838
<< metal5 >>
rect 1904 20838 22236 20880
rect 1904 20602 4450 20838
rect 4686 20602 9778 20838
rect 10014 20602 15106 20838
rect 15342 20602 20434 20838
rect 20670 20602 22236 20838
rect 1904 20560 22236 20602
rect 1904 2838 22236 2880
rect 1904 2602 7114 2838
rect 7350 2602 12442 2838
rect 12678 2602 17770 2838
rect 18006 2602 22236 2838
rect 1904 2560 22236 2602
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2732 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1996 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_2
timestamp 1607194113
transform 1 0 1904 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_0
timestamp 1607194113
transform 1 0 2732 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_1
timestamp 1607194113
transform 1 0 1996 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_0
timestamp 1607194113
transform 1 0 1904 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3100 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2824 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_0
timestamp 1607194113
transform 1 0 3100 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_0
timestamp 1607194113
transform 1 0 2824 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_30
timestamp 1607194113
transform 1 0 4296 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_1
timestamp 1607194113
transform 1 0 4020 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_1
timestamp 1607194113
transform 1 0 3928 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_1
timestamp 1607194113
transform 1 0 4296 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_1
timestamp 1607194113
transform 1 0 4020 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_1
timestamp 1607194113
transform 1 0 3928 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_29
timestamp 1607194113
transform 1 0 5492 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_2
timestamp 1607194113
transform 1 0 5216 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_2
timestamp 1607194113
transform 1 0 5124 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_2
timestamp 1607194113
transform 1 0 5492 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_2
timestamp 1607194113
transform 1 0 5216 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_2
timestamp 1607194113
transform 1 0 5124 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_3
timestamp 1607194113
transform 1 0 6412 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_3
timestamp 1607194113
transform 1 0 6320 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_3
timestamp 1607194113
transform 1 0 6412 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_3
timestamp 1607194113
transform 1 0 6320 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_28
timestamp 1607194113
transform 1 0 6688 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_3
timestamp 1607194113
transform 1 0 6688 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_27
timestamp 1607194113
transform 1 0 7884 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_4
timestamp 1607194113
transform 1 0 7608 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_4
timestamp 1607194113
transform 1 0 7516 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_4
timestamp 1607194113
transform 1 0 7884 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_4
timestamp 1607194113
transform 1 0 7608 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_4
timestamp 1607194113
transform 1 0 7516 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_26
timestamp 1607194113
transform 1 0 9080 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_5
timestamp 1607194113
transform 1 0 8804 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_5
timestamp 1607194113
transform 1 0 8712 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_5
timestamp 1607194113
transform 1 0 9080 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_5
timestamp 1607194113
transform 1 0 8804 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_5
timestamp 1607194113
transform 1 0 8712 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_6
timestamp 1607194113
transform 1 0 10000 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_6
timestamp 1607194113
transform 1 0 9908 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_6
timestamp 1607194113
transform 1 0 10000 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_6
timestamp 1607194113
transform 1 0 9908 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_25
timestamp 1607194113
transform 1 0 10276 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_6
timestamp 1607194113
transform 1 0 10276 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_24
timestamp 1607194113
transform 1 0 11472 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_7
timestamp 1607194113
transform 1 0 11196 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_7
timestamp 1607194113
transform 1 0 11104 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_7
timestamp 1607194113
transform 1 0 11472 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_7
timestamp 1607194113
transform 1 0 11196 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_7
timestamp 1607194113
transform 1 0 11104 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_23
timestamp 1607194113
transform 1 0 12668 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_8
timestamp 1607194113
transform 1 0 12392 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_8
timestamp 1607194113
transform 1 0 12300 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_8
timestamp 1607194113
transform 1 0 12668 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_8
timestamp 1607194113
transform 1 0 12392 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_8
timestamp 1607194113
transform 1 0 12300 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_9
timestamp 1607194113
transform 1 0 13588 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_9
timestamp 1607194113
transform 1 0 13496 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_9
timestamp 1607194113
transform 1 0 13588 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_9
timestamp 1607194113
transform 1 0 13496 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_22
timestamp 1607194113
transform 1 0 13864 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_9
timestamp 1607194113
transform 1 0 13864 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_21
timestamp 1607194113
transform 1 0 15060 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_10
timestamp 1607194113
transform 1 0 14784 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_10
timestamp 1607194113
transform 1 0 14692 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_10
timestamp 1607194113
transform 1 0 15060 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_10
timestamp 1607194113
transform 1 0 14784 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_10
timestamp 1607194113
transform 1 0 14692 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_20
timestamp 1607194113
transform 1 0 16256 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_11
timestamp 1607194113
transform 1 0 15980 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_11
timestamp 1607194113
transform 1 0 15888 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_11
timestamp 1607194113
transform 1 0 16256 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_11
timestamp 1607194113
transform 1 0 15980 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_11
timestamp 1607194113
transform 1 0 15888 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_12
timestamp 1607194113
transform 1 0 17176 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_12
timestamp 1607194113
transform 1 0 17084 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_12
timestamp 1607194113
transform 1 0 17176 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_12
timestamp 1607194113
transform 1 0 17084 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_19
timestamp 1607194113
transform 1 0 17452 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_12
timestamp 1607194113
transform 1 0 17452 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_18
timestamp 1607194113
transform 1 0 18648 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_13
timestamp 1607194113
transform 1 0 18372 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_13
timestamp 1607194113
transform 1 0 18280 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_13
timestamp 1607194113
transform 1 0 18648 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_13
timestamp 1607194113
transform 1 0 18372 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_13
timestamp 1607194113
transform 1 0 18280 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_17
timestamp 1607194113
transform 1 0 19844 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_14
timestamp 1607194113
transform 1 0 19568 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_14
timestamp 1607194113
transform 1 0 19476 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_14
timestamp 1607194113
transform 1 0 19844 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap0_14
timestamp 1607194113
transform 1 0 19568 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_14
timestamp 1607194113
transform 1 0 19476 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_15
timestamp 1607194113
transform 1 0 20764 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_15
timestamp 1607194113
transform 1 0 20672 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_15
timestamp 1607194113
transform 1 0 20764 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_15
timestamp 1607194113
transform 1 0 20672 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_16
timestamp 1607194113
transform 1 0 21040 0 1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_15
timestamp 1607194113
transform 1 0 21040 0 -1 1472
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap1_16
timestamp 1607194113
transform 1 0 21960 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_16
timestamp 1607194113
transform 1 0 21868 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_16
timestamp 1607194113
transform 1 0 21960 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_16
timestamp 1607194113
transform 1 0 21868 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_0
timestamp 1607194113
transform 1 0 2732 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_5
timestamp 1607194113
transform 1 0 1996 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_4
timestamp 1607194113
transform 1 0 1904 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_32
timestamp 1607194113
transform 1 0 3100 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_0
timestamp 1607194113
transform 1 0 2824 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_33
timestamp 1607194113
transform 1 0 4296 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_1
timestamp 1607194113
transform 1 0 4020 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_1
timestamp 1607194113
transform 1 0 3928 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_34
timestamp 1607194113
transform 1 0 5492 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_2
timestamp 1607194113
transform 1 0 5216 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_2
timestamp 1607194113
transform 1 0 5124 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_3
timestamp 1607194113
transform 1 0 6412 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_3
timestamp 1607194113
transform 1 0 6320 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_35
timestamp 1607194113
transform 1 0 6688 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_36
timestamp 1607194113
transform 1 0 7884 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_4
timestamp 1607194113
transform 1 0 7608 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_4
timestamp 1607194113
transform 1 0 7516 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_37
timestamp 1607194113
transform 1 0 9080 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_5
timestamp 1607194113
transform 1 0 8804 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_5
timestamp 1607194113
transform 1 0 8712 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_6
timestamp 1607194113
transform 1 0 10000 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_6
timestamp 1607194113
transform 1 0 9908 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_38
timestamp 1607194113
transform 1 0 10276 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_39
timestamp 1607194113
transform 1 0 11472 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_7
timestamp 1607194113
transform 1 0 11196 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_7
timestamp 1607194113
transform 1 0 11104 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_40
timestamp 1607194113
transform 1 0 12668 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_8
timestamp 1607194113
transform 1 0 12392 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_8
timestamp 1607194113
transform 1 0 12300 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_9
timestamp 1607194113
transform 1 0 13588 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_9
timestamp 1607194113
transform 1 0 13496 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_41
timestamp 1607194113
transform 1 0 13864 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_42
timestamp 1607194113
transform 1 0 15060 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_10
timestamp 1607194113
transform 1 0 14784 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_10
timestamp 1607194113
transform 1 0 14692 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_43
timestamp 1607194113
transform 1 0 16256 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_11
timestamp 1607194113
transform 1 0 15980 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_11
timestamp 1607194113
transform 1 0 15888 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_12
timestamp 1607194113
transform 1 0 17176 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_12
timestamp 1607194113
transform 1 0 17084 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_44
timestamp 1607194113
transform 1 0 17452 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_45
timestamp 1607194113
transform 1 0 18648 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_13
timestamp 1607194113
transform 1 0 18372 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_13
timestamp 1607194113
transform 1 0 18280 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_46
timestamp 1607194113
transform 1 0 19844 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_14
timestamp 1607194113
transform 1 0 19568 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_14
timestamp 1607194113
transform 1 0 19476 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_15
timestamp 1607194113
transform 1 0 20764 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_15
timestamp 1607194113
transform 1 0 20672 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_47
timestamp 1607194113
transform 1 0 21040 0 -1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap2_16
timestamp 1607194113
transform 1 0 21960 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_16
timestamp 1607194113
transform 1 0 21868 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_0
timestamp 1607194113
transform 1 0 2732 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_7
timestamp 1607194113
transform 1 0 1996 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_6
timestamp 1607194113
transform 1 0 1904 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_63
timestamp 1607194113
transform 1 0 3100 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_0
timestamp 1607194113
transform 1 0 2824 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_62
timestamp 1607194113
transform 1 0 4296 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_1
timestamp 1607194113
transform 1 0 4020 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_1
timestamp 1607194113
transform 1 0 3928 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_61
timestamp 1607194113
transform 1 0 5492 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_2
timestamp 1607194113
transform 1 0 5216 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_2
timestamp 1607194113
transform 1 0 5124 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_3
timestamp 1607194113
transform 1 0 6412 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_3
timestamp 1607194113
transform 1 0 6320 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_60
timestamp 1607194113
transform 1 0 6688 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_59
timestamp 1607194113
transform 1 0 7884 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_4
timestamp 1607194113
transform 1 0 7608 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_4
timestamp 1607194113
transform 1 0 7516 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_58
timestamp 1607194113
transform 1 0 9080 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_5
timestamp 1607194113
transform 1 0 8804 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_5
timestamp 1607194113
transform 1 0 8712 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_6
timestamp 1607194113
transform 1 0 10000 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_6
timestamp 1607194113
transform 1 0 9908 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_57
timestamp 1607194113
transform 1 0 10276 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_56
timestamp 1607194113
transform 1 0 11472 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_7
timestamp 1607194113
transform 1 0 11196 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_7
timestamp 1607194113
transform 1 0 11104 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_55
timestamp 1607194113
transform 1 0 12668 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_8
timestamp 1607194113
transform 1 0 12392 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_8
timestamp 1607194113
transform 1 0 12300 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_9
timestamp 1607194113
transform 1 0 13588 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_9
timestamp 1607194113
transform 1 0 13496 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_54
timestamp 1607194113
transform 1 0 13864 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_53
timestamp 1607194113
transform 1 0 15060 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_10
timestamp 1607194113
transform 1 0 14784 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_10
timestamp 1607194113
transform 1 0 14692 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_52
timestamp 1607194113
transform 1 0 16256 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_11
timestamp 1607194113
transform 1 0 15980 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_11
timestamp 1607194113
transform 1 0 15888 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_12
timestamp 1607194113
transform 1 0 17176 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_12
timestamp 1607194113
transform 1 0 17084 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_51
timestamp 1607194113
transform 1 0 17452 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_50
timestamp 1607194113
transform 1 0 18648 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_13
timestamp 1607194113
transform 1 0 18372 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_13
timestamp 1607194113
transform 1 0 18280 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_49
timestamp 1607194113
transform 1 0 19844 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_14
timestamp 1607194113
transform 1 0 19568 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_14
timestamp 1607194113
transform 1 0 19476 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_15
timestamp 1607194113
transform 1 0 20764 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_15
timestamp 1607194113
transform 1 0 20672 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_48
timestamp 1607194113
transform 1 0 21040 0 1 2560
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap3_16
timestamp 1607194113
transform 1 0 21960 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_16
timestamp 1607194113
transform 1 0 21868 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_0
timestamp 1607194113
transform 1 0 2732 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_9
timestamp 1607194113
transform 1 0 1996 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_8
timestamp 1607194113
transform 1 0 1904 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_64
timestamp 1607194113
transform 1 0 3100 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_0
timestamp 1607194113
transform 1 0 2824 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_65
timestamp 1607194113
transform 1 0 4296 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_1
timestamp 1607194113
transform 1 0 4020 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_1
timestamp 1607194113
transform 1 0 3928 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_66
timestamp 1607194113
transform 1 0 5492 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_2
timestamp 1607194113
transform 1 0 5216 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_2
timestamp 1607194113
transform 1 0 5124 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_3
timestamp 1607194113
transform 1 0 6412 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_3
timestamp 1607194113
transform 1 0 6320 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_67
timestamp 1607194113
transform 1 0 6688 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_68
timestamp 1607194113
transform 1 0 7884 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_4
timestamp 1607194113
transform 1 0 7608 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_4
timestamp 1607194113
transform 1 0 7516 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_69
timestamp 1607194113
transform 1 0 9080 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_5
timestamp 1607194113
transform 1 0 8804 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_5
timestamp 1607194113
transform 1 0 8712 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_6
timestamp 1607194113
transform 1 0 10000 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_6
timestamp 1607194113
transform 1 0 9908 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_70
timestamp 1607194113
transform 1 0 10276 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_71
timestamp 1607194113
transform 1 0 11472 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_7
timestamp 1607194113
transform 1 0 11196 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_7
timestamp 1607194113
transform 1 0 11104 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_72
timestamp 1607194113
transform 1 0 12668 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_8
timestamp 1607194113
transform 1 0 12392 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_8
timestamp 1607194113
transform 1 0 12300 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_9
timestamp 1607194113
transform 1 0 13588 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_9
timestamp 1607194113
transform 1 0 13496 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_73
timestamp 1607194113
transform 1 0 13864 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_74
timestamp 1607194113
transform 1 0 15060 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_10
timestamp 1607194113
transform 1 0 14784 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_10
timestamp 1607194113
transform 1 0 14692 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_75
timestamp 1607194113
transform 1 0 16256 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_11
timestamp 1607194113
transform 1 0 15980 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_11
timestamp 1607194113
transform 1 0 15888 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_12
timestamp 1607194113
transform 1 0 17176 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_12
timestamp 1607194113
transform 1 0 17084 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_76
timestamp 1607194113
transform 1 0 17452 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_77
timestamp 1607194113
transform 1 0 18648 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_13
timestamp 1607194113
transform 1 0 18372 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_13
timestamp 1607194113
transform 1 0 18280 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_78
timestamp 1607194113
transform 1 0 19844 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_14
timestamp 1607194113
transform 1 0 19568 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_14
timestamp 1607194113
transform 1 0 19476 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_15
timestamp 1607194113
transform 1 0 20764 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_15
timestamp 1607194113
transform 1 0 20672 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_79
timestamp 1607194113
transform 1 0 21040 0 -1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap4_16
timestamp 1607194113
transform 1 0 21960 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_16
timestamp 1607194113
transform 1 0 21868 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_0
timestamp 1607194113
transform 1 0 2732 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_11
timestamp 1607194113
transform 1 0 1996 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_10
timestamp 1607194113
transform 1 0 1904 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_95
timestamp 1607194113
transform 1 0 3100 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_0
timestamp 1607194113
transform 1 0 2824 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_94
timestamp 1607194113
transform 1 0 4296 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_1
timestamp 1607194113
transform 1 0 4020 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_1
timestamp 1607194113
transform 1 0 3928 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_93
timestamp 1607194113
transform 1 0 5492 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_2
timestamp 1607194113
transform 1 0 5216 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_2
timestamp 1607194113
transform 1 0 5124 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_3
timestamp 1607194113
transform 1 0 6412 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_3
timestamp 1607194113
transform 1 0 6320 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_92
timestamp 1607194113
transform 1 0 6688 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_91
timestamp 1607194113
transform 1 0 7884 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_4
timestamp 1607194113
transform 1 0 7608 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_4
timestamp 1607194113
transform 1 0 7516 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_90
timestamp 1607194113
transform 1 0 9080 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_5
timestamp 1607194113
transform 1 0 8804 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_5
timestamp 1607194113
transform 1 0 8712 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_6
timestamp 1607194113
transform 1 0 10000 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_6
timestamp 1607194113
transform 1 0 9908 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_89
timestamp 1607194113
transform 1 0 10276 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_88
timestamp 1607194113
transform 1 0 11472 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_7
timestamp 1607194113
transform 1 0 11196 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_7
timestamp 1607194113
transform 1 0 11104 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_87
timestamp 1607194113
transform 1 0 12668 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_8
timestamp 1607194113
transform 1 0 12392 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_8
timestamp 1607194113
transform 1 0 12300 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_9
timestamp 1607194113
transform 1 0 13588 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_9
timestamp 1607194113
transform 1 0 13496 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_86
timestamp 1607194113
transform 1 0 13864 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_85
timestamp 1607194113
transform 1 0 15060 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_10
timestamp 1607194113
transform 1 0 14784 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_10
timestamp 1607194113
transform 1 0 14692 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_84
timestamp 1607194113
transform 1 0 16256 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_11
timestamp 1607194113
transform 1 0 15980 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_11
timestamp 1607194113
transform 1 0 15888 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_12
timestamp 1607194113
transform 1 0 17176 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_12
timestamp 1607194113
transform 1 0 17084 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_83
timestamp 1607194113
transform 1 0 17452 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_82
timestamp 1607194113
transform 1 0 18648 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_13
timestamp 1607194113
transform 1 0 18372 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_13
timestamp 1607194113
transform 1 0 18280 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_81
timestamp 1607194113
transform 1 0 19844 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_14
timestamp 1607194113
transform 1 0 19568 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_14
timestamp 1607194113
transform 1 0 19476 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_15
timestamp 1607194113
transform 1 0 20764 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_15
timestamp 1607194113
transform 1 0 20672 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_80
timestamp 1607194113
transform 1 0 21040 0 1 3648
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap5_16
timestamp 1607194113
transform 1 0 21960 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_16
timestamp 1607194113
transform 1 0 21868 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_0
timestamp 1607194113
transform 1 0 2732 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_15
timestamp 1607194113
transform 1 0 1996 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_14
timestamp 1607194113
transform 1 0 1904 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_0
timestamp 1607194113
transform 1 0 2732 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_13
timestamp 1607194113
transform 1 0 1996 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_12
timestamp 1607194113
transform 1 0 1904 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_127
timestamp 1607194113
transform 1 0 3100 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_0
timestamp 1607194113
transform 1 0 2824 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_96
timestamp 1607194113
transform 1 0 3100 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_0
timestamp 1607194113
transform 1 0 2824 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_126
timestamp 1607194113
transform 1 0 4296 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_1
timestamp 1607194113
transform 1 0 4020 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_1
timestamp 1607194113
transform 1 0 3928 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_97
timestamp 1607194113
transform 1 0 4296 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_1
timestamp 1607194113
transform 1 0 4020 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_1
timestamp 1607194113
transform 1 0 3928 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_125
timestamp 1607194113
transform 1 0 5492 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_2
timestamp 1607194113
transform 1 0 5216 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_2
timestamp 1607194113
transform 1 0 5124 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_98
timestamp 1607194113
transform 1 0 5492 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_2
timestamp 1607194113
transform 1 0 5216 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_2
timestamp 1607194113
transform 1 0 5124 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_3
timestamp 1607194113
transform 1 0 6412 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_3
timestamp 1607194113
transform 1 0 6320 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_3
timestamp 1607194113
transform 1 0 6412 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_3
timestamp 1607194113
transform 1 0 6320 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_124
timestamp 1607194113
transform 1 0 6688 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_99
timestamp 1607194113
transform 1 0 6688 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_123
timestamp 1607194113
transform 1 0 7884 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_4
timestamp 1607194113
transform 1 0 7608 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_4
timestamp 1607194113
transform 1 0 7516 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_100
timestamp 1607194113
transform 1 0 7884 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_4
timestamp 1607194113
transform 1 0 7608 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_4
timestamp 1607194113
transform 1 0 7516 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_122
timestamp 1607194113
transform 1 0 9080 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_5
timestamp 1607194113
transform 1 0 8804 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_5
timestamp 1607194113
transform 1 0 8712 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_101
timestamp 1607194113
transform 1 0 9080 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_5
timestamp 1607194113
transform 1 0 8804 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_5
timestamp 1607194113
transform 1 0 8712 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_6
timestamp 1607194113
transform 1 0 10000 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_6
timestamp 1607194113
transform 1 0 9908 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_6
timestamp 1607194113
transform 1 0 10000 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_6
timestamp 1607194113
transform 1 0 9908 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_121
timestamp 1607194113
transform 1 0 10276 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_102
timestamp 1607194113
transform 1 0 10276 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_120
timestamp 1607194113
transform 1 0 11472 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_7
timestamp 1607194113
transform 1 0 11196 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_7
timestamp 1607194113
transform 1 0 11104 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_103
timestamp 1607194113
transform 1 0 11472 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_7
timestamp 1607194113
transform 1 0 11196 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_7
timestamp 1607194113
transform 1 0 11104 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_119
timestamp 1607194113
transform 1 0 12668 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_8
timestamp 1607194113
transform 1 0 12392 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_8
timestamp 1607194113
transform 1 0 12300 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_104
timestamp 1607194113
transform 1 0 12668 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_8
timestamp 1607194113
transform 1 0 12392 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_8
timestamp 1607194113
transform 1 0 12300 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_9
timestamp 1607194113
transform 1 0 13588 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_9
timestamp 1607194113
transform 1 0 13496 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_9
timestamp 1607194113
transform 1 0 13588 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_9
timestamp 1607194113
transform 1 0 13496 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_118
timestamp 1607194113
transform 1 0 13864 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_105
timestamp 1607194113
transform 1 0 13864 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_117
timestamp 1607194113
transform 1 0 15060 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_10
timestamp 1607194113
transform 1 0 14784 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_10
timestamp 1607194113
transform 1 0 14692 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_106
timestamp 1607194113
transform 1 0 15060 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_10
timestamp 1607194113
transform 1 0 14784 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_10
timestamp 1607194113
transform 1 0 14692 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_116
timestamp 1607194113
transform 1 0 16256 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_11
timestamp 1607194113
transform 1 0 15980 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_11
timestamp 1607194113
transform 1 0 15888 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_107
timestamp 1607194113
transform 1 0 16256 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_11
timestamp 1607194113
transform 1 0 15980 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_11
timestamp 1607194113
transform 1 0 15888 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_12
timestamp 1607194113
transform 1 0 17176 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_12
timestamp 1607194113
transform 1 0 17084 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_12
timestamp 1607194113
transform 1 0 17176 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_12
timestamp 1607194113
transform 1 0 17084 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_115
timestamp 1607194113
transform 1 0 17452 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_108
timestamp 1607194113
transform 1 0 17452 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_114
timestamp 1607194113
transform 1 0 18648 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_13
timestamp 1607194113
transform 1 0 18372 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_13
timestamp 1607194113
transform 1 0 18280 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_109
timestamp 1607194113
transform 1 0 18648 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_13
timestamp 1607194113
transform 1 0 18372 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_13
timestamp 1607194113
transform 1 0 18280 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_113
timestamp 1607194113
transform 1 0 19844 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_14
timestamp 1607194113
transform 1 0 19568 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_14
timestamp 1607194113
transform 1 0 19476 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_110
timestamp 1607194113
transform 1 0 19844 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap6_14
timestamp 1607194113
transform 1 0 19568 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_14
timestamp 1607194113
transform 1 0 19476 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_15
timestamp 1607194113
transform 1 0 20764 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_15
timestamp 1607194113
transform 1 0 20672 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_15
timestamp 1607194113
transform 1 0 20764 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_15
timestamp 1607194113
transform 1 0 20672 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_112
timestamp 1607194113
transform 1 0 21040 0 1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_111
timestamp 1607194113
transform 1 0 21040 0 -1 4736
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap7_16
timestamp 1607194113
transform 1 0 21960 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_16
timestamp 1607194113
transform 1 0 21868 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_16
timestamp 1607194113
transform 1 0 21960 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_16
timestamp 1607194113
transform 1 0 21868 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_0
timestamp 1607194113
transform 1 0 2732 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_17
timestamp 1607194113
transform 1 0 1996 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_16
timestamp 1607194113
transform 1 0 1904 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_128
timestamp 1607194113
transform 1 0 3100 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_0
timestamp 1607194113
transform 1 0 2824 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_129
timestamp 1607194113
transform 1 0 4296 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_1
timestamp 1607194113
transform 1 0 4020 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_1
timestamp 1607194113
transform 1 0 3928 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_130
timestamp 1607194113
transform 1 0 5492 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_2
timestamp 1607194113
transform 1 0 5216 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_2
timestamp 1607194113
transform 1 0 5124 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_3
timestamp 1607194113
transform 1 0 6412 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_3
timestamp 1607194113
transform 1 0 6320 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_131
timestamp 1607194113
transform 1 0 6688 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_132
timestamp 1607194113
transform 1 0 7884 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_4
timestamp 1607194113
transform 1 0 7608 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_4
timestamp 1607194113
transform 1 0 7516 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_133
timestamp 1607194113
transform 1 0 9080 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_5
timestamp 1607194113
transform 1 0 8804 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_5
timestamp 1607194113
transform 1 0 8712 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_6
timestamp 1607194113
transform 1 0 10000 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_6
timestamp 1607194113
transform 1 0 9908 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_134
timestamp 1607194113
transform 1 0 10276 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_135
timestamp 1607194113
transform 1 0 11472 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_7
timestamp 1607194113
transform 1 0 11196 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_7
timestamp 1607194113
transform 1 0 11104 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_136
timestamp 1607194113
transform 1 0 12668 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_8
timestamp 1607194113
transform 1 0 12392 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_8
timestamp 1607194113
transform 1 0 12300 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_9
timestamp 1607194113
transform 1 0 13588 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_9
timestamp 1607194113
transform 1 0 13496 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_137
timestamp 1607194113
transform 1 0 13864 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_138
timestamp 1607194113
transform 1 0 15060 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_10
timestamp 1607194113
transform 1 0 14784 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_10
timestamp 1607194113
transform 1 0 14692 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_139
timestamp 1607194113
transform 1 0 16256 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_11
timestamp 1607194113
transform 1 0 15980 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_11
timestamp 1607194113
transform 1 0 15888 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_12
timestamp 1607194113
transform 1 0 17176 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_12
timestamp 1607194113
transform 1 0 17084 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_140
timestamp 1607194113
transform 1 0 17452 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_141
timestamp 1607194113
transform 1 0 18648 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_13
timestamp 1607194113
transform 1 0 18372 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_13
timestamp 1607194113
transform 1 0 18280 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_142
timestamp 1607194113
transform 1 0 19844 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_14
timestamp 1607194113
transform 1 0 19568 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_14
timestamp 1607194113
transform 1 0 19476 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_15
timestamp 1607194113
transform 1 0 20764 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_15
timestamp 1607194113
transform 1 0 20672 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_143
timestamp 1607194113
transform 1 0 21040 0 -1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap8_16
timestamp 1607194113
transform 1 0 21960 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_16
timestamp 1607194113
transform 1 0 21868 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_0
timestamp 1607194113
transform 1 0 2732 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_19
timestamp 1607194113
transform 1 0 1996 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_18
timestamp 1607194113
transform 1 0 1904 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_159
timestamp 1607194113
transform 1 0 3100 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_0
timestamp 1607194113
transform 1 0 2824 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_158
timestamp 1607194113
transform 1 0 4296 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_1
timestamp 1607194113
transform 1 0 4020 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_1
timestamp 1607194113
transform 1 0 3928 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_157
timestamp 1607194113
transform 1 0 5492 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_2
timestamp 1607194113
transform 1 0 5216 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_2
timestamp 1607194113
transform 1 0 5124 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_3
timestamp 1607194113
transform 1 0 6412 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_3
timestamp 1607194113
transform 1 0 6320 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_156
timestamp 1607194113
transform 1 0 6688 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_155
timestamp 1607194113
transform 1 0 7884 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_4
timestamp 1607194113
transform 1 0 7608 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_4
timestamp 1607194113
transform 1 0 7516 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_154
timestamp 1607194113
transform 1 0 9080 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_5
timestamp 1607194113
transform 1 0 8804 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_5
timestamp 1607194113
transform 1 0 8712 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_6
timestamp 1607194113
transform 1 0 10000 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_6
timestamp 1607194113
transform 1 0 9908 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_153
timestamp 1607194113
transform 1 0 10276 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_152
timestamp 1607194113
transform 1 0 11472 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_7
timestamp 1607194113
transform 1 0 11196 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_7
timestamp 1607194113
transform 1 0 11104 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_151
timestamp 1607194113
transform 1 0 12668 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_8
timestamp 1607194113
transform 1 0 12392 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_8
timestamp 1607194113
transform 1 0 12300 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_9
timestamp 1607194113
transform 1 0 13588 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_9
timestamp 1607194113
transform 1 0 13496 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_150
timestamp 1607194113
transform 1 0 13864 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_149
timestamp 1607194113
transform 1 0 15060 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_10
timestamp 1607194113
transform 1 0 14784 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_10
timestamp 1607194113
transform 1 0 14692 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_148
timestamp 1607194113
transform 1 0 16256 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_11
timestamp 1607194113
transform 1 0 15980 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_11
timestamp 1607194113
transform 1 0 15888 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_12
timestamp 1607194113
transform 1 0 17176 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_12
timestamp 1607194113
transform 1 0 17084 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_147
timestamp 1607194113
transform 1 0 17452 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_146
timestamp 1607194113
transform 1 0 18648 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_13
timestamp 1607194113
transform 1 0 18372 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_13
timestamp 1607194113
transform 1 0 18280 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_145
timestamp 1607194113
transform 1 0 19844 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_14
timestamp 1607194113
transform 1 0 19568 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_14
timestamp 1607194113
transform 1 0 19476 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_15
timestamp 1607194113
transform 1 0 20764 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_15
timestamp 1607194113
transform 1 0 20672 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_144
timestamp 1607194113
transform 1 0 21040 0 1 5824
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap9_16
timestamp 1607194113
transform 1 0 21960 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_16
timestamp 1607194113
transform 1 0 21868 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_0
timestamp 1607194113
transform 1 0 2732 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_21
timestamp 1607194113
transform 1 0 1996 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_20
timestamp 1607194113
transform 1 0 1904 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_160
timestamp 1607194113
transform 1 0 3100 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_0
timestamp 1607194113
transform 1 0 2824 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_161
timestamp 1607194113
transform 1 0 4296 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_1
timestamp 1607194113
transform 1 0 4020 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_1
timestamp 1607194113
transform 1 0 3928 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_162
timestamp 1607194113
transform 1 0 5492 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_2
timestamp 1607194113
transform 1 0 5216 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_2
timestamp 1607194113
transform 1 0 5124 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_3
timestamp 1607194113
transform 1 0 6412 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_3
timestamp 1607194113
transform 1 0 6320 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_163
timestamp 1607194113
transform 1 0 6688 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_164
timestamp 1607194113
transform 1 0 7884 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_4
timestamp 1607194113
transform 1 0 7608 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_4
timestamp 1607194113
transform 1 0 7516 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_165
timestamp 1607194113
transform 1 0 9080 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_5
timestamp 1607194113
transform 1 0 8804 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_5
timestamp 1607194113
transform 1 0 8712 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_6
timestamp 1607194113
transform 1 0 10000 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_6
timestamp 1607194113
transform 1 0 9908 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_166
timestamp 1607194113
transform 1 0 10276 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_167
timestamp 1607194113
transform 1 0 11472 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_7
timestamp 1607194113
transform 1 0 11196 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_7
timestamp 1607194113
transform 1 0 11104 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_168
timestamp 1607194113
transform 1 0 12668 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_8
timestamp 1607194113
transform 1 0 12392 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_8
timestamp 1607194113
transform 1 0 12300 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_9
timestamp 1607194113
transform 1 0 13588 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_9
timestamp 1607194113
transform 1 0 13496 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_169
timestamp 1607194113
transform 1 0 13864 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_170
timestamp 1607194113
transform 1 0 15060 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_10
timestamp 1607194113
transform 1 0 14784 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_10
timestamp 1607194113
transform 1 0 14692 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_171
timestamp 1607194113
transform 1 0 16256 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_11
timestamp 1607194113
transform 1 0 15980 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_11
timestamp 1607194113
transform 1 0 15888 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_12
timestamp 1607194113
transform 1 0 17176 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_12
timestamp 1607194113
transform 1 0 17084 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_172
timestamp 1607194113
transform 1 0 17452 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_173
timestamp 1607194113
transform 1 0 18648 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_13
timestamp 1607194113
transform 1 0 18372 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_13
timestamp 1607194113
transform 1 0 18280 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_174
timestamp 1607194113
transform 1 0 19844 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_14
timestamp 1607194113
transform 1 0 19568 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_14
timestamp 1607194113
transform 1 0 19476 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_15
timestamp 1607194113
transform 1 0 20764 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_15
timestamp 1607194113
transform 1 0 20672 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_175
timestamp 1607194113
transform 1 0 21040 0 -1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap10_16
timestamp 1607194113
transform 1 0 21960 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_16
timestamp 1607194113
transform 1 0 21868 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_0
timestamp 1607194113
transform 1 0 2732 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_23
timestamp 1607194113
transform 1 0 1996 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_22
timestamp 1607194113
transform 1 0 1904 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_191
timestamp 1607194113
transform 1 0 3100 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_0
timestamp 1607194113
transform 1 0 2824 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_190
timestamp 1607194113
transform 1 0 4296 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_1
timestamp 1607194113
transform 1 0 4020 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_1
timestamp 1607194113
transform 1 0 3928 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_189
timestamp 1607194113
transform 1 0 5492 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_2
timestamp 1607194113
transform 1 0 5216 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_2
timestamp 1607194113
transform 1 0 5124 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_3
timestamp 1607194113
transform 1 0 6412 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_3
timestamp 1607194113
transform 1 0 6320 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_188
timestamp 1607194113
transform 1 0 6688 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_187
timestamp 1607194113
transform 1 0 7884 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_4
timestamp 1607194113
transform 1 0 7608 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_4
timestamp 1607194113
transform 1 0 7516 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_186
timestamp 1607194113
transform 1 0 9080 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_5
timestamp 1607194113
transform 1 0 8804 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_5
timestamp 1607194113
transform 1 0 8712 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_6
timestamp 1607194113
transform 1 0 10000 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_6
timestamp 1607194113
transform 1 0 9908 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_185
timestamp 1607194113
transform 1 0 10276 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_184
timestamp 1607194113
transform 1 0 11472 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_7
timestamp 1607194113
transform 1 0 11196 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_7
timestamp 1607194113
transform 1 0 11104 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_183
timestamp 1607194113
transform 1 0 12668 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_8
timestamp 1607194113
transform 1 0 12392 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_8
timestamp 1607194113
transform 1 0 12300 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_9
timestamp 1607194113
transform 1 0 13588 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_9
timestamp 1607194113
transform 1 0 13496 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_182
timestamp 1607194113
transform 1 0 13864 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_181
timestamp 1607194113
transform 1 0 15060 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_10
timestamp 1607194113
transform 1 0 14784 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_10
timestamp 1607194113
transform 1 0 14692 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_180
timestamp 1607194113
transform 1 0 16256 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_11
timestamp 1607194113
transform 1 0 15980 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_11
timestamp 1607194113
transform 1 0 15888 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_12
timestamp 1607194113
transform 1 0 17176 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_12
timestamp 1607194113
transform 1 0 17084 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_179
timestamp 1607194113
transform 1 0 17452 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_178
timestamp 1607194113
transform 1 0 18648 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_13
timestamp 1607194113
transform 1 0 18372 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_13
timestamp 1607194113
transform 1 0 18280 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_177
timestamp 1607194113
transform 1 0 19844 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_14
timestamp 1607194113
transform 1 0 19568 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_14
timestamp 1607194113
transform 1 0 19476 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_15
timestamp 1607194113
transform 1 0 20764 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_15
timestamp 1607194113
transform 1 0 20672 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_176
timestamp 1607194113
transform 1 0 21040 0 1 6912
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap11_16
timestamp 1607194113
transform 1 0 21960 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_16
timestamp 1607194113
transform 1 0 21868 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_0
timestamp 1607194113
transform 1 0 2732 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_25
timestamp 1607194113
transform 1 0 1996 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_24
timestamp 1607194113
transform 1 0 1904 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_192
timestamp 1607194113
transform 1 0 3100 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_0
timestamp 1607194113
transform 1 0 2824 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_193
timestamp 1607194113
transform 1 0 4296 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_1
timestamp 1607194113
transform 1 0 4020 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_1
timestamp 1607194113
transform 1 0 3928 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_194
timestamp 1607194113
transform 1 0 5492 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_2
timestamp 1607194113
transform 1 0 5216 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_2
timestamp 1607194113
transform 1 0 5124 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_3
timestamp 1607194113
transform 1 0 6412 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_3
timestamp 1607194113
transform 1 0 6320 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_195
timestamp 1607194113
transform 1 0 6688 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_196
timestamp 1607194113
transform 1 0 7884 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_4
timestamp 1607194113
transform 1 0 7608 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_4
timestamp 1607194113
transform 1 0 7516 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_197
timestamp 1607194113
transform 1 0 9080 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_5
timestamp 1607194113
transform 1 0 8804 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_5
timestamp 1607194113
transform 1 0 8712 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_6
timestamp 1607194113
transform 1 0 10000 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_6
timestamp 1607194113
transform 1 0 9908 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_198
timestamp 1607194113
transform 1 0 10276 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_199
timestamp 1607194113
transform 1 0 11472 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_7
timestamp 1607194113
transform 1 0 11196 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_7
timestamp 1607194113
transform 1 0 11104 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_200
timestamp 1607194113
transform 1 0 12668 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_8
timestamp 1607194113
transform 1 0 12392 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_8
timestamp 1607194113
transform 1 0 12300 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_9
timestamp 1607194113
transform 1 0 13588 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_9
timestamp 1607194113
transform 1 0 13496 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_201
timestamp 1607194113
transform 1 0 13864 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_202
timestamp 1607194113
transform 1 0 15060 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_10
timestamp 1607194113
transform 1 0 14784 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_10
timestamp 1607194113
transform 1 0 14692 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_203
timestamp 1607194113
transform 1 0 16256 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_11
timestamp 1607194113
transform 1 0 15980 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_11
timestamp 1607194113
transform 1 0 15888 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_12
timestamp 1607194113
transform 1 0 17176 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_12
timestamp 1607194113
transform 1 0 17084 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_204
timestamp 1607194113
transform 1 0 17452 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_205
timestamp 1607194113
transform 1 0 18648 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_13
timestamp 1607194113
transform 1 0 18372 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_13
timestamp 1607194113
transform 1 0 18280 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_206
timestamp 1607194113
transform 1 0 19844 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_14
timestamp 1607194113
transform 1 0 19568 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_14
timestamp 1607194113
transform 1 0 19476 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_15
timestamp 1607194113
transform 1 0 20764 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_15
timestamp 1607194113
transform 1 0 20672 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_207
timestamp 1607194113
transform 1 0 21040 0 -1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap12_16
timestamp 1607194113
transform 1 0 21960 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_16
timestamp 1607194113
transform 1 0 21868 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_0
timestamp 1607194113
transform 1 0 2732 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_29
timestamp 1607194113
transform 1 0 1996 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_28
timestamp 1607194113
transform 1 0 1904 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_0
timestamp 1607194113
transform 1 0 2732 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_27
timestamp 1607194113
transform 1 0 1996 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_26
timestamp 1607194113
transform 1 0 1904 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_224
timestamp 1607194113
transform 1 0 3100 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_0
timestamp 1607194113
transform 1 0 2824 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_223
timestamp 1607194113
transform 1 0 3100 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_0
timestamp 1607194113
transform 1 0 2824 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_225
timestamp 1607194113
transform 1 0 4296 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_1
timestamp 1607194113
transform 1 0 4020 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_1
timestamp 1607194113
transform 1 0 3928 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_222
timestamp 1607194113
transform 1 0 4296 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_1
timestamp 1607194113
transform 1 0 4020 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_1
timestamp 1607194113
transform 1 0 3928 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_226
timestamp 1607194113
transform 1 0 5492 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_2
timestamp 1607194113
transform 1 0 5216 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_2
timestamp 1607194113
transform 1 0 5124 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_221
timestamp 1607194113
transform 1 0 5492 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_2
timestamp 1607194113
transform 1 0 5216 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_2
timestamp 1607194113
transform 1 0 5124 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_3
timestamp 1607194113
transform 1 0 6412 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_3
timestamp 1607194113
transform 1 0 6320 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_3
timestamp 1607194113
transform 1 0 6412 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_3
timestamp 1607194113
transform 1 0 6320 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_227
timestamp 1607194113
transform 1 0 6688 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_220
timestamp 1607194113
transform 1 0 6688 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_228
timestamp 1607194113
transform 1 0 7884 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_4
timestamp 1607194113
transform 1 0 7608 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_4
timestamp 1607194113
transform 1 0 7516 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_219
timestamp 1607194113
transform 1 0 7884 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_4
timestamp 1607194113
transform 1 0 7608 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_4
timestamp 1607194113
transform 1 0 7516 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_229
timestamp 1607194113
transform 1 0 9080 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_5
timestamp 1607194113
transform 1 0 8804 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_5
timestamp 1607194113
transform 1 0 8712 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_218
timestamp 1607194113
transform 1 0 9080 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_5
timestamp 1607194113
transform 1 0 8804 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_5
timestamp 1607194113
transform 1 0 8712 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_6
timestamp 1607194113
transform 1 0 10000 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_6
timestamp 1607194113
transform 1 0 9908 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_6
timestamp 1607194113
transform 1 0 10000 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_6
timestamp 1607194113
transform 1 0 9908 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_230
timestamp 1607194113
transform 1 0 10276 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_217
timestamp 1607194113
transform 1 0 10276 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_231
timestamp 1607194113
transform 1 0 11472 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_7
timestamp 1607194113
transform 1 0 11196 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_7
timestamp 1607194113
transform 1 0 11104 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_216
timestamp 1607194113
transform 1 0 11472 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_7
timestamp 1607194113
transform 1 0 11196 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_7
timestamp 1607194113
transform 1 0 11104 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_232
timestamp 1607194113
transform 1 0 12668 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_8
timestamp 1607194113
transform 1 0 12392 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_8
timestamp 1607194113
transform 1 0 12300 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_215
timestamp 1607194113
transform 1 0 12668 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_8
timestamp 1607194113
transform 1 0 12392 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_8
timestamp 1607194113
transform 1 0 12300 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_9
timestamp 1607194113
transform 1 0 13588 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_9
timestamp 1607194113
transform 1 0 13496 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_9
timestamp 1607194113
transform 1 0 13588 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_9
timestamp 1607194113
transform 1 0 13496 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_233
timestamp 1607194113
transform 1 0 13864 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_214
timestamp 1607194113
transform 1 0 13864 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_234
timestamp 1607194113
transform 1 0 15060 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_10
timestamp 1607194113
transform 1 0 14784 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_10
timestamp 1607194113
transform 1 0 14692 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_213
timestamp 1607194113
transform 1 0 15060 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_10
timestamp 1607194113
transform 1 0 14784 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_10
timestamp 1607194113
transform 1 0 14692 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_235
timestamp 1607194113
transform 1 0 16256 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_11
timestamp 1607194113
transform 1 0 15980 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_11
timestamp 1607194113
transform 1 0 15888 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_212
timestamp 1607194113
transform 1 0 16256 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_11
timestamp 1607194113
transform 1 0 15980 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_11
timestamp 1607194113
transform 1 0 15888 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_12
timestamp 1607194113
transform 1 0 17176 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_12
timestamp 1607194113
transform 1 0 17084 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_12
timestamp 1607194113
transform 1 0 17176 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_12
timestamp 1607194113
transform 1 0 17084 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_236
timestamp 1607194113
transform 1 0 17452 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_211
timestamp 1607194113
transform 1 0 17452 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_237
timestamp 1607194113
transform 1 0 18648 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_13
timestamp 1607194113
transform 1 0 18372 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_13
timestamp 1607194113
transform 1 0 18280 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_210
timestamp 1607194113
transform 1 0 18648 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_13
timestamp 1607194113
transform 1 0 18372 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_13
timestamp 1607194113
transform 1 0 18280 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_238
timestamp 1607194113
transform 1 0 19844 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_14
timestamp 1607194113
transform 1 0 19568 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_14
timestamp 1607194113
transform 1 0 19476 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_209
timestamp 1607194113
transform 1 0 19844 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap13_14
timestamp 1607194113
transform 1 0 19568 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_14
timestamp 1607194113
transform 1 0 19476 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_15
timestamp 1607194113
transform 1 0 20764 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_15
timestamp 1607194113
transform 1 0 20672 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_15
timestamp 1607194113
transform 1 0 20764 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_15
timestamp 1607194113
transform 1 0 20672 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_239
timestamp 1607194113
transform 1 0 21040 0 -1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_208
timestamp 1607194113
transform 1 0 21040 0 1 8000
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap14_16
timestamp 1607194113
transform 1 0 21960 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_16
timestamp 1607194113
transform 1 0 21868 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_16
timestamp 1607194113
transform 1 0 21960 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_16
timestamp 1607194113
transform 1 0 21868 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_0
timestamp 1607194113
transform 1 0 2732 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1904 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_255
timestamp 1607194113
transform 1 0 3100 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_0
timestamp 1607194113
transform 1 0 2824 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_254
timestamp 1607194113
transform 1 0 4296 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_1
timestamp 1607194113
transform 1 0 4020 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_1
timestamp 1607194113
transform 1 0 3928 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_253
timestamp 1607194113
transform 1 0 5492 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_2
timestamp 1607194113
transform 1 0 5216 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_2
timestamp 1607194113
transform 1 0 5124 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_3
timestamp 1607194113
transform 1 0 6412 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_3
timestamp 1607194113
transform 1 0 6320 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_252
timestamp 1607194113
transform 1 0 6688 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_251
timestamp 1607194113
transform 1 0 7884 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_4
timestamp 1607194113
transform 1 0 7608 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_4
timestamp 1607194113
transform 1 0 7516 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_250
timestamp 1607194113
transform 1 0 9080 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_5
timestamp 1607194113
transform 1 0 8804 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_5
timestamp 1607194113
transform 1 0 8712 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_6
timestamp 1607194113
transform 1 0 10000 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_6
timestamp 1607194113
transform 1 0 9908 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_249
timestamp 1607194113
transform 1 0 10276 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_248
timestamp 1607194113
transform 1 0 11472 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_7
timestamp 1607194113
transform 1 0 11196 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_7
timestamp 1607194113
transform 1 0 11104 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_247
timestamp 1607194113
transform 1 0 12668 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_8
timestamp 1607194113
transform 1 0 12392 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_8
timestamp 1607194113
transform 1 0 12300 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_9
timestamp 1607194113
transform 1 0 13588 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_9
timestamp 1607194113
transform 1 0 13496 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_246
timestamp 1607194113
transform 1 0 13864 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_245
timestamp 1607194113
transform 1 0 15060 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_10
timestamp 1607194113
transform 1 0 14784 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_10
timestamp 1607194113
transform 1 0 14692 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_244
timestamp 1607194113
transform 1 0 16256 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_11
timestamp 1607194113
transform 1 0 15980 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_11
timestamp 1607194113
transform 1 0 15888 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_12
timestamp 1607194113
transform 1 0 17176 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_12
timestamp 1607194113
transform 1 0 17084 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_243
timestamp 1607194113
transform 1 0 17452 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_242
timestamp 1607194113
transform 1 0 18648 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_13
timestamp 1607194113
transform 1 0 18372 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_13
timestamp 1607194113
transform 1 0 18280 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_241
timestamp 1607194113
transform 1 0 19844 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_14
timestamp 1607194113
transform 1 0 19568 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_14
timestamp 1607194113
transform 1 0 19476 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_15
timestamp 1607194113
transform 1 0 20764 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_15
timestamp 1607194113
transform 1 0 20672 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_8_240
timestamp 1607194113
transform 1 0 21040 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap15_16
timestamp 1607194113
transform 1 0 21960 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_16
timestamp 1607194113
transform 1 0 21868 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_0
timestamp 1607194113
transform 1 0 2732 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_31
timestamp 1607194113
transform 1 0 1996 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_30
timestamp 1607194113
transform 1 0 1904 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_0
timestamp 1607194113
transform 1 0 3100 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_0
timestamp 1607194113
transform 1 0 2824 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_1
timestamp 1607194113
transform 1 0 4296 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_1
timestamp 1607194113
transform 1 0 4020 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_1
timestamp 1607194113
transform 1 0 3928 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_2
timestamp 1607194113
transform 1 0 5492 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_2
timestamp 1607194113
transform 1 0 5216 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_2
timestamp 1607194113
transform 1 0 5124 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_3
timestamp 1607194113
transform 1 0 6412 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_3
timestamp 1607194113
transform 1 0 6320 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_3
timestamp 1607194113
transform 1 0 6688 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_4
timestamp 1607194113
transform 1 0 7884 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_4
timestamp 1607194113
transform 1 0 7608 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_4
timestamp 1607194113
transform 1 0 7516 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_5
timestamp 1607194113
transform 1 0 9080 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_5
timestamp 1607194113
transform 1 0 8804 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_5
timestamp 1607194113
transform 1 0 8712 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_6
timestamp 1607194113
transform 1 0 10000 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_6
timestamp 1607194113
transform 1 0 9908 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_6
timestamp 1607194113
transform 1 0 10276 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_7
timestamp 1607194113
transform 1 0 11472 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_7
timestamp 1607194113
transform 1 0 11196 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_7
timestamp 1607194113
transform 1 0 11104 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_8
timestamp 1607194113
transform 1 0 12668 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_8
timestamp 1607194113
transform 1 0 12392 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_8
timestamp 1607194113
transform 1 0 12300 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_9
timestamp 1607194113
transform 1 0 13588 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_9
timestamp 1607194113
transform 1 0 13496 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_9
timestamp 1607194113
transform 1 0 13864 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_10
timestamp 1607194113
transform 1 0 15060 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_10
timestamp 1607194113
transform 1 0 14784 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_10
timestamp 1607194113
transform 1 0 14692 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_11
timestamp 1607194113
transform 1 0 16256 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_11
timestamp 1607194113
transform 1 0 15980 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_11
timestamp 1607194113
transform 1 0 15888 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_12
timestamp 1607194113
transform 1 0 17176 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_12
timestamp 1607194113
transform 1 0 17084 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_12
timestamp 1607194113
transform 1 0 17452 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_13
timestamp 1607194113
transform 1 0 18648 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_13
timestamp 1607194113
transform 1 0 18372 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_13
timestamp 1607194113
transform 1 0 18280 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_14
timestamp 1607194113
transform 1 0 19844 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_14
timestamp 1607194113
transform 1 0 19568 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_14
timestamp 1607194113
transform 1 0 19476 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_15
timestamp 1607194113
transform 1 0 20764 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_15
timestamp 1607194113
transform 1 0 20672 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_15
timestamp 1607194113
transform 1 0 21040 0 -1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap16_16
timestamp 1607194113
transform 1 0 21960 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_16
timestamp 1607194113
transform 1 0 21868 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_0
timestamp 1607194113
transform 1 0 2732 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_33
timestamp 1607194113
transform 1 0 1996 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_32
timestamp 1607194113
transform 1 0 1904 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_31
timestamp 1607194113
transform 1 0 3100 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_0
timestamp 1607194113
transform 1 0 2824 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_30
timestamp 1607194113
transform 1 0 4296 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_1
timestamp 1607194113
transform 1 0 4020 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_1
timestamp 1607194113
transform 1 0 3928 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_29
timestamp 1607194113
transform 1 0 5492 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_2
timestamp 1607194113
transform 1 0 5216 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_2
timestamp 1607194113
transform 1 0 5124 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_3
timestamp 1607194113
transform 1 0 6412 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_3
timestamp 1607194113
transform 1 0 6320 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_28
timestamp 1607194113
transform 1 0 6688 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_27
timestamp 1607194113
transform 1 0 7884 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_4
timestamp 1607194113
transform 1 0 7608 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_4
timestamp 1607194113
transform 1 0 7516 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_26
timestamp 1607194113
transform 1 0 9080 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_5
timestamp 1607194113
transform 1 0 8804 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_5
timestamp 1607194113
transform 1 0 8712 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_6
timestamp 1607194113
transform 1 0 10000 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_6
timestamp 1607194113
transform 1 0 9908 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_25
timestamp 1607194113
transform 1 0 10276 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_24
timestamp 1607194113
transform 1 0 11472 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_7
timestamp 1607194113
transform 1 0 11196 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_7
timestamp 1607194113
transform 1 0 11104 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_23
timestamp 1607194113
transform 1 0 12668 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_8
timestamp 1607194113
transform 1 0 12392 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_8
timestamp 1607194113
transform 1 0 12300 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_9
timestamp 1607194113
transform 1 0 13588 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_9
timestamp 1607194113
transform 1 0 13496 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_22
timestamp 1607194113
transform 1 0 13864 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_21
timestamp 1607194113
transform 1 0 15060 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_10
timestamp 1607194113
transform 1 0 14784 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_10
timestamp 1607194113
transform 1 0 14692 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_20
timestamp 1607194113
transform 1 0 16256 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_11
timestamp 1607194113
transform 1 0 15980 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_11
timestamp 1607194113
transform 1 0 15888 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_12
timestamp 1607194113
transform 1 0 17176 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_12
timestamp 1607194113
transform 1 0 17084 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_19
timestamp 1607194113
transform 1 0 17452 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_18
timestamp 1607194113
transform 1 0 18648 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_13
timestamp 1607194113
transform 1 0 18372 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_13
timestamp 1607194113
transform 1 0 18280 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_17
timestamp 1607194113
transform 1 0 19844 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_14
timestamp 1607194113
transform 1 0 19568 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_14
timestamp 1607194113
transform 1 0 19476 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_15
timestamp 1607194113
transform 1 0 20764 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_15
timestamp 1607194113
transform 1 0 20672 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_16
timestamp 1607194113
transform 1 0 21040 0 1 10176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap17_16
timestamp 1607194113
transform 1 0 21960 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_16
timestamp 1607194113
transform 1 0 21868 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_0
timestamp 1607194113
transform 1 0 2732 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_35
timestamp 1607194113
transform 1 0 1996 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_34
timestamp 1607194113
transform 1 0 1904 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_32
timestamp 1607194113
transform 1 0 3100 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_0
timestamp 1607194113
transform 1 0 2824 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_33
timestamp 1607194113
transform 1 0 4296 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_1
timestamp 1607194113
transform 1 0 4020 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_1
timestamp 1607194113
transform 1 0 3928 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_34
timestamp 1607194113
transform 1 0 5492 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_2
timestamp 1607194113
transform 1 0 5216 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_2
timestamp 1607194113
transform 1 0 5124 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_3
timestamp 1607194113
transform 1 0 6412 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_3
timestamp 1607194113
transform 1 0 6320 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_35
timestamp 1607194113
transform 1 0 6688 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_36
timestamp 1607194113
transform 1 0 7884 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_4
timestamp 1607194113
transform 1 0 7608 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_4
timestamp 1607194113
transform 1 0 7516 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_37
timestamp 1607194113
transform 1 0 9080 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_5
timestamp 1607194113
transform 1 0 8804 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_5
timestamp 1607194113
transform 1 0 8712 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_6
timestamp 1607194113
transform 1 0 10000 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_6
timestamp 1607194113
transform 1 0 9908 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_38
timestamp 1607194113
transform 1 0 10276 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_39
timestamp 1607194113
transform 1 0 11472 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_7
timestamp 1607194113
transform 1 0 11196 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_7
timestamp 1607194113
transform 1 0 11104 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_40
timestamp 1607194113
transform 1 0 12668 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_8
timestamp 1607194113
transform 1 0 12392 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_8
timestamp 1607194113
transform 1 0 12300 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_9
timestamp 1607194113
transform 1 0 13588 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_9
timestamp 1607194113
transform 1 0 13496 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_41
timestamp 1607194113
transform 1 0 13864 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_42
timestamp 1607194113
transform 1 0 15060 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_10
timestamp 1607194113
transform 1 0 14784 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_10
timestamp 1607194113
transform 1 0 14692 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_43
timestamp 1607194113
transform 1 0 16256 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_11
timestamp 1607194113
transform 1 0 15980 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_11
timestamp 1607194113
transform 1 0 15888 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_12
timestamp 1607194113
transform 1 0 17176 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_12
timestamp 1607194113
transform 1 0 17084 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_44
timestamp 1607194113
transform 1 0 17452 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_45
timestamp 1607194113
transform 1 0 18648 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_13
timestamp 1607194113
transform 1 0 18372 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_13
timestamp 1607194113
transform 1 0 18280 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_46
timestamp 1607194113
transform 1 0 19844 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_14
timestamp 1607194113
transform 1 0 19568 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_14
timestamp 1607194113
transform 1 0 19476 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_15
timestamp 1607194113
transform 1 0 20764 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_15
timestamp 1607194113
transform 1 0 20672 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_47
timestamp 1607194113
transform 1 0 21040 0 -1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap18_16
timestamp 1607194113
transform 1 0 21960 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_16
timestamp 1607194113
transform 1 0 21868 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_0
timestamp 1607194113
transform 1 0 2732 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_39
timestamp 1607194113
transform 1 0 1996 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_38
timestamp 1607194113
transform 1 0 1904 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_0
timestamp 1607194113
transform 1 0 2732 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_37
timestamp 1607194113
transform 1 0 1996 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_36
timestamp 1607194113
transform 1 0 1904 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_64
timestamp 1607194113
transform 1 0 3100 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_0
timestamp 1607194113
transform 1 0 2824 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_63
timestamp 1607194113
transform 1 0 3100 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_0
timestamp 1607194113
transform 1 0 2824 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_65
timestamp 1607194113
transform 1 0 4296 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_1
timestamp 1607194113
transform 1 0 4020 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_1
timestamp 1607194113
transform 1 0 3928 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_62
timestamp 1607194113
transform 1 0 4296 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_1
timestamp 1607194113
transform 1 0 4020 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_1
timestamp 1607194113
transform 1 0 3928 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_66
timestamp 1607194113
transform 1 0 5492 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_2
timestamp 1607194113
transform 1 0 5216 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_2
timestamp 1607194113
transform 1 0 5124 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_61
timestamp 1607194113
transform 1 0 5492 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_2
timestamp 1607194113
transform 1 0 5216 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_2
timestamp 1607194113
transform 1 0 5124 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_3
timestamp 1607194113
transform 1 0 6412 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_3
timestamp 1607194113
transform 1 0 6320 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_3
timestamp 1607194113
transform 1 0 6412 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_3
timestamp 1607194113
transform 1 0 6320 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_67
timestamp 1607194113
transform 1 0 6688 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_60
timestamp 1607194113
transform 1 0 6688 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_68
timestamp 1607194113
transform 1 0 7884 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_4
timestamp 1607194113
transform 1 0 7608 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_4
timestamp 1607194113
transform 1 0 7516 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_59
timestamp 1607194113
transform 1 0 7884 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_4
timestamp 1607194113
transform 1 0 7608 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_4
timestamp 1607194113
transform 1 0 7516 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_69
timestamp 1607194113
transform 1 0 9080 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_5
timestamp 1607194113
transform 1 0 8804 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_5
timestamp 1607194113
transform 1 0 8712 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_58
timestamp 1607194113
transform 1 0 9080 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_5
timestamp 1607194113
transform 1 0 8804 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_5
timestamp 1607194113
transform 1 0 8712 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_6
timestamp 1607194113
transform 1 0 10000 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_6
timestamp 1607194113
transform 1 0 9908 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_6
timestamp 1607194113
transform 1 0 10000 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_6
timestamp 1607194113
transform 1 0 9908 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_70
timestamp 1607194113
transform 1 0 10276 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_57
timestamp 1607194113
transform 1 0 10276 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_71
timestamp 1607194113
transform 1 0 11472 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_7
timestamp 1607194113
transform 1 0 11196 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_7
timestamp 1607194113
transform 1 0 11104 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_56
timestamp 1607194113
transform 1 0 11472 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_7
timestamp 1607194113
transform 1 0 11196 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_7
timestamp 1607194113
transform 1 0 11104 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_72
timestamp 1607194113
transform 1 0 12668 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_8
timestamp 1607194113
transform 1 0 12392 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_8
timestamp 1607194113
transform 1 0 12300 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_55
timestamp 1607194113
transform 1 0 12668 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_8
timestamp 1607194113
transform 1 0 12392 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_8
timestamp 1607194113
transform 1 0 12300 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_9
timestamp 1607194113
transform 1 0 13588 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_9
timestamp 1607194113
transform 1 0 13496 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_9
timestamp 1607194113
transform 1 0 13588 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_9
timestamp 1607194113
transform 1 0 13496 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_73
timestamp 1607194113
transform 1 0 13864 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_54
timestamp 1607194113
transform 1 0 13864 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_74
timestamp 1607194113
transform 1 0 15060 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_10
timestamp 1607194113
transform 1 0 14784 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_10
timestamp 1607194113
transform 1 0 14692 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_53
timestamp 1607194113
transform 1 0 15060 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_10
timestamp 1607194113
transform 1 0 14784 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_10
timestamp 1607194113
transform 1 0 14692 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_75
timestamp 1607194113
transform 1 0 16256 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_11
timestamp 1607194113
transform 1 0 15980 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_11
timestamp 1607194113
transform 1 0 15888 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_52
timestamp 1607194113
transform 1 0 16256 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_11
timestamp 1607194113
transform 1 0 15980 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_11
timestamp 1607194113
transform 1 0 15888 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_12
timestamp 1607194113
transform 1 0 17176 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_12
timestamp 1607194113
transform 1 0 17084 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_12
timestamp 1607194113
transform 1 0 17176 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_12
timestamp 1607194113
transform 1 0 17084 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_76
timestamp 1607194113
transform 1 0 17452 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_51
timestamp 1607194113
transform 1 0 17452 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_77
timestamp 1607194113
transform 1 0 18648 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_13
timestamp 1607194113
transform 1 0 18372 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_13
timestamp 1607194113
transform 1 0 18280 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_50
timestamp 1607194113
transform 1 0 18648 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_13
timestamp 1607194113
transform 1 0 18372 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_13
timestamp 1607194113
transform 1 0 18280 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_78
timestamp 1607194113
transform 1 0 19844 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_14
timestamp 1607194113
transform 1 0 19568 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_14
timestamp 1607194113
transform 1 0 19476 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_49
timestamp 1607194113
transform 1 0 19844 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap19_14
timestamp 1607194113
transform 1 0 19568 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_14
timestamp 1607194113
transform 1 0 19476 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_15
timestamp 1607194113
transform 1 0 20764 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_15
timestamp 1607194113
transform 1 0 20672 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_15
timestamp 1607194113
transform 1 0 20764 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_15
timestamp 1607194113
transform 1 0 20672 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_79
timestamp 1607194113
transform 1 0 21040 0 -1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_48
timestamp 1607194113
transform 1 0 21040 0 1 11264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap20_16
timestamp 1607194113
transform 1 0 21960 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_16
timestamp 1607194113
transform 1 0 21868 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_16
timestamp 1607194113
transform 1 0 21960 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_16
timestamp 1607194113
transform 1 0 21868 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_0
timestamp 1607194113
transform 1 0 2732 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_41
timestamp 1607194113
transform 1 0 1996 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_40
timestamp 1607194113
transform 1 0 1904 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_95
timestamp 1607194113
transform 1 0 3100 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_0
timestamp 1607194113
transform 1 0 2824 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_94
timestamp 1607194113
transform 1 0 4296 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_1
timestamp 1607194113
transform 1 0 4020 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_1
timestamp 1607194113
transform 1 0 3928 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_93
timestamp 1607194113
transform 1 0 5492 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_2
timestamp 1607194113
transform 1 0 5216 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_2
timestamp 1607194113
transform 1 0 5124 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_3
timestamp 1607194113
transform 1 0 6412 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_3
timestamp 1607194113
transform 1 0 6320 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_92
timestamp 1607194113
transform 1 0 6688 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_91
timestamp 1607194113
transform 1 0 7884 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_4
timestamp 1607194113
transform 1 0 7608 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_4
timestamp 1607194113
transform 1 0 7516 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_90
timestamp 1607194113
transform 1 0 9080 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_5
timestamp 1607194113
transform 1 0 8804 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_5
timestamp 1607194113
transform 1 0 8712 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_6
timestamp 1607194113
transform 1 0 10000 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_6
timestamp 1607194113
transform 1 0 9908 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_89
timestamp 1607194113
transform 1 0 10276 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_88
timestamp 1607194113
transform 1 0 11472 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_7
timestamp 1607194113
transform 1 0 11196 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_7
timestamp 1607194113
transform 1 0 11104 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_87
timestamp 1607194113
transform 1 0 12668 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_8
timestamp 1607194113
transform 1 0 12392 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_8
timestamp 1607194113
transform 1 0 12300 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_9
timestamp 1607194113
transform 1 0 13588 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_9
timestamp 1607194113
transform 1 0 13496 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_86
timestamp 1607194113
transform 1 0 13864 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_85
timestamp 1607194113
transform 1 0 15060 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_10
timestamp 1607194113
transform 1 0 14784 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_10
timestamp 1607194113
transform 1 0 14692 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_84
timestamp 1607194113
transform 1 0 16256 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_11
timestamp 1607194113
transform 1 0 15980 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_11
timestamp 1607194113
transform 1 0 15888 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_12
timestamp 1607194113
transform 1 0 17176 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_12
timestamp 1607194113
transform 1 0 17084 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_83
timestamp 1607194113
transform 1 0 17452 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_82
timestamp 1607194113
transform 1 0 18648 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_13
timestamp 1607194113
transform 1 0 18372 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_13
timestamp 1607194113
transform 1 0 18280 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_81
timestamp 1607194113
transform 1 0 19844 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_14
timestamp 1607194113
transform 1 0 19568 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_14
timestamp 1607194113
transform 1 0 19476 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_15
timestamp 1607194113
transform 1 0 20764 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_15
timestamp 1607194113
transform 1 0 20672 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_80
timestamp 1607194113
transform 1 0 21040 0 1 12352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap21_16
timestamp 1607194113
transform 1 0 21960 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_16
timestamp 1607194113
transform 1 0 21868 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_0
timestamp 1607194113
transform 1 0 2732 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_43
timestamp 1607194113
transform 1 0 1996 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_42
timestamp 1607194113
transform 1 0 1904 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_96
timestamp 1607194113
transform 1 0 3100 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_0
timestamp 1607194113
transform 1 0 2824 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_97
timestamp 1607194113
transform 1 0 4296 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_1
timestamp 1607194113
transform 1 0 4020 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_1
timestamp 1607194113
transform 1 0 3928 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_98
timestamp 1607194113
transform 1 0 5492 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_2
timestamp 1607194113
transform 1 0 5216 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_2
timestamp 1607194113
transform 1 0 5124 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_3
timestamp 1607194113
transform 1 0 6412 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_3
timestamp 1607194113
transform 1 0 6320 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_99
timestamp 1607194113
transform 1 0 6688 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_100
timestamp 1607194113
transform 1 0 7884 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_4
timestamp 1607194113
transform 1 0 7608 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_4
timestamp 1607194113
transform 1 0 7516 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_101
timestamp 1607194113
transform 1 0 9080 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_5
timestamp 1607194113
transform 1 0 8804 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_5
timestamp 1607194113
transform 1 0 8712 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_6
timestamp 1607194113
transform 1 0 10000 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_6
timestamp 1607194113
transform 1 0 9908 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_102
timestamp 1607194113
transform 1 0 10276 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_103
timestamp 1607194113
transform 1 0 11472 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_7
timestamp 1607194113
transform 1 0 11196 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_7
timestamp 1607194113
transform 1 0 11104 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_104
timestamp 1607194113
transform 1 0 12668 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_8
timestamp 1607194113
transform 1 0 12392 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_8
timestamp 1607194113
transform 1 0 12300 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_9
timestamp 1607194113
transform 1 0 13588 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_9
timestamp 1607194113
transform 1 0 13496 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_105
timestamp 1607194113
transform 1 0 13864 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_106
timestamp 1607194113
transform 1 0 15060 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_10
timestamp 1607194113
transform 1 0 14784 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_10
timestamp 1607194113
transform 1 0 14692 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_107
timestamp 1607194113
transform 1 0 16256 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_11
timestamp 1607194113
transform 1 0 15980 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_11
timestamp 1607194113
transform 1 0 15888 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_12
timestamp 1607194113
transform 1 0 17176 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_12
timestamp 1607194113
transform 1 0 17084 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_108
timestamp 1607194113
transform 1 0 17452 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_109
timestamp 1607194113
transform 1 0 18648 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_13
timestamp 1607194113
transform 1 0 18372 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_13
timestamp 1607194113
transform 1 0 18280 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_110
timestamp 1607194113
transform 1 0 19844 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_14
timestamp 1607194113
transform 1 0 19568 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_14
timestamp 1607194113
transform 1 0 19476 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_15
timestamp 1607194113
transform 1 0 20764 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_15
timestamp 1607194113
transform 1 0 20672 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_111
timestamp 1607194113
transform 1 0 21040 0 -1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap22_16
timestamp 1607194113
transform 1 0 21960 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_16
timestamp 1607194113
transform 1 0 21868 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_0
timestamp 1607194113
transform 1 0 2732 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_7
timestamp 1607194113
transform 1 0 1904 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_127
timestamp 1607194113
transform 1 0 3100 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_0
timestamp 1607194113
transform 1 0 2824 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_126
timestamp 1607194113
transform 1 0 4296 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_1
timestamp 1607194113
transform 1 0 4020 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_1
timestamp 1607194113
transform 1 0 3928 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_125
timestamp 1607194113
transform 1 0 5492 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_2
timestamp 1607194113
transform 1 0 5216 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_2
timestamp 1607194113
transform 1 0 5124 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_3
timestamp 1607194113
transform 1 0 6412 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_3
timestamp 1607194113
transform 1 0 6320 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_124
timestamp 1607194113
transform 1 0 6688 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_123
timestamp 1607194113
transform 1 0 7884 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_4
timestamp 1607194113
transform 1 0 7608 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_4
timestamp 1607194113
transform 1 0 7516 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_122
timestamp 1607194113
transform 1 0 9080 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_5
timestamp 1607194113
transform 1 0 8804 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_5
timestamp 1607194113
transform 1 0 8712 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_6
timestamp 1607194113
transform 1 0 10000 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_6
timestamp 1607194113
transform 1 0 9908 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_121
timestamp 1607194113
transform 1 0 10276 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_120
timestamp 1607194113
transform 1 0 11472 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_7
timestamp 1607194113
transform 1 0 11196 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_7
timestamp 1607194113
transform 1 0 11104 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_119
timestamp 1607194113
transform 1 0 12668 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_8
timestamp 1607194113
transform 1 0 12392 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_8
timestamp 1607194113
transform 1 0 12300 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_9
timestamp 1607194113
transform 1 0 13588 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_9
timestamp 1607194113
transform 1 0 13496 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_118
timestamp 1607194113
transform 1 0 13864 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_117
timestamp 1607194113
transform 1 0 15060 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_10
timestamp 1607194113
transform 1 0 14784 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_10
timestamp 1607194113
transform 1 0 14692 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_116
timestamp 1607194113
transform 1 0 16256 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_11
timestamp 1607194113
transform 1 0 15980 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_11
timestamp 1607194113
transform 1 0 15888 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_12
timestamp 1607194113
transform 1 0 17176 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_12
timestamp 1607194113
transform 1 0 17084 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_115
timestamp 1607194113
transform 1 0 17452 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_114
timestamp 1607194113
transform 1 0 18648 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_13
timestamp 1607194113
transform 1 0 18372 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_13
timestamp 1607194113
transform 1 0 18280 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_113
timestamp 1607194113
transform 1 0 19844 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_14
timestamp 1607194113
transform 1 0 19568 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_14
timestamp 1607194113
transform 1 0 19476 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_15
timestamp 1607194113
transform 1 0 20764 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_15
timestamp 1607194113
transform 1 0 20672 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_7_112
timestamp 1607194113
transform 1 0 21040 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap23_16
timestamp 1607194113
transform 1 0 21960 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_16
timestamp 1607194113
transform 1 0 21868 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_0
timestamp 1607194113
transform 1 0 2732 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_45
timestamp 1607194113
transform 1 0 1996 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_44
timestamp 1607194113
transform 1 0 1904 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_0
timestamp 1607194113
transform 1 0 3100 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_0
timestamp 1607194113
transform 1 0 2824 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_1
timestamp 1607194113
transform 1 0 4296 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_1
timestamp 1607194113
transform 1 0 4020 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_1
timestamp 1607194113
transform 1 0 3928 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_2
timestamp 1607194113
transform 1 0 5492 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_2
timestamp 1607194113
transform 1 0 5216 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_2
timestamp 1607194113
transform 1 0 5124 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_3
timestamp 1607194113
transform 1 0 6412 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_3
timestamp 1607194113
transform 1 0 6320 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_3
timestamp 1607194113
transform 1 0 6688 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_4
timestamp 1607194113
transform 1 0 7884 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_4
timestamp 1607194113
transform 1 0 7608 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_4
timestamp 1607194113
transform 1 0 7516 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_5
timestamp 1607194113
transform 1 0 9080 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_5
timestamp 1607194113
transform 1 0 8804 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_5
timestamp 1607194113
transform 1 0 8712 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_6
timestamp 1607194113
transform 1 0 10000 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_6
timestamp 1607194113
transform 1 0 9908 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_6
timestamp 1607194113
transform 1 0 10276 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_7
timestamp 1607194113
transform 1 0 11472 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_7
timestamp 1607194113
transform 1 0 11196 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_7
timestamp 1607194113
transform 1 0 11104 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_8
timestamp 1607194113
transform 1 0 12668 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_8
timestamp 1607194113
transform 1 0 12392 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_8
timestamp 1607194113
transform 1 0 12300 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_9
timestamp 1607194113
transform 1 0 13588 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_9
timestamp 1607194113
transform 1 0 13496 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_9
timestamp 1607194113
transform 1 0 13864 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_10
timestamp 1607194113
transform 1 0 15060 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_10
timestamp 1607194113
transform 1 0 14784 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_10
timestamp 1607194113
transform 1 0 14692 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_11
timestamp 1607194113
transform 1 0 16256 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_11
timestamp 1607194113
transform 1 0 15980 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_11
timestamp 1607194113
transform 1 0 15888 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_12
timestamp 1607194113
transform 1 0 17176 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_12
timestamp 1607194113
transform 1 0 17084 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_12
timestamp 1607194113
transform 1 0 17452 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_13
timestamp 1607194113
transform 1 0 18648 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_13
timestamp 1607194113
transform 1 0 18372 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_13
timestamp 1607194113
transform 1 0 18280 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_14
timestamp 1607194113
transform 1 0 19844 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_14
timestamp 1607194113
transform 1 0 19568 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_14
timestamp 1607194113
transform 1 0 19476 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_15
timestamp 1607194113
transform 1 0 20764 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_15
timestamp 1607194113
transform 1 0 20672 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_15
timestamp 1607194113
transform 1 0 21040 0 -1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap24_16
timestamp 1607194113
transform 1 0 21960 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_16
timestamp 1607194113
transform 1 0 21868 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_0
timestamp 1607194113
transform 1 0 2732 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_47
timestamp 1607194113
transform 1 0 1996 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_46
timestamp 1607194113
transform 1 0 1904 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_31
timestamp 1607194113
transform 1 0 3100 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_0
timestamp 1607194113
transform 1 0 2824 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_30
timestamp 1607194113
transform 1 0 4296 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_1
timestamp 1607194113
transform 1 0 4020 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_1
timestamp 1607194113
transform 1 0 3928 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_29
timestamp 1607194113
transform 1 0 5492 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_2
timestamp 1607194113
transform 1 0 5216 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_2
timestamp 1607194113
transform 1 0 5124 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_3
timestamp 1607194113
transform 1 0 6412 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_3
timestamp 1607194113
transform 1 0 6320 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_28
timestamp 1607194113
transform 1 0 6688 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_27
timestamp 1607194113
transform 1 0 7884 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_4
timestamp 1607194113
transform 1 0 7608 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_4
timestamp 1607194113
transform 1 0 7516 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_26
timestamp 1607194113
transform 1 0 9080 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_5
timestamp 1607194113
transform 1 0 8804 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_5
timestamp 1607194113
transform 1 0 8712 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_6
timestamp 1607194113
transform 1 0 10000 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_6
timestamp 1607194113
transform 1 0 9908 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_25
timestamp 1607194113
transform 1 0 10276 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_24
timestamp 1607194113
transform 1 0 11472 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_7
timestamp 1607194113
transform 1 0 11196 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_7
timestamp 1607194113
transform 1 0 11104 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_23
timestamp 1607194113
transform 1 0 12668 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_8
timestamp 1607194113
transform 1 0 12392 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_8
timestamp 1607194113
transform 1 0 12300 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_9
timestamp 1607194113
transform 1 0 13588 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_9
timestamp 1607194113
transform 1 0 13496 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_22
timestamp 1607194113
transform 1 0 13864 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_21
timestamp 1607194113
transform 1 0 15060 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_10
timestamp 1607194113
transform 1 0 14784 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_10
timestamp 1607194113
transform 1 0 14692 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_20
timestamp 1607194113
transform 1 0 16256 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_11
timestamp 1607194113
transform 1 0 15980 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_11
timestamp 1607194113
transform 1 0 15888 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_12
timestamp 1607194113
transform 1 0 17176 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_12
timestamp 1607194113
transform 1 0 17084 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_19
timestamp 1607194113
transform 1 0 17452 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_18
timestamp 1607194113
transform 1 0 18648 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_13
timestamp 1607194113
transform 1 0 18372 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_13
timestamp 1607194113
transform 1 0 18280 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_17
timestamp 1607194113
transform 1 0 19844 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_14
timestamp 1607194113
transform 1 0 19568 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_14
timestamp 1607194113
transform 1 0 19476 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_15
timestamp 1607194113
transform 1 0 20764 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_15
timestamp 1607194113
transform 1 0 20672 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_16
timestamp 1607194113
transform 1 0 21040 0 1 14528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap25_16
timestamp 1607194113
transform 1 0 21960 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_16
timestamp 1607194113
transform 1 0 21868 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_0
timestamp 1607194113
transform 1 0 2732 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_6
timestamp 1607194113
transform 1 0 1904 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_0
timestamp 1607194113
transform 1 0 2732 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_49
timestamp 1607194113
transform 1 0 1996 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_48
timestamp 1607194113
transform 1 0 1904 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_63
timestamp 1607194113
transform 1 0 3100 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_0
timestamp 1607194113
transform 1 0 2824 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_32
timestamp 1607194113
transform 1 0 3100 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_0
timestamp 1607194113
transform 1 0 2824 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_62
timestamp 1607194113
transform 1 0 4296 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_1
timestamp 1607194113
transform 1 0 4020 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_1
timestamp 1607194113
transform 1 0 3928 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_33
timestamp 1607194113
transform 1 0 4296 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_1
timestamp 1607194113
transform 1 0 4020 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_1
timestamp 1607194113
transform 1 0 3928 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_61
timestamp 1607194113
transform 1 0 5492 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_2
timestamp 1607194113
transform 1 0 5216 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_2
timestamp 1607194113
transform 1 0 5124 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_34
timestamp 1607194113
transform 1 0 5492 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_2
timestamp 1607194113
transform 1 0 5216 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_2
timestamp 1607194113
transform 1 0 5124 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_3
timestamp 1607194113
transform 1 0 6412 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_3
timestamp 1607194113
transform 1 0 6320 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_3
timestamp 1607194113
transform 1 0 6412 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_3
timestamp 1607194113
transform 1 0 6320 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_60
timestamp 1607194113
transform 1 0 6688 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_35
timestamp 1607194113
transform 1 0 6688 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_59
timestamp 1607194113
transform 1 0 7884 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_4
timestamp 1607194113
transform 1 0 7608 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_4
timestamp 1607194113
transform 1 0 7516 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_36
timestamp 1607194113
transform 1 0 7884 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_4
timestamp 1607194113
transform 1 0 7608 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_4
timestamp 1607194113
transform 1 0 7516 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_58
timestamp 1607194113
transform 1 0 9080 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_5
timestamp 1607194113
transform 1 0 8804 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_5
timestamp 1607194113
transform 1 0 8712 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_37
timestamp 1607194113
transform 1 0 9080 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_5
timestamp 1607194113
transform 1 0 8804 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_5
timestamp 1607194113
transform 1 0 8712 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_6
timestamp 1607194113
transform 1 0 10000 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_6
timestamp 1607194113
transform 1 0 9908 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_6
timestamp 1607194113
transform 1 0 10000 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_6
timestamp 1607194113
transform 1 0 9908 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_57
timestamp 1607194113
transform 1 0 10276 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_38
timestamp 1607194113
transform 1 0 10276 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_56
timestamp 1607194113
transform 1 0 11472 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_7
timestamp 1607194113
transform 1 0 11196 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_7
timestamp 1607194113
transform 1 0 11104 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_39
timestamp 1607194113
transform 1 0 11472 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_7
timestamp 1607194113
transform 1 0 11196 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_7
timestamp 1607194113
transform 1 0 11104 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_55
timestamp 1607194113
transform 1 0 12668 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_8
timestamp 1607194113
transform 1 0 12392 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_8
timestamp 1607194113
transform 1 0 12300 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_40
timestamp 1607194113
transform 1 0 12668 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_8
timestamp 1607194113
transform 1 0 12392 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_8
timestamp 1607194113
transform 1 0 12300 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_9
timestamp 1607194113
transform 1 0 13588 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_9
timestamp 1607194113
transform 1 0 13496 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_9
timestamp 1607194113
transform 1 0 13588 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_9
timestamp 1607194113
transform 1 0 13496 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_54
timestamp 1607194113
transform 1 0 13864 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_41
timestamp 1607194113
transform 1 0 13864 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_53
timestamp 1607194113
transform 1 0 15060 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_10
timestamp 1607194113
transform 1 0 14784 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_10
timestamp 1607194113
transform 1 0 14692 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_42
timestamp 1607194113
transform 1 0 15060 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_10
timestamp 1607194113
transform 1 0 14784 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_10
timestamp 1607194113
transform 1 0 14692 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_52
timestamp 1607194113
transform 1 0 16256 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_11
timestamp 1607194113
transform 1 0 15980 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_11
timestamp 1607194113
transform 1 0 15888 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_43
timestamp 1607194113
transform 1 0 16256 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_11
timestamp 1607194113
transform 1 0 15980 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_11
timestamp 1607194113
transform 1 0 15888 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_12
timestamp 1607194113
transform 1 0 17176 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_12
timestamp 1607194113
transform 1 0 17084 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_12
timestamp 1607194113
transform 1 0 17176 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_12
timestamp 1607194113
transform 1 0 17084 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_51
timestamp 1607194113
transform 1 0 17452 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_44
timestamp 1607194113
transform 1 0 17452 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_50
timestamp 1607194113
transform 1 0 18648 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_13
timestamp 1607194113
transform 1 0 18372 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_13
timestamp 1607194113
transform 1 0 18280 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_45
timestamp 1607194113
transform 1 0 18648 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_13
timestamp 1607194113
transform 1 0 18372 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_13
timestamp 1607194113
transform 1 0 18280 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_49
timestamp 1607194113
transform 1 0 19844 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_14
timestamp 1607194113
transform 1 0 19568 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_14
timestamp 1607194113
transform 1 0 19476 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_46
timestamp 1607194113
transform 1 0 19844 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap26_14
timestamp 1607194113
transform 1 0 19568 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_14
timestamp 1607194113
transform 1 0 19476 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_15
timestamp 1607194113
transform 1 0 20764 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_15
timestamp 1607194113
transform 1 0 20672 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_15
timestamp 1607194113
transform 1 0 20764 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_15
timestamp 1607194113
transform 1 0 20672 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_48
timestamp 1607194113
transform 1 0 21040 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_6_47
timestamp 1607194113
transform 1 0 21040 0 -1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap27_16
timestamp 1607194113
transform 1 0 21960 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_16
timestamp 1607194113
transform 1 0 21868 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_16
timestamp 1607194113
transform 1 0 21960 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_16
timestamp 1607194113
transform 1 0 21868 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_0
timestamp 1607194113
transform 1 0 2732 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_51
timestamp 1607194113
transform 1 0 1996 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_50
timestamp 1607194113
transform 1 0 1904 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_0
timestamp 1607194113
transform 1 0 3100 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_0
timestamp 1607194113
transform 1 0 2824 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_1
timestamp 1607194113
transform 1 0 4296 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_1
timestamp 1607194113
transform 1 0 4020 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_1
timestamp 1607194113
transform 1 0 3928 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_2
timestamp 1607194113
transform 1 0 5492 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_2
timestamp 1607194113
transform 1 0 5216 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_2
timestamp 1607194113
transform 1 0 5124 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_3
timestamp 1607194113
transform 1 0 6412 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_3
timestamp 1607194113
transform 1 0 6320 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_3
timestamp 1607194113
transform 1 0 6688 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_4
timestamp 1607194113
transform 1 0 7884 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_4
timestamp 1607194113
transform 1 0 7608 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_4
timestamp 1607194113
transform 1 0 7516 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_5
timestamp 1607194113
transform 1 0 9080 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_5
timestamp 1607194113
transform 1 0 8804 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_5
timestamp 1607194113
transform 1 0 8712 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_6
timestamp 1607194113
transform 1 0 10000 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_6
timestamp 1607194113
transform 1 0 9908 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_6
timestamp 1607194113
transform 1 0 10276 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_7
timestamp 1607194113
transform 1 0 11472 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_7
timestamp 1607194113
transform 1 0 11196 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_7
timestamp 1607194113
transform 1 0 11104 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_8
timestamp 1607194113
transform 1 0 12668 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_8
timestamp 1607194113
transform 1 0 12392 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_8
timestamp 1607194113
transform 1 0 12300 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_9
timestamp 1607194113
transform 1 0 13588 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_9
timestamp 1607194113
transform 1 0 13496 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_9
timestamp 1607194113
transform 1 0 13864 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_10
timestamp 1607194113
transform 1 0 15060 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_10
timestamp 1607194113
transform 1 0 14784 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_10
timestamp 1607194113
transform 1 0 14692 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_11
timestamp 1607194113
transform 1 0 16256 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_11
timestamp 1607194113
transform 1 0 15980 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_11
timestamp 1607194113
transform 1 0 15888 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_12
timestamp 1607194113
transform 1 0 17176 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_12
timestamp 1607194113
transform 1 0 17084 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_12
timestamp 1607194113
transform 1 0 17452 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_13
timestamp 1607194113
transform 1 0 18648 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_13
timestamp 1607194113
transform 1 0 18372 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_13
timestamp 1607194113
transform 1 0 18280 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_14
timestamp 1607194113
transform 1 0 19844 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_14
timestamp 1607194113
transform 1 0 19568 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_14
timestamp 1607194113
transform 1 0 19476 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_15
timestamp 1607194113
transform 1 0 20764 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_15
timestamp 1607194113
transform 1 0 20672 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_15
timestamp 1607194113
transform 1 0 21040 0 -1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap28_16
timestamp 1607194113
transform 1 0 21960 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_16
timestamp 1607194113
transform 1 0 21868 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_0
timestamp 1607194113
transform 1 0 2732 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_5
timestamp 1607194113
transform 1 0 1904 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_31
timestamp 1607194113
transform 1 0 3100 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_0
timestamp 1607194113
transform 1 0 2824 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_30
timestamp 1607194113
transform 1 0 4296 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_1
timestamp 1607194113
transform 1 0 4020 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_1
timestamp 1607194113
transform 1 0 3928 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_29
timestamp 1607194113
transform 1 0 5492 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_2
timestamp 1607194113
transform 1 0 5216 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_2
timestamp 1607194113
transform 1 0 5124 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_3
timestamp 1607194113
transform 1 0 6412 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_3
timestamp 1607194113
transform 1 0 6320 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_28
timestamp 1607194113
transform 1 0 6688 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_27
timestamp 1607194113
transform 1 0 7884 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_4
timestamp 1607194113
transform 1 0 7608 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_4
timestamp 1607194113
transform 1 0 7516 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_26
timestamp 1607194113
transform 1 0 9080 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_5
timestamp 1607194113
transform 1 0 8804 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_5
timestamp 1607194113
transform 1 0 8712 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_6
timestamp 1607194113
transform 1 0 10000 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_6
timestamp 1607194113
transform 1 0 9908 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_25
timestamp 1607194113
transform 1 0 10276 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_24
timestamp 1607194113
transform 1 0 11472 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_7
timestamp 1607194113
transform 1 0 11196 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_7
timestamp 1607194113
transform 1 0 11104 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_23
timestamp 1607194113
transform 1 0 12668 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_8
timestamp 1607194113
transform 1 0 12392 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_8
timestamp 1607194113
transform 1 0 12300 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_9
timestamp 1607194113
transform 1 0 13588 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_9
timestamp 1607194113
transform 1 0 13496 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_22
timestamp 1607194113
transform 1 0 13864 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_21
timestamp 1607194113
transform 1 0 15060 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_10
timestamp 1607194113
transform 1 0 14784 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_10
timestamp 1607194113
transform 1 0 14692 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_20
timestamp 1607194113
transform 1 0 16256 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_11
timestamp 1607194113
transform 1 0 15980 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_11
timestamp 1607194113
transform 1 0 15888 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_12
timestamp 1607194113
transform 1 0 17176 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_12
timestamp 1607194113
transform 1 0 17084 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_19
timestamp 1607194113
transform 1 0 17452 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_18
timestamp 1607194113
transform 1 0 18648 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_13
timestamp 1607194113
transform 1 0 18372 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_13
timestamp 1607194113
transform 1 0 18280 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_17
timestamp 1607194113
transform 1 0 19844 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_14
timestamp 1607194113
transform 1 0 19568 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_14
timestamp 1607194113
transform 1 0 19476 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_15
timestamp 1607194113
transform 1 0 20764 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_15
timestamp 1607194113
transform 1 0 20672 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_5_16
timestamp 1607194113
transform 1 0 21040 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap29_16
timestamp 1607194113
transform 1 0 21960 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_16
timestamp 1607194113
transform 1 0 21868 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_0
timestamp 1607194113
transform 1 0 2732 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_53
timestamp 1607194113
transform 1 0 1996 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_52
timestamp 1607194113
transform 1 0 1904 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_0
timestamp 1607194113
transform 1 0 3100 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap30_0
timestamp 1607194113
transform 1 0 2824 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_1
timestamp 1607194113
transform 1 0 4296 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap30_1
timestamp 1607194113
transform 1 0 4020 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_1
timestamp 1607194113
transform 1 0 3928 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_2
timestamp 1607194113
transform 1 0 5492 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap30_2
timestamp 1607194113
transform 1 0 5216 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_2
timestamp 1607194113
transform 1 0 5124 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap30_3
timestamp 1607194113
transform 1 0 6412 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_3
timestamp 1607194113
transform 1 0 6320 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_3
timestamp 1607194113
transform 1 0 6688 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_4
timestamp 1607194113
transform 1 0 7884 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap30_4
timestamp 1607194113
transform 1 0 7608 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_4
timestamp 1607194113
transform 1 0 7516 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_5
timestamp 1607194113
transform 1 0 9080 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap30_5
timestamp 1607194113
transform 1 0 8804 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_5
timestamp 1607194113
transform 1 0 8712 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap30_6
timestamp 1607194113
transform 1 0 10000 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_6
timestamp 1607194113
transform 1 0 9908 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_6
timestamp 1607194113
transform 1 0 10276 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_7
timestamp 1607194113
transform 1 0 11472 0 -1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap30_7
timestamp 1607194113
transform 1 0 11196 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_7
timestamp 1607194113
transform 1 0 11104 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_61
timestamp 1607194113
transform 1 0 12760 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_60
timestamp 1607194113
transform 1 0 12668 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap30_8
timestamp 1607194113
transform 1 0 12392 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_8
timestamp 1607194113
transform 1 0 12300 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_63
timestamp 1607194113
transform 1 0 13588 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_62
timestamp 1607194113
transform 1 0 13496 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_65
timestamp 1607194113
transform 1 0 14416 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_64
timestamp 1607194113
transform 1 0 14324 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_67
timestamp 1607194113
transform 1 0 15244 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_66
timestamp 1607194113
transform 1 0 15152 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_69
timestamp 1607194113
transform 1 0 16072 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_68
timestamp 1607194113
transform 1 0 15980 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_71
timestamp 1607194113
transform 1 0 16900 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_70
timestamp 1607194113
transform 1 0 16808 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_73
timestamp 1607194113
transform 1 0 17728 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_72
timestamp 1607194113
transform 1 0 17636 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_75
timestamp 1607194113
transform 1 0 18556 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_74
timestamp 1607194113
transform 1 0 18464 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_77
timestamp 1607194113
transform 1 0 19384 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_76
timestamp 1607194113
transform 1 0 19292 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_79
timestamp 1607194113
transform 1 0 20212 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_78
timestamp 1607194113
transform 1 0 20120 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 21776 0 -1 17792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILL_81
timestamp 1607194113
transform 1 0 21040 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_80
timestamp 1607194113
transform 1 0 20948 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 22144 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_0
timestamp 1607194113
transform 1 0 2732 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_4
timestamp 1607194113
transform 1 0 1904 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_15
timestamp 1607194113
transform 1 0 3100 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap31_0
timestamp 1607194113
transform 1 0 2824 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_14
timestamp 1607194113
transform 1 0 4296 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap31_1
timestamp 1607194113
transform 1 0 4020 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_1
timestamp 1607194113
transform 1 0 3928 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_13
timestamp 1607194113
transform 1 0 5492 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap31_2
timestamp 1607194113
transform 1 0 5216 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_2
timestamp 1607194113
transform 1 0 5124 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap31_3
timestamp 1607194113
transform 1 0 6412 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_3
timestamp 1607194113
transform 1 0 6320 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_12
timestamp 1607194113
transform 1 0 6688 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_11
timestamp 1607194113
transform 1 0 7884 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap31_4
timestamp 1607194113
transform 1 0 7608 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_4
timestamp 1607194113
transform 1 0 7516 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_10
timestamp 1607194113
transform 1 0 9080 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap31_5
timestamp 1607194113
transform 1 0 8804 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_5
timestamp 1607194113
transform 1 0 8712 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap31_6
timestamp 1607194113
transform 1 0 10000 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_6
timestamp 1607194113
transform 1 0 9908 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_9
timestamp 1607194113
transform 1 0 10276 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_4_8
timestamp 1607194113
transform 1 0 11472 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap31_7
timestamp 1607194113
transform 1 0 11196 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_7
timestamp 1607194113
transform 1 0 11104 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_85
timestamp 1607194113
transform 1 0 12760 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_84
timestamp 1607194113
transform 1 0 12668 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap31_8
timestamp 1607194113
transform 1 0 12392 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_8
timestamp 1607194113
transform 1 0 12300 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_87
timestamp 1607194113
transform 1 0 13588 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_86
timestamp 1607194113
transform 1 0 13496 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_89
timestamp 1607194113
transform 1 0 14416 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_88
timestamp 1607194113
transform 1 0 14324 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_91
timestamp 1607194113
transform 1 0 15244 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_90
timestamp 1607194113
transform 1 0 15152 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_93
timestamp 1607194113
transform 1 0 16072 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_92
timestamp 1607194113
transform 1 0 15980 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_95
timestamp 1607194113
transform 1 0 16900 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_94
timestamp 1607194113
transform 1 0 16808 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_97
timestamp 1607194113
transform 1 0 17728 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_96
timestamp 1607194113
transform 1 0 17636 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_99
timestamp 1607194113
transform 1 0 18556 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_98
timestamp 1607194113
transform 1 0 18464 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_101
timestamp 1607194113
transform 1 0 19384 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_100
timestamp 1607194113
transform 1 0 19292 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_103
timestamp 1607194113
transform 1 0 20212 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_102
timestamp 1607194113
transform 1 0 20120 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_106
timestamp 1607194113
transform 1 0 21776 0 1 17792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILL_105
timestamp 1607194113
transform 1 0 21040 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_104
timestamp 1607194113
transform 1 0 20948 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_107
timestamp 1607194113
transform 1 0 22144 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_0
timestamp 1607194113
transform 1 0 2732 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_55
timestamp 1607194113
transform 1 0 1996 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_54
timestamp 1607194113
transform 1 0 1904 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_0
timestamp 1607194113
transform 1 0 3100 0 -1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap32_0
timestamp 1607194113
transform 1 0 2824 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_1
timestamp 1607194113
transform 1 0 4296 0 -1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap32_1
timestamp 1607194113
transform 1 0 4020 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_1
timestamp 1607194113
transform 1 0 3928 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_2
timestamp 1607194113
transform 1 0 5492 0 -1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap32_2
timestamp 1607194113
transform 1 0 5216 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_2
timestamp 1607194113
transform 1 0 5124 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap32_3
timestamp 1607194113
transform 1 0 6412 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_3
timestamp 1607194113
transform 1 0 6320 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_3
timestamp 1607194113
transform 1 0 6688 0 -1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_8  FILL_109
timestamp 1607194113
transform 1 0 7976 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_108
timestamp 1607194113
transform 1 0 7884 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap32_4
timestamp 1607194113
transform 1 0 7608 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_4
timestamp 1607194113
transform 1 0 7516 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_111
timestamp 1607194113
transform 1 0 8804 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_110
timestamp 1607194113
transform 1 0 8712 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_113
timestamp 1607194113
transform 1 0 9632 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_112
timestamp 1607194113
transform 1 0 9540 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_115
timestamp 1607194113
transform 1 0 10460 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_114
timestamp 1607194113
transform 1 0 10368 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_117
timestamp 1607194113
transform 1 0 11288 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_116
timestamp 1607194113
transform 1 0 11196 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_119
timestamp 1607194113
transform 1 0 12116 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_118
timestamp 1607194113
transform 1 0 12024 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_121
timestamp 1607194113
transform 1 0 12944 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_120
timestamp 1607194113
transform 1 0 12852 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_124
timestamp 1607194113
transform 1 0 14508 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_123
timestamp 1607194113
transform 1 0 13772 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_122
timestamp 1607194113
transform 1 0 13680 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_127
timestamp 1607194113
transform 1 0 15428 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_126
timestamp 1607194113
transform 1 0 15336 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_125
timestamp 1607194113
transform 1 0 14600 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_129
timestamp 1607194113
transform 1 0 16256 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_128
timestamp 1607194113
transform 1 0 16164 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_131
timestamp 1607194113
transform 1 0 17084 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_130
timestamp 1607194113
transform 1 0 16992 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_133
timestamp 1607194113
transform 1 0 17912 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_132
timestamp 1607194113
transform 1 0 17820 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_135
timestamp 1607194113
transform 1 0 18740 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_134
timestamp 1607194113
transform 1 0 18648 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_137
timestamp 1607194113
transform 1 0 19568 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_136
timestamp 1607194113
transform 1 0 19476 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_139
timestamp 1607194113
transform 1 0 20396 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_138
timestamp 1607194113
transform 1 0 20304 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_141
timestamp 1607194113
transform 1 0 21224 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_140
timestamp 1607194113
transform 1 0 21132 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_143
timestamp 1607194113
transform 1 0 22144 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_142 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 21960 0 -1 18880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap34_0
timestamp 1607194113
transform 1 0 2732 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_57
timestamp 1607194113
transform 1 0 1996 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_56
timestamp 1607194113
transform 1 0 1904 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_0
timestamp 1607194113
transform 1 0 2732 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_3
timestamp 1607194113
transform 1 0 1904 0 1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_2_0
timestamp 1607194113
transform 1 0 3100 0 -1 19968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap34_0
timestamp 1607194113
transform 1 0 2824 0 -1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_7
timestamp 1607194113
transform 1 0 3100 0 1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap33_0
timestamp 1607194113
transform 1 0 2824 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_2_1
timestamp 1607194113
transform 1 0 4296 0 -1 19968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap34_1
timestamp 1607194113
transform 1 0 4020 0 -1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap34_1
timestamp 1607194113
transform 1 0 3928 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_6
timestamp 1607194113
transform 1 0 4296 0 1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap33_1
timestamp 1607194113
transform 1 0 4020 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_1
timestamp 1607194113
transform 1 0 3928 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_180
timestamp 1607194113
transform 1 0 5492 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap34_2
timestamp 1607194113
transform 1 0 5216 0 -1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap34_2
timestamp 1607194113
transform 1 0 5124 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_5
timestamp 1607194113
transform 1 0 5492 0 1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap33_2
timestamp 1607194113
transform 1 0 5216 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_2
timestamp 1607194113
transform 1 0 5124 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_183
timestamp 1607194113
transform 1 0 6412 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_182
timestamp 1607194113
transform 1 0 6320 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_181
timestamp 1607194113
transform 1 0 5584 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap33_3
timestamp 1607194113
transform 1 0 6412 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_3
timestamp 1607194113
transform 1 0 6320 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_185
timestamp 1607194113
transform 1 0 7240 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_184
timestamp 1607194113
transform 1 0 7148 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_3_4
timestamp 1607194113
transform 1 0 6688 0 1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_8  FILL_187
timestamp 1607194113
transform 1 0 8068 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_186
timestamp 1607194113
transform 1 0 7976 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_145
timestamp 1607194113
transform 1 0 7976 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_144
timestamp 1607194113
transform 1 0 7884 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap33_4
timestamp 1607194113
transform 1 0 7608 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_4
timestamp 1607194113
transform 1 0 7516 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_189
timestamp 1607194113
transform 1 0 8896 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_188
timestamp 1607194113
transform 1 0 8804 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_147
timestamp 1607194113
transform 1 0 8804 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_146
timestamp 1607194113
transform 1 0 8712 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_191
timestamp 1607194113
transform 1 0 9724 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_190
timestamp 1607194113
transform 1 0 9632 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_149
timestamp 1607194113
transform 1 0 9632 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_148
timestamp 1607194113
transform 1 0 9540 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_193
timestamp 1607194113
transform 1 0 10552 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_192
timestamp 1607194113
transform 1 0 10460 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_151
timestamp 1607194113
transform 1 0 10460 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_150
timestamp 1607194113
transform 1 0 10368 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_195
timestamp 1607194113
transform 1 0 11380 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_194
timestamp 1607194113
transform 1 0 11288 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_153
timestamp 1607194113
transform 1 0 11288 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_152
timestamp 1607194113
transform 1 0 11196 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_197
timestamp 1607194113
transform 1 0 12208 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_196
timestamp 1607194113
transform 1 0 12116 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_155
timestamp 1607194113
transform 1 0 12116 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_154
timestamp 1607194113
transform 1 0 12024 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_199
timestamp 1607194113
transform 1 0 13036 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_198
timestamp 1607194113
transform 1 0 12944 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_157
timestamp 1607194113
transform 1 0 12944 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_156
timestamp 1607194113
transform 1 0 12852 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_201
timestamp 1607194113
transform 1 0 13864 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_200
timestamp 1607194113
transform 1 0 13772 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_160
timestamp 1607194113
transform 1 0 14508 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_159
timestamp 1607194113
transform 1 0 13772 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_158
timestamp 1607194113
transform 1 0 13680 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_204
timestamp 1607194113
transform 1 0 15428 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_203
timestamp 1607194113
transform 1 0 14692 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_202
timestamp 1607194113
transform 1 0 14600 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_163
timestamp 1607194113
transform 1 0 15428 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_162
timestamp 1607194113
transform 1 0 15336 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_161
timestamp 1607194113
transform 1 0 14600 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_207
timestamp 1607194113
transform 1 0 16348 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_206
timestamp 1607194113
transform 1 0 16256 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_205
timestamp 1607194113
transform 1 0 15520 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_165
timestamp 1607194113
transform 1 0 16256 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_164
timestamp 1607194113
transform 1 0 16164 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_209
timestamp 1607194113
transform 1 0 17176 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_208
timestamp 1607194113
transform 1 0 17084 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_167
timestamp 1607194113
transform 1 0 17084 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_166
timestamp 1607194113
transform 1 0 16992 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_211
timestamp 1607194113
transform 1 0 18004 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_210
timestamp 1607194113
transform 1 0 17912 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_169
timestamp 1607194113
transform 1 0 17912 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_168
timestamp 1607194113
transform 1 0 17820 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_213
timestamp 1607194113
transform 1 0 18832 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_212
timestamp 1607194113
transform 1 0 18740 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_171
timestamp 1607194113
transform 1 0 18740 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_170
timestamp 1607194113
transform 1 0 18648 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_215
timestamp 1607194113
transform 1 0 19660 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_214
timestamp 1607194113
transform 1 0 19568 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_173
timestamp 1607194113
transform 1 0 19568 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_172
timestamp 1607194113
transform 1 0 19476 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_217
timestamp 1607194113
transform 1 0 20488 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_216
timestamp 1607194113
transform 1 0 20396 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_175
timestamp 1607194113
transform 1 0 20396 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_174
timestamp 1607194113
transform 1 0 20304 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_219
timestamp 1607194113
transform 1 0 21316 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_218
timestamp 1607194113
transform 1 0 21224 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_177
timestamp 1607194113
transform 1 0 21224 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_176
timestamp 1607194113
transform 1 0 21132 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_220
timestamp 1607194113
transform 1 0 22052 0 -1 19968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_179
timestamp 1607194113
transform 1 0 22144 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_178
timestamp 1607194113
transform 1 0 21960 0 1 18880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap35_0
timestamp 1607194113
transform 1 0 2732 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_2
timestamp 1607194113
transform 1 0 1904 0 1 19968
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_2_3
timestamp 1607194113
transform 1 0 3100 0 1 19968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap35_0
timestamp 1607194113
transform 1 0 2824 0 1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_2_2
timestamp 1607194113
transform 1 0 4296 0 1 19968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap35_1
timestamp 1607194113
transform 1 0 4020 0 1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap35_1
timestamp 1607194113
transform 1 0 3928 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_221
timestamp 1607194113
transform 1 0 5492 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap35_2
timestamp 1607194113
transform 1 0 5216 0 1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap35_2
timestamp 1607194113
transform 1 0 5124 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_224
timestamp 1607194113
transform 1 0 6412 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_223
timestamp 1607194113
transform 1 0 6320 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_222
timestamp 1607194113
transform 1 0 5584 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_226
timestamp 1607194113
transform 1 0 7240 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_225
timestamp 1607194113
transform 1 0 7148 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_228
timestamp 1607194113
transform 1 0 8068 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_227
timestamp 1607194113
transform 1 0 7976 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_230
timestamp 1607194113
transform 1 0 8896 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_229
timestamp 1607194113
transform 1 0 8804 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_232
timestamp 1607194113
transform 1 0 9724 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_231
timestamp 1607194113
transform 1 0 9632 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_234
timestamp 1607194113
transform 1 0 10552 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_233
timestamp 1607194113
transform 1 0 10460 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_236
timestamp 1607194113
transform 1 0 11380 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_235
timestamp 1607194113
transform 1 0 11288 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_238
timestamp 1607194113
transform 1 0 12208 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_237
timestamp 1607194113
transform 1 0 12116 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_240
timestamp 1607194113
transform 1 0 13036 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_239
timestamp 1607194113
transform 1 0 12944 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_242
timestamp 1607194113
transform 1 0 13864 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_241
timestamp 1607194113
transform 1 0 13772 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_245
timestamp 1607194113
transform 1 0 15428 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_244
timestamp 1607194113
transform 1 0 14692 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_243
timestamp 1607194113
transform 1 0 14600 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_248
timestamp 1607194113
transform 1 0 16348 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_247
timestamp 1607194113
transform 1 0 16256 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_246
timestamp 1607194113
transform 1 0 15520 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_250
timestamp 1607194113
transform 1 0 17176 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_249
timestamp 1607194113
transform 1 0 17084 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_252
timestamp 1607194113
transform 1 0 18004 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_251
timestamp 1607194113
transform 1 0 17912 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_254
timestamp 1607194113
transform 1 0 18832 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_253
timestamp 1607194113
transform 1 0 18740 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_256
timestamp 1607194113
transform 1 0 19660 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_255
timestamp 1607194113
transform 1 0 19568 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_258
timestamp 1607194113
transform 1 0 20488 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_257
timestamp 1607194113
transform 1 0 20396 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_260
timestamp 1607194113
transform 1 0 21316 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_259
timestamp 1607194113
transform 1 0 21224 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_261
timestamp 1607194113
transform 1 0 22052 0 1 19968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap36_0
timestamp 1607194113
transform 1 0 2732 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_59
timestamp 1607194113
transform 1 0 1996 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_58
timestamp 1607194113
transform 1 0 1904 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_1_0
timestamp 1607194113
transform 1 0 3100 0 -1 21056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap36_0
timestamp 1607194113
transform 1 0 2824 0 -1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_263
timestamp 1607194113
transform 1 0 4388 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_262
timestamp 1607194113
transform 1 0 4296 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap36_1
timestamp 1607194113
transform 1 0 4020 0 -1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap36_1
timestamp 1607194113
transform 1 0 3928 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_265
timestamp 1607194113
transform 1 0 5216 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_264
timestamp 1607194113
transform 1 0 5124 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_267
timestamp 1607194113
transform 1 0 6044 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_266
timestamp 1607194113
transform 1 0 5952 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_269
timestamp 1607194113
transform 1 0 6872 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_268
timestamp 1607194113
transform 1 0 6780 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_271
timestamp 1607194113
transform 1 0 7700 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_270
timestamp 1607194113
transform 1 0 7608 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_273
timestamp 1607194113
transform 1 0 8528 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_272
timestamp 1607194113
transform 1 0 8436 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_275
timestamp 1607194113
transform 1 0 9356 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_274
timestamp 1607194113
transform 1 0 9264 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_278
timestamp 1607194113
transform 1 0 10920 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_277
timestamp 1607194113
transform 1 0 10184 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_276
timestamp 1607194113
transform 1 0 10092 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_281
timestamp 1607194113
transform 1 0 11840 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_280
timestamp 1607194113
transform 1 0 11748 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_279
timestamp 1607194113
transform 1 0 11012 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_283
timestamp 1607194113
transform 1 0 12668 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_282
timestamp 1607194113
transform 1 0 12576 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_285
timestamp 1607194113
transform 1 0 13496 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_284
timestamp 1607194113
transform 1 0 13404 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_287
timestamp 1607194113
transform 1 0 14324 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_286
timestamp 1607194113
transform 1 0 14232 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_289
timestamp 1607194113
transform 1 0 15152 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_288
timestamp 1607194113
transform 1 0 15060 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_291
timestamp 1607194113
transform 1 0 15980 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_290
timestamp 1607194113
transform 1 0 15888 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_293
timestamp 1607194113
transform 1 0 16808 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_292
timestamp 1607194113
transform 1 0 16716 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_295
timestamp 1607194113
transform 1 0 17636 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_294
timestamp 1607194113
transform 1 0 17544 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_297
timestamp 1607194113
transform 1 0 18464 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_296
timestamp 1607194113
transform 1 0 18372 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_299
timestamp 1607194113
transform 1 0 19292 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_298
timestamp 1607194113
transform 1 0 19200 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_302
timestamp 1607194113
transform 1 0 20856 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_301
timestamp 1607194113
transform 1 0 20120 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_300
timestamp 1607194113
transform 1 0 20028 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_304
timestamp 1607194113
transform 1 0 21684 0 -1 21056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILL_303
timestamp 1607194113
transform 1 0 20948 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILL_305
timestamp 1607194113
transform 1 0 22052 0 -1 21056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap37_0
timestamp 1607194113
transform 1 0 2732 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_1
timestamp 1607194113
transform 1 0 1904 0 1 21056
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_1_1
timestamp 1607194113
transform 1 0 3100 0 1 21056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap37_0
timestamp 1607194113
transform 1 0 2824 0 1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_307
timestamp 1607194113
transform 1 0 4388 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_306
timestamp 1607194113
transform 1 0 4296 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap37_1
timestamp 1607194113
transform 1 0 4020 0 1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap37_1
timestamp 1607194113
transform 1 0 3928 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_309
timestamp 1607194113
transform 1 0 5216 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_308
timestamp 1607194113
transform 1 0 5124 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_311
timestamp 1607194113
transform 1 0 6044 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_310
timestamp 1607194113
transform 1 0 5952 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_313
timestamp 1607194113
transform 1 0 6872 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_312
timestamp 1607194113
transform 1 0 6780 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_315
timestamp 1607194113
transform 1 0 7700 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_314
timestamp 1607194113
transform 1 0 7608 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_317
timestamp 1607194113
transform 1 0 8528 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_316
timestamp 1607194113
transform 1 0 8436 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_319
timestamp 1607194113
transform 1 0 9356 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_318
timestamp 1607194113
transform 1 0 9264 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_322
timestamp 1607194113
transform 1 0 10920 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_321
timestamp 1607194113
transform 1 0 10184 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_320
timestamp 1607194113
transform 1 0 10092 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_325
timestamp 1607194113
transform 1 0 11840 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_324
timestamp 1607194113
transform 1 0 11748 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_323
timestamp 1607194113
transform 1 0 11012 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_327
timestamp 1607194113
transform 1 0 12668 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_326
timestamp 1607194113
transform 1 0 12576 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_329
timestamp 1607194113
transform 1 0 13496 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_328
timestamp 1607194113
transform 1 0 13404 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_331
timestamp 1607194113
transform 1 0 14324 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_330
timestamp 1607194113
transform 1 0 14232 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_333
timestamp 1607194113
transform 1 0 15152 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_332
timestamp 1607194113
transform 1 0 15060 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_335
timestamp 1607194113
transform 1 0 15980 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_334
timestamp 1607194113
transform 1 0 15888 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_337
timestamp 1607194113
transform 1 0 16808 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_336
timestamp 1607194113
transform 1 0 16716 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_339
timestamp 1607194113
transform 1 0 17636 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_338
timestamp 1607194113
transform 1 0 17544 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_341
timestamp 1607194113
transform 1 0 18464 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_340
timestamp 1607194113
transform 1 0 18372 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_343
timestamp 1607194113
transform 1 0 19292 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_342
timestamp 1607194113
transform 1 0 19200 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_346
timestamp 1607194113
transform 1 0 20856 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_345
timestamp 1607194113
transform 1 0 20120 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_344
timestamp 1607194113
transform 1 0 20028 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_348
timestamp 1607194113
transform 1 0 21684 0 1 21056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILL_347
timestamp 1607194113
transform 1 0 20948 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILL_349
timestamp 1607194113
transform 1 0 22052 0 1 21056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap38_0
timestamp 1607194113
transform 1 0 2732 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_0
timestamp 1607194113
transform 1 0 1904 0 -1 22144
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  delay_0_0
timestamp 1607194113
transform 1 0 3100 0 -1 22144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  decap38_0
timestamp 1607194113
transform 1 0 2824 0 -1 22144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_351
timestamp 1607194113
transform 1 0 4388 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_350
timestamp 1607194113
transform 1 0 4296 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap38_1
timestamp 1607194113
transform 1 0 4020 0 -1 22144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap38_1
timestamp 1607194113
transform 1 0 3928 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_353
timestamp 1607194113
transform 1 0 5216 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_352
timestamp 1607194113
transform 1 0 5124 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_355
timestamp 1607194113
transform 1 0 6044 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_354
timestamp 1607194113
transform 1 0 5952 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_357
timestamp 1607194113
transform 1 0 6872 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_356
timestamp 1607194113
transform 1 0 6780 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_359
timestamp 1607194113
transform 1 0 7700 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_358
timestamp 1607194113
transform 1 0 7608 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_361
timestamp 1607194113
transform 1 0 8528 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_360
timestamp 1607194113
transform 1 0 8436 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_363
timestamp 1607194113
transform 1 0 9356 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_362
timestamp 1607194113
transform 1 0 9264 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_366
timestamp 1607194113
transform 1 0 10920 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_365
timestamp 1607194113
transform 1 0 10184 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_364
timestamp 1607194113
transform 1 0 10092 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_369
timestamp 1607194113
transform 1 0 11840 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_368
timestamp 1607194113
transform 1 0 11748 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_367
timestamp 1607194113
transform 1 0 11012 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_371
timestamp 1607194113
transform 1 0 12668 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_370
timestamp 1607194113
transform 1 0 12576 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_373
timestamp 1607194113
transform 1 0 13496 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_372
timestamp 1607194113
transform 1 0 13404 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_375
timestamp 1607194113
transform 1 0 14324 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_374
timestamp 1607194113
transform 1 0 14232 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_377
timestamp 1607194113
transform 1 0 15152 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_376
timestamp 1607194113
transform 1 0 15060 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_379
timestamp 1607194113
transform 1 0 15980 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_378
timestamp 1607194113
transform 1 0 15888 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_381
timestamp 1607194113
transform 1 0 16808 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_380
timestamp 1607194113
transform 1 0 16716 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_383
timestamp 1607194113
transform 1 0 17636 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_382
timestamp 1607194113
transform 1 0 17544 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_385
timestamp 1607194113
transform 1 0 18464 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_384
timestamp 1607194113
transform 1 0 18372 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_387
timestamp 1607194113
transform 1 0 19292 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_386
timestamp 1607194113
transform 1 0 19200 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_390
timestamp 1607194113
transform 1 0 20856 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_389
timestamp 1607194113
transform 1 0 20120 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_388
timestamp 1607194113
transform 1 0 20028 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_392
timestamp 1607194113
transform 1 0 21684 0 -1 22144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILL_391
timestamp 1607194113
transform 1 0 20948 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILL_393
timestamp 1607194113
transform 1 0 22052 0 -1 22144
box -38 -48 222 592
<< labels >>
rlabel metal3 s 800 800 920 920 6 inp_i
port 0 nsew default input
rlabel metal3 s 800 22016 920 22136 6 out_o
port 1 nsew default tristate
rlabel metal3 s 800 8960 920 9080 6 en_i[8]
port 2 nsew default input
rlabel metal3 s 800 13312 920 13432 6 en_i[7]
port 3 nsew default input
rlabel metal3 s 800 15488 920 15608 6 en_i[6]
port 4 nsew default input
rlabel metal3 s 800 16576 920 16696 6 en_i[5]
port 5 nsew default input
rlabel metal3 s 800 17664 920 17784 6 en_i[4]
port 6 nsew default input
rlabel metal3 s 800 18752 920 18872 6 en_i[3]
port 7 nsew default input
rlabel metal3 s 800 19840 920 19960 6 en_i[2]
port 8 nsew default input
rlabel metal3 s 800 20928 920 21048 6 en_i[1]
port 9 nsew default input
rlabel metal3 s 800 21472 920 21592 6 en_i[0]
port 10 nsew default input
rlabel metal5 s 1904 2560 22236 2880 6 VPWR
port 11 nsew default input
rlabel metal5 s 1904 20560 22236 20880 6 VGND
port 12 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23074 23185
<< end >>
